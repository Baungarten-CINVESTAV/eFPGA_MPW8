magic
tech sky130A
magscale 1 2
timestamp 1672417322
<< viali >>
rect 3985 37349 4019 37383
rect 25329 37349 25363 37383
rect 1593 37281 1627 37315
rect 11989 37281 12023 37315
rect 22017 37281 22051 37315
rect 23581 37281 23615 37315
rect 34897 37281 34931 37315
rect 38301 37281 38335 37315
rect 1869 37213 1903 37247
rect 2881 37213 2915 37247
rect 4169 37213 4203 37247
rect 4813 37213 4847 37247
rect 6009 37213 6043 37247
rect 6745 37213 6779 37247
rect 7573 37213 7607 37247
rect 8309 37213 8343 37247
rect 9781 37213 9815 37247
rect 11161 37213 11195 37247
rect 13093 37213 13127 37247
rect 13737 37213 13771 37247
rect 14289 37213 14323 37247
rect 15393 37213 15427 37247
rect 16037 37213 16071 37247
rect 16865 37213 16899 37247
rect 17509 37213 17543 37247
rect 18705 37213 18739 37247
rect 18797 37213 18831 37247
rect 19441 37213 19475 37247
rect 20085 37213 20119 37247
rect 21373 37213 21407 37247
rect 22293 37213 22327 37247
rect 23397 37213 23431 37247
rect 24593 37213 24627 37247
rect 25513 37213 25547 37247
rect 27353 37213 27387 37247
rect 27813 37213 27847 37247
rect 28733 37213 28767 37247
rect 29929 37213 29963 37247
rect 30573 37213 30607 37247
rect 31217 37213 31251 37247
rect 32321 37213 32355 37247
rect 33241 37213 33275 37247
rect 35173 37213 35207 37247
rect 36185 37213 36219 37247
rect 38117 37213 38151 37247
rect 11805 37145 11839 37179
rect 3065 37077 3099 37111
rect 4629 37077 4663 37111
rect 5825 37077 5859 37111
rect 6561 37077 6595 37111
rect 7757 37077 7791 37111
rect 8493 37077 8527 37111
rect 9965 37077 9999 37111
rect 10977 37077 11011 37111
rect 12909 37077 12943 37111
rect 13553 37077 13587 37111
rect 14473 37077 14507 37111
rect 15485 37077 15519 37111
rect 16221 37077 16255 37111
rect 16957 37077 16991 37111
rect 17693 37077 17727 37111
rect 19533 37077 19567 37111
rect 20269 37077 20303 37111
rect 21189 37077 21223 37111
rect 24777 37077 24811 37111
rect 25973 37077 26007 37111
rect 27169 37077 27203 37111
rect 27997 37077 28031 37111
rect 28549 37077 28583 37111
rect 29745 37077 29779 37111
rect 30389 37077 30423 37111
rect 31033 37077 31067 37111
rect 32505 37077 32539 37111
rect 33057 37077 33091 37111
rect 36369 37077 36403 37111
rect 1777 36873 1811 36907
rect 2329 36873 2363 36907
rect 22201 36873 22235 36907
rect 26157 36873 26191 36907
rect 35725 36873 35759 36907
rect 36829 36873 36863 36907
rect 8677 36805 8711 36839
rect 10241 36805 10275 36839
rect 15577 36805 15611 36839
rect 25145 36805 25179 36839
rect 27537 36805 27571 36839
rect 38117 36805 38151 36839
rect 1593 36737 1627 36771
rect 2513 36737 2547 36771
rect 2973 36737 3007 36771
rect 3801 36737 3835 36771
rect 4261 36737 4295 36771
rect 6745 36737 6779 36771
rect 10149 36737 10183 36771
rect 10977 36737 11011 36771
rect 12265 36737 12299 36771
rect 12909 36737 12943 36771
rect 13553 36737 13587 36771
rect 14197 36737 14231 36771
rect 14841 36737 14875 36771
rect 15485 36737 15519 36771
rect 16129 36737 16163 36771
rect 19349 36737 19383 36771
rect 20361 36737 20395 36771
rect 21005 36737 21039 36771
rect 22017 36737 22051 36771
rect 22937 36737 22971 36771
rect 23397 36737 23431 36771
rect 24041 36737 24075 36771
rect 26341 36737 26375 36771
rect 29101 36737 29135 36771
rect 29561 36737 29595 36771
rect 35081 36737 35115 36771
rect 35173 36737 35207 36771
rect 35909 36737 35943 36771
rect 36645 36737 36679 36771
rect 4905 36669 4939 36703
rect 8585 36669 8619 36703
rect 8861 36669 8895 36703
rect 16865 36669 16899 36703
rect 19441 36669 19475 36703
rect 24133 36669 24167 36703
rect 25053 36669 25087 36703
rect 25329 36669 25363 36703
rect 27445 36669 27479 36703
rect 28365 36669 28399 36703
rect 4353 36601 4387 36635
rect 12357 36601 12391 36635
rect 22753 36601 22787 36635
rect 28917 36601 28951 36635
rect 3065 36533 3099 36567
rect 3617 36533 3651 36567
rect 6837 36533 6871 36567
rect 11069 36533 11103 36567
rect 13001 36533 13035 36567
rect 13645 36533 13679 36567
rect 14289 36533 14323 36567
rect 14933 36533 14967 36567
rect 16221 36533 16255 36567
rect 17128 36533 17162 36567
rect 18613 36533 18647 36567
rect 20453 36533 20487 36567
rect 21097 36533 21131 36567
rect 23489 36533 23523 36567
rect 29653 36533 29687 36567
rect 38209 36533 38243 36567
rect 1593 36329 1627 36363
rect 3985 36329 4019 36363
rect 7941 36329 7975 36363
rect 26709 36329 26743 36363
rect 37473 36329 37507 36363
rect 4813 36193 4847 36227
rect 5825 36193 5859 36227
rect 6377 36193 6411 36227
rect 11989 36193 12023 36227
rect 15853 36193 15887 36227
rect 25513 36193 25547 36227
rect 25789 36193 25823 36227
rect 27537 36193 27571 36227
rect 1777 36125 1811 36159
rect 2881 36125 2915 36159
rect 4169 36125 4203 36159
rect 7849 36125 7883 36159
rect 11713 36125 11747 36159
rect 14565 36125 14599 36159
rect 15209 36125 15243 36159
rect 18705 36125 18739 36159
rect 19901 36125 19935 36159
rect 20637 36125 20671 36159
rect 24593 36125 24627 36159
rect 26617 36125 26651 36159
rect 28641 36125 28675 36159
rect 36369 36125 36403 36159
rect 37289 36125 37323 36159
rect 38025 36125 38059 36159
rect 4905 36057 4939 36091
rect 6469 36057 6503 36091
rect 7389 36057 7423 36091
rect 13737 36057 13771 36091
rect 14657 36057 14691 36091
rect 16129 36057 16163 36091
rect 21373 36057 21407 36091
rect 21465 36057 21499 36091
rect 22017 36057 22051 36091
rect 22569 36057 22603 36091
rect 22661 36057 22695 36091
rect 23581 36057 23615 36091
rect 25605 36057 25639 36091
rect 27629 36057 27663 36091
rect 28181 36057 28215 36091
rect 2697 35989 2731 36023
rect 9137 35989 9171 36023
rect 15301 35989 15335 36023
rect 17601 35989 17635 36023
rect 18797 35989 18831 36023
rect 19993 35989 20027 36023
rect 20729 35989 20763 36023
rect 24685 35989 24719 36023
rect 28733 35989 28767 36023
rect 36185 35989 36219 36023
rect 38209 35989 38243 36023
rect 3341 35785 3375 35819
rect 5917 35785 5951 35819
rect 14013 35785 14047 35819
rect 28825 35785 28859 35819
rect 7205 35717 7239 35751
rect 9413 35717 9447 35751
rect 20821 35717 20855 35751
rect 20913 35717 20947 35751
rect 23213 35717 23247 35751
rect 23305 35717 23339 35751
rect 25421 35717 25455 35751
rect 27261 35717 27295 35751
rect 5825 35649 5859 35683
rect 12449 35649 12483 35683
rect 13921 35649 13955 35683
rect 16865 35649 16899 35683
rect 19257 35649 19291 35683
rect 19901 35649 19935 35683
rect 21465 35649 21499 35683
rect 22477 35649 22511 35683
rect 24317 35649 24351 35683
rect 26433 35649 26467 35683
rect 27169 35649 27203 35683
rect 28089 35649 28123 35683
rect 28733 35649 28767 35683
rect 38025 35649 38059 35683
rect 1593 35581 1627 35615
rect 1869 35581 1903 35615
rect 6929 35581 6963 35615
rect 9137 35581 9171 35615
rect 11161 35581 11195 35615
rect 14565 35581 14599 35615
rect 14841 35581 14875 35615
rect 17141 35581 17175 35615
rect 23489 35581 23523 35615
rect 25329 35581 25363 35615
rect 25605 35581 25639 35615
rect 12541 35513 12575 35547
rect 16313 35513 16347 35547
rect 8677 35445 8711 35479
rect 18613 35445 18647 35479
rect 19349 35445 19383 35479
rect 19993 35445 20027 35479
rect 22569 35445 22603 35479
rect 24409 35445 24443 35479
rect 26525 35445 26559 35479
rect 28181 35445 28215 35479
rect 38209 35445 38243 35479
rect 1777 35241 1811 35275
rect 24685 35241 24719 35275
rect 35081 35241 35115 35275
rect 9781 35173 9815 35207
rect 14289 35173 14323 35207
rect 25421 35173 25455 35207
rect 4629 35105 4663 35139
rect 6377 35105 6411 35139
rect 9229 35105 9263 35139
rect 11989 35105 12023 35139
rect 15761 35105 15795 35139
rect 26341 35105 26375 35139
rect 26617 35105 26651 35139
rect 28457 35105 28491 35139
rect 1593 35037 1627 35071
rect 8585 35037 8619 35071
rect 11713 35037 11747 35071
rect 14473 35037 14507 35071
rect 18705 35037 18739 35071
rect 19901 35037 19935 35071
rect 20545 35037 20579 35071
rect 21189 35037 21223 35071
rect 21833 35037 21867 35071
rect 24593 35037 24627 35071
rect 25329 35037 25363 35071
rect 35265 35037 35299 35071
rect 37657 35037 37691 35071
rect 4905 34969 4939 35003
rect 9321 34969 9355 35003
rect 13737 34969 13771 35003
rect 16037 34969 16071 35003
rect 17785 34969 17819 35003
rect 23029 34969 23063 35003
rect 23121 34969 23155 35003
rect 24041 34969 24075 35003
rect 26433 34969 26467 35003
rect 28181 34969 28215 35003
rect 28273 34969 28307 35003
rect 8401 34901 8435 34935
rect 18797 34901 18831 34935
rect 19993 34901 20027 34935
rect 20637 34901 20671 34935
rect 21281 34901 21315 34935
rect 21925 34901 21959 34935
rect 37473 34901 37507 34935
rect 1593 34697 1627 34731
rect 9597 34697 9631 34731
rect 19349 34697 19383 34731
rect 24041 34697 24075 34731
rect 26525 34697 26559 34731
rect 28365 34697 28399 34731
rect 5641 34629 5675 34663
rect 20177 34629 20211 34663
rect 22477 34629 22511 34663
rect 22569 34629 22603 34663
rect 24685 34629 24719 34663
rect 24777 34629 24811 34663
rect 25329 34629 25363 34663
rect 27353 34629 27387 34663
rect 1777 34561 1811 34595
rect 5549 34561 5583 34595
rect 9781 34561 9815 34595
rect 17325 34561 17359 34595
rect 17417 34561 17451 34595
rect 17969 34561 18003 34595
rect 18613 34561 18647 34595
rect 19257 34561 19291 34595
rect 20085 34561 20119 34595
rect 20729 34561 20763 34595
rect 23949 34561 23983 34595
rect 26433 34561 26467 34595
rect 38025 34561 38059 34595
rect 3249 34493 3283 34527
rect 11713 34493 11747 34527
rect 11989 34493 12023 34527
rect 13737 34493 13771 34527
rect 18061 34493 18095 34527
rect 18705 34493 18739 34527
rect 20821 34493 20855 34527
rect 23489 34493 23523 34527
rect 27261 34493 27295 34527
rect 27905 34493 27939 34527
rect 3512 34357 3546 34391
rect 4997 34357 5031 34391
rect 38209 34357 38243 34391
rect 18797 34153 18831 34187
rect 22109 34153 22143 34187
rect 36645 34153 36679 34187
rect 27813 34085 27847 34119
rect 5641 34017 5675 34051
rect 9413 34017 9447 34051
rect 9689 34017 9723 34051
rect 11886 34017 11920 34051
rect 15301 34017 15335 34051
rect 17325 34017 17359 34051
rect 23397 34017 23431 34051
rect 27261 34017 27295 34051
rect 1593 33949 1627 33983
rect 2513 33949 2547 33983
rect 18061 33949 18095 33983
rect 18153 33949 18187 33983
rect 18705 33949 18739 33983
rect 19533 33949 19567 33983
rect 20821 33949 20855 33983
rect 22017 33949 22051 33983
rect 25237 33949 25271 33983
rect 28365 33949 28399 33983
rect 36829 33949 36863 33983
rect 5917 33881 5951 33915
rect 12173 33881 12207 33915
rect 15577 33881 15611 33915
rect 22753 33881 22787 33915
rect 22845 33881 22879 33915
rect 27353 33881 27387 33915
rect 1777 33813 1811 33847
rect 2329 33813 2363 33847
rect 7389 33813 7423 33847
rect 11161 33813 11195 33847
rect 13645 33813 13679 33847
rect 19625 33813 19659 33847
rect 20177 33813 20211 33847
rect 20913 33813 20947 33847
rect 25329 33813 25363 33847
rect 28457 33813 28491 33847
rect 6009 33609 6043 33643
rect 23857 33609 23891 33643
rect 25145 33609 25179 33643
rect 25789 33609 25823 33643
rect 28457 33609 28491 33643
rect 10425 33541 10459 33575
rect 13001 33541 13035 33575
rect 20453 33541 20487 33575
rect 20545 33541 20579 33575
rect 22845 33541 22879 33575
rect 23765 33541 23799 33575
rect 27353 33541 27387 33575
rect 2053 33473 2087 33507
rect 4261 33473 4295 33507
rect 7481 33473 7515 33507
rect 9689 33473 9723 33507
rect 16865 33473 16899 33507
rect 19533 33473 19567 33507
rect 22753 33473 22787 33507
rect 24409 33473 24443 33507
rect 25053 33473 25087 33507
rect 25697 33473 25731 33507
rect 28365 33473 28399 33507
rect 29009 33473 29043 33507
rect 29653 33473 29687 33507
rect 2329 33405 2363 33439
rect 3801 33405 3835 33439
rect 4537 33405 4571 33439
rect 7757 33405 7791 33439
rect 12725 33405 12759 33439
rect 14749 33405 14783 33439
rect 17141 33405 17175 33439
rect 21465 33405 21499 33439
rect 27261 33405 27295 33439
rect 27905 33405 27939 33439
rect 9229 33269 9263 33303
rect 18613 33269 18647 33303
rect 19625 33269 19659 33303
rect 24501 33269 24535 33303
rect 29101 33269 29135 33303
rect 29745 33269 29779 33303
rect 2053 33065 2087 33099
rect 8493 33065 8527 33099
rect 25329 33065 25363 33099
rect 19901 32997 19935 33031
rect 24685 32997 24719 33031
rect 6745 32929 6779 32963
rect 15209 32929 15243 32963
rect 15853 32929 15887 32963
rect 20545 32929 20579 32963
rect 21281 32929 21315 32963
rect 26433 32929 26467 32963
rect 27721 32929 27755 32963
rect 2053 32861 2087 32895
rect 10977 32861 11011 32895
rect 19809 32861 19843 32895
rect 20453 32861 20487 32895
rect 23305 32861 23339 32895
rect 24593 32861 24627 32895
rect 25237 32861 25271 32895
rect 38025 32861 38059 32895
rect 7021 32793 7055 32827
rect 11253 32793 11287 32827
rect 13001 32793 13035 32827
rect 14473 32793 14507 32827
rect 16129 32793 16163 32827
rect 21373 32793 21407 32827
rect 22293 32793 22327 32827
rect 26157 32793 26191 32827
rect 26249 32793 26283 32827
rect 27813 32793 27847 32827
rect 28733 32793 28767 32827
rect 17601 32725 17635 32759
rect 23397 32725 23431 32759
rect 38209 32725 38243 32759
rect 7297 32453 7331 32487
rect 9689 32453 9723 32487
rect 11989 32453 12023 32487
rect 14749 32453 14783 32487
rect 19970 32453 20004 32487
rect 23581 32453 23615 32487
rect 25145 32453 25179 32487
rect 27261 32453 27295 32487
rect 29009 32453 29043 32487
rect 1685 32385 1719 32419
rect 6561 32385 6595 32419
rect 9413 32385 9447 32419
rect 14473 32385 14507 32419
rect 16865 32385 16899 32419
rect 19165 32385 19199 32419
rect 22017 32385 22051 32419
rect 22845 32385 22879 32419
rect 26249 32385 26283 32419
rect 27169 32385 27203 32419
rect 28917 32385 28951 32419
rect 38025 32385 38059 32419
rect 12725 32317 12759 32351
rect 17141 32317 17175 32351
rect 19901 32317 19935 32351
rect 20269 32317 20303 32351
rect 23489 32317 23523 32351
rect 24041 32317 24075 32351
rect 25053 32317 25087 32351
rect 27813 32317 27847 32351
rect 27997 32317 28031 32351
rect 1869 32249 1903 32283
rect 22109 32249 22143 32283
rect 22661 32249 22695 32283
rect 25605 32249 25639 32283
rect 11161 32181 11195 32215
rect 16221 32181 16255 32215
rect 18613 32181 18647 32215
rect 19257 32181 19291 32215
rect 26341 32181 26375 32215
rect 28181 32181 28215 32215
rect 38209 32181 38243 32215
rect 27629 31977 27663 32011
rect 29009 31977 29043 32011
rect 7021 31909 7055 31943
rect 5273 31841 5307 31875
rect 5549 31841 5583 31875
rect 9137 31841 9171 31875
rect 9413 31841 9447 31875
rect 16037 31841 16071 31875
rect 17785 31841 17819 31875
rect 19533 31841 19567 31875
rect 20177 31841 20211 31875
rect 23305 31841 23339 31875
rect 26065 31841 26099 31875
rect 27077 31841 27111 31875
rect 1593 31773 1627 31807
rect 2329 31773 2363 31807
rect 2421 31773 2455 31807
rect 11989 31773 12023 31807
rect 18705 31773 18739 31807
rect 20637 31773 20671 31807
rect 25329 31773 25363 31807
rect 27537 31773 27571 31807
rect 28917 31773 28951 31807
rect 11161 31705 11195 31739
rect 12265 31705 12299 31739
rect 16313 31705 16347 31739
rect 19625 31705 19659 31739
rect 20729 31705 20763 31739
rect 23029 31705 23063 31739
rect 23121 31705 23155 31739
rect 26157 31705 26191 31739
rect 1777 31637 1811 31671
rect 13737 31637 13771 31671
rect 18797 31637 18831 31671
rect 25421 31637 25455 31671
rect 28181 31637 28215 31671
rect 20545 31433 20579 31467
rect 21373 31433 21407 31467
rect 23949 31433 23983 31467
rect 28089 31433 28123 31467
rect 29837 31433 29871 31467
rect 3341 31365 3375 31399
rect 13737 31365 13771 31399
rect 17877 31365 17911 31399
rect 25329 31365 25363 31399
rect 3065 31297 3099 31331
rect 11713 31297 11747 31331
rect 19809 31297 19843 31331
rect 20453 31297 20487 31331
rect 21281 31297 21315 31331
rect 22017 31297 22051 31331
rect 23397 31297 23431 31331
rect 23857 31297 23891 31331
rect 27445 31297 27479 31331
rect 30021 31297 30055 31331
rect 30665 31297 30699 31331
rect 7665 31229 7699 31263
rect 7941 31229 7975 31263
rect 11989 31229 12023 31263
rect 17049 31229 17083 31263
rect 17785 31229 17819 31263
rect 18797 31229 18831 31263
rect 22201 31229 22235 31263
rect 25237 31229 25271 31263
rect 26157 31229 26191 31263
rect 27629 31229 27663 31263
rect 23213 31161 23247 31195
rect 30481 31161 30515 31195
rect 4813 31093 4847 31127
rect 9413 31093 9447 31127
rect 19901 31093 19935 31127
rect 22569 31093 22603 31127
rect 19901 30889 19935 30923
rect 23765 30889 23799 30923
rect 12173 30821 12207 30855
rect 4261 30753 4295 30787
rect 6377 30753 6411 30787
rect 6653 30753 6687 30787
rect 10425 30753 10459 30787
rect 15853 30753 15887 30787
rect 16129 30753 16163 30787
rect 21649 30753 21683 30787
rect 22109 30753 22143 30787
rect 26249 30753 26283 30787
rect 27905 30753 27939 30787
rect 3985 30685 4019 30719
rect 18705 30685 18739 30719
rect 19809 30685 19843 30719
rect 20913 30685 20947 30719
rect 23121 30685 23155 30719
rect 23949 30685 23983 30719
rect 28089 30685 28123 30719
rect 38301 30685 38335 30719
rect 10701 30617 10735 30651
rect 21741 30617 21775 30651
rect 26341 30617 26375 30651
rect 27261 30617 27295 30651
rect 5733 30549 5767 30583
rect 8125 30549 8159 30583
rect 17601 30549 17635 30583
rect 18797 30549 18831 30583
rect 21005 30549 21039 30583
rect 23213 30549 23247 30583
rect 28549 30549 28583 30583
rect 38117 30549 38151 30583
rect 29285 30345 29319 30379
rect 9873 30277 9907 30311
rect 16129 30277 16163 30311
rect 24225 30277 24259 30311
rect 24961 30277 24995 30311
rect 27261 30277 27295 30311
rect 1593 30209 1627 30243
rect 7573 30209 7607 30243
rect 15393 30209 15427 30243
rect 16865 30209 16899 30243
rect 19441 30209 19475 30243
rect 20085 30209 20119 30243
rect 20729 30209 20763 30243
rect 22201 30209 22235 30243
rect 22293 30209 22327 30243
rect 23397 30209 23431 30243
rect 24133 30209 24167 30243
rect 26341 30209 26375 30243
rect 27169 30209 27203 30243
rect 28641 30209 28675 30243
rect 29469 30209 29503 30243
rect 10609 30141 10643 30175
rect 12817 30141 12851 30175
rect 13093 30141 13127 30175
rect 17141 30141 17175 30175
rect 20177 30141 20211 30175
rect 23489 30141 23523 30175
rect 24869 30141 24903 30175
rect 25789 30141 25823 30175
rect 1777 30005 1811 30039
rect 7836 30005 7870 30039
rect 9321 30005 9355 30039
rect 14565 30005 14599 30039
rect 18613 30005 18647 30039
rect 19533 30005 19567 30039
rect 20821 30005 20855 30039
rect 26433 30005 26467 30039
rect 28733 30005 28767 30039
rect 4721 29801 4755 29835
rect 22385 29801 22419 29835
rect 28549 29801 28583 29835
rect 29745 29801 29779 29835
rect 34897 29801 34931 29835
rect 10885 29733 10919 29767
rect 16037 29665 16071 29699
rect 21097 29665 21131 29699
rect 24961 29665 24995 29699
rect 25973 29665 26007 29699
rect 28181 29665 28215 29699
rect 37749 29665 37783 29699
rect 4629 29597 4663 29631
rect 9137 29597 9171 29631
rect 11345 29597 11379 29631
rect 18705 29597 18739 29631
rect 18797 29597 18831 29631
rect 19441 29597 19475 29631
rect 20269 29597 20303 29631
rect 21005 29597 21039 29631
rect 21649 29597 21683 29631
rect 22293 29597 22327 29631
rect 22937 29597 22971 29631
rect 23581 29597 23615 29631
rect 26433 29597 26467 29631
rect 27077 29597 27111 29631
rect 27997 29597 28031 29631
rect 29929 29597 29963 29631
rect 30757 29597 30791 29631
rect 30849 29597 30883 29631
rect 35081 29597 35115 29631
rect 37473 29597 37507 29631
rect 9413 29529 9447 29563
rect 12081 29529 12115 29563
rect 16313 29529 16347 29563
rect 21741 29529 21775 29563
rect 25053 29529 25087 29563
rect 17785 29461 17819 29495
rect 19533 29461 19567 29495
rect 20085 29461 20119 29495
rect 23029 29461 23063 29495
rect 23673 29461 23707 29495
rect 26525 29461 26559 29495
rect 27169 29461 27203 29495
rect 13461 29257 13495 29291
rect 4997 29189 5031 29223
rect 18153 29189 18187 29223
rect 20545 29189 20579 29223
rect 21465 29189 21499 29223
rect 23949 29189 23983 29223
rect 25697 29189 25731 29223
rect 1777 29121 1811 29155
rect 2421 29121 2455 29155
rect 4445 29121 4479 29155
rect 9321 29121 9355 29155
rect 11713 29121 11747 29155
rect 14473 29121 14507 29155
rect 19717 29121 19751 29155
rect 22661 29121 22695 29155
rect 27169 29121 27203 29155
rect 5733 29053 5767 29087
rect 11069 29053 11103 29087
rect 18061 29053 18095 29087
rect 18429 29053 18463 29087
rect 19809 29053 19843 29087
rect 20453 29053 20487 29087
rect 23857 29053 23891 29087
rect 24869 29053 24903 29087
rect 25605 29053 25639 29087
rect 26617 29053 26651 29087
rect 27261 29053 27295 29087
rect 27813 29053 27847 29087
rect 27997 29053 28031 29087
rect 22753 28985 22787 29019
rect 28457 28985 28491 29019
rect 1593 28917 1627 28951
rect 2684 28917 2718 28951
rect 9584 28917 9618 28951
rect 11976 28917 12010 28951
rect 14736 28917 14770 28951
rect 16221 28917 16255 28951
rect 13369 28713 13403 28747
rect 17601 28713 17635 28747
rect 21189 28713 21223 28747
rect 22385 28713 22419 28747
rect 19533 28645 19567 28679
rect 6929 28577 6963 28611
rect 11621 28577 11655 28611
rect 15853 28577 15887 28611
rect 23029 28577 23063 28611
rect 25329 28577 25363 28611
rect 25973 28577 26007 28611
rect 27813 28577 27847 28611
rect 31309 28577 31343 28611
rect 1869 28509 1903 28543
rect 4905 28509 4939 28543
rect 19441 28509 19475 28543
rect 20085 28509 20119 28543
rect 21097 28509 21131 28543
rect 21741 28509 21775 28543
rect 21925 28509 21959 28543
rect 24593 28509 24627 28543
rect 24685 28509 24719 28543
rect 25237 28509 25271 28543
rect 28641 28509 28675 28543
rect 31217 28509 31251 28543
rect 5181 28441 5215 28475
rect 11897 28441 11931 28475
rect 16129 28441 16163 28475
rect 23121 28441 23155 28475
rect 24041 28441 24075 28475
rect 26065 28441 26099 28475
rect 26985 28441 27019 28475
rect 27537 28441 27571 28475
rect 27629 28441 27663 28475
rect 28733 28441 28767 28475
rect 31953 28441 31987 28475
rect 32045 28441 32079 28475
rect 32965 28441 32999 28475
rect 1961 28373 1995 28407
rect 20177 28373 20211 28407
rect 11069 28169 11103 28203
rect 21281 28169 21315 28203
rect 24961 28169 24995 28203
rect 25605 28169 25639 28203
rect 27353 28101 27387 28135
rect 9321 28033 9355 28067
rect 15853 28033 15887 28067
rect 19257 28033 19291 28067
rect 19901 28033 19935 28067
rect 20545 28033 20579 28067
rect 21189 28033 21223 28067
rect 22845 28033 22879 28067
rect 23305 28033 23339 28067
rect 24225 28033 24259 28067
rect 24869 28033 24903 28067
rect 25513 28033 25547 28067
rect 26341 28033 26375 28067
rect 38301 28033 38335 28067
rect 3249 27965 3283 27999
rect 3525 27965 3559 27999
rect 4997 27965 5031 27999
rect 9597 27965 9631 27999
rect 13829 27965 13863 27999
rect 15577 27965 15611 27999
rect 19993 27965 20027 27999
rect 22201 27965 22235 27999
rect 22385 27965 22419 27999
rect 24317 27965 24351 27999
rect 27261 27965 27295 27999
rect 23397 27897 23431 27931
rect 27813 27897 27847 27931
rect 13553 27829 13587 27863
rect 19349 27829 19383 27863
rect 20637 27829 20671 27863
rect 26157 27829 26191 27863
rect 38117 27829 38151 27863
rect 10590 27625 10624 27659
rect 7021 27557 7055 27591
rect 29837 27557 29871 27591
rect 5273 27489 5307 27523
rect 10333 27489 10367 27523
rect 12357 27489 12391 27523
rect 17601 27489 17635 27523
rect 22109 27489 22143 27523
rect 23121 27489 23155 27523
rect 25881 27489 25915 27523
rect 1593 27421 1627 27455
rect 21189 27421 21223 27455
rect 23581 27421 23615 27455
rect 24593 27421 24627 27455
rect 29745 27421 29779 27455
rect 38025 27421 38059 27455
rect 5549 27353 5583 27387
rect 17693 27353 17727 27387
rect 18613 27353 18647 27387
rect 19717 27353 19751 27387
rect 19809 27353 19843 27387
rect 20729 27353 20763 27387
rect 22194 27353 22228 27387
rect 25973 27353 26007 27387
rect 26893 27353 26927 27387
rect 1777 27285 1811 27319
rect 21281 27285 21315 27319
rect 23673 27285 23707 27319
rect 24685 27285 24719 27319
rect 38209 27285 38243 27319
rect 1593 27081 1627 27115
rect 17417 27081 17451 27115
rect 20913 27081 20947 27115
rect 34161 27081 34195 27115
rect 4537 27013 4571 27047
rect 9413 27013 9447 27047
rect 10977 27013 11011 27047
rect 18153 27013 18187 27047
rect 22109 27013 22143 27047
rect 23857 27013 23891 27047
rect 24961 27013 24995 27047
rect 27353 27013 27387 27047
rect 1777 26945 1811 26979
rect 17325 26945 17359 26979
rect 19533 26945 19567 26979
rect 20177 26945 20211 26979
rect 20821 26945 20855 26979
rect 22017 26945 22051 26979
rect 22661 26945 22695 26979
rect 25789 26945 25823 26979
rect 28365 26945 28399 26979
rect 29193 26945 29227 26979
rect 34345 26945 34379 26979
rect 4261 26877 4295 26911
rect 7205 26877 7239 26911
rect 7481 26877 7515 26911
rect 18061 26877 18095 26911
rect 19073 26877 19107 26911
rect 23765 26877 23799 26911
rect 24041 26877 24075 26911
rect 27261 26877 27295 26911
rect 29285 26877 29319 26911
rect 22753 26809 22787 26843
rect 25605 26809 25639 26843
rect 27813 26809 27847 26843
rect 6009 26741 6043 26775
rect 8953 26741 8987 26775
rect 19625 26741 19659 26775
rect 20269 26741 20303 26775
rect 25053 26741 25087 26775
rect 28457 26741 28491 26775
rect 8493 26537 8527 26571
rect 16024 26537 16058 26571
rect 18797 26537 18831 26571
rect 25053 26537 25087 26571
rect 25697 26537 25731 26571
rect 31953 26537 31987 26571
rect 38117 26537 38151 26571
rect 13737 26469 13771 26503
rect 26893 26469 26927 26503
rect 2145 26401 2179 26435
rect 7021 26401 7055 26435
rect 23213 26401 23247 26435
rect 26341 26401 26375 26435
rect 6745 26333 6779 26367
rect 11989 26333 12023 26367
rect 15761 26333 15795 26367
rect 18705 26333 18739 26367
rect 23121 26333 23155 26367
rect 23765 26333 23799 26367
rect 23857 26333 23891 26367
rect 24961 26333 24995 26367
rect 25605 26333 25639 26367
rect 31861 26333 31895 26367
rect 38301 26333 38335 26367
rect 2237 26265 2271 26299
rect 3157 26265 3191 26299
rect 12265 26265 12299 26299
rect 17785 26265 17819 26299
rect 19533 26265 19567 26299
rect 19625 26265 19659 26299
rect 20545 26265 20579 26299
rect 26433 26265 26467 26299
rect 32597 26265 32631 26299
rect 32689 26265 32723 26299
rect 33241 26265 33275 26299
rect 3065 25993 3099 26027
rect 5365 25993 5399 26027
rect 19717 25993 19751 26027
rect 22201 25993 22235 26027
rect 32689 25993 32723 26027
rect 2973 25857 3007 25891
rect 7941 25857 7975 25891
rect 19625 25857 19659 25891
rect 20269 25857 20303 25891
rect 21281 25857 21315 25891
rect 22109 25857 22143 25891
rect 22937 25857 22971 25891
rect 23397 25857 23431 25891
rect 28273 25857 28307 25891
rect 29101 25857 29135 25891
rect 29193 25857 29227 25891
rect 31217 25857 31251 25891
rect 3617 25789 3651 25823
rect 3893 25789 3927 25823
rect 8677 25789 8711 25823
rect 9321 25789 9355 25823
rect 9597 25789 9631 25823
rect 11713 25789 11747 25823
rect 11989 25789 12023 25823
rect 13461 25789 13495 25823
rect 16865 25789 16899 25823
rect 17141 25789 17175 25823
rect 23489 25789 23523 25823
rect 29929 25789 29963 25823
rect 30113 25789 30147 25823
rect 31033 25789 31067 25823
rect 22753 25721 22787 25755
rect 11069 25653 11103 25687
rect 18613 25653 18647 25687
rect 20361 25653 20395 25687
rect 21373 25653 21407 25687
rect 28089 25653 28123 25687
rect 30573 25653 30607 25687
rect 31401 25653 31435 25687
rect 10885 25449 10919 25483
rect 21925 25449 21959 25483
rect 29745 25449 29779 25483
rect 17693 25381 17727 25415
rect 27169 25381 27203 25415
rect 6745 25313 6779 25347
rect 7021 25313 7055 25347
rect 9137 25313 9171 25347
rect 9413 25313 9447 25347
rect 12081 25313 12115 25347
rect 21281 25313 21315 25347
rect 1685 25245 1719 25279
rect 11805 25245 11839 25279
rect 15945 25245 15979 25279
rect 18705 25245 18739 25279
rect 19441 25245 19475 25279
rect 20637 25245 20671 25279
rect 21465 25245 21499 25279
rect 27353 25245 27387 25279
rect 28549 25245 28583 25279
rect 29193 25245 29227 25279
rect 29929 25245 29963 25279
rect 1869 25177 1903 25211
rect 16221 25177 16255 25211
rect 19717 25177 19751 25211
rect 8493 25109 8527 25143
rect 13553 25109 13587 25143
rect 18797 25109 18831 25143
rect 20729 25109 20763 25143
rect 28365 25109 28399 25143
rect 29009 25109 29043 25143
rect 17049 24837 17083 24871
rect 22937 24837 22971 24871
rect 27537 24837 27571 24871
rect 1777 24769 1811 24803
rect 4721 24769 4755 24803
rect 8401 24769 8435 24803
rect 11713 24769 11747 24803
rect 13093 24769 13127 24803
rect 13185 24769 13219 24803
rect 18797 24769 18831 24803
rect 19073 24769 19107 24803
rect 20269 24769 20303 24803
rect 20905 24769 20939 24803
rect 21005 24769 21039 24803
rect 23949 24769 23983 24803
rect 25605 24769 25639 24803
rect 38025 24769 38059 24803
rect 5457 24701 5491 24735
rect 8677 24701 8711 24735
rect 12449 24701 12483 24735
rect 14105 24701 14139 24735
rect 14381 24701 14415 24735
rect 16957 24701 16991 24735
rect 17233 24701 17267 24735
rect 22845 24701 22879 24735
rect 24041 24701 24075 24735
rect 27445 24701 27479 24735
rect 28365 24701 28399 24735
rect 29009 24701 29043 24735
rect 10149 24633 10183 24667
rect 23397 24633 23431 24667
rect 1593 24565 1627 24599
rect 15853 24565 15887 24599
rect 20361 24565 20395 24599
rect 25697 24565 25731 24599
rect 38209 24565 38243 24599
rect 1685 24225 1719 24259
rect 3985 24225 4019 24259
rect 20269 24225 20303 24259
rect 22845 24225 22879 24259
rect 28549 24225 28583 24259
rect 29193 24225 29227 24259
rect 6009 24157 6043 24191
rect 6469 24157 6503 24191
rect 15393 24157 15427 24191
rect 21097 24157 21131 24191
rect 24593 24157 24627 24191
rect 27997 24157 28031 24191
rect 38025 24157 38059 24191
rect 1961 24089 1995 24123
rect 4261 24089 4295 24123
rect 6745 24089 6779 24123
rect 15669 24089 15703 24123
rect 19625 24089 19659 24123
rect 19717 24089 19751 24123
rect 21833 24089 21867 24123
rect 21925 24089 21959 24123
rect 28641 24089 28675 24123
rect 3433 24021 3467 24055
rect 8217 24021 8251 24055
rect 17141 24021 17175 24055
rect 18245 24021 18279 24055
rect 21189 24021 21223 24055
rect 24685 24021 24719 24055
rect 27813 24021 27847 24055
rect 38209 24021 38243 24055
rect 16957 23817 16991 23851
rect 23673 23817 23707 23851
rect 4537 23749 4571 23783
rect 15393 23749 15427 23783
rect 18153 23749 18187 23783
rect 18254 23749 18288 23783
rect 18797 23749 18831 23783
rect 20637 23749 20671 23783
rect 24317 23749 24351 23783
rect 25605 23749 25639 23783
rect 25697 23749 25731 23783
rect 27721 23749 27755 23783
rect 27813 23749 27847 23783
rect 1961 23681 1995 23715
rect 2605 23681 2639 23715
rect 4261 23681 4295 23715
rect 7941 23681 7975 23715
rect 16865 23681 16899 23715
rect 20545 23681 20579 23715
rect 22017 23681 22051 23715
rect 22661 23681 22695 23715
rect 23581 23681 23615 23715
rect 34253 23681 34287 23715
rect 8217 23613 8251 23647
rect 16129 23613 16163 23647
rect 22109 23613 22143 23647
rect 26617 23613 26651 23647
rect 27997 23613 28031 23647
rect 29377 23613 29411 23647
rect 22753 23545 22787 23579
rect 1777 23477 1811 23511
rect 2421 23477 2455 23511
rect 6009 23477 6043 23511
rect 9689 23477 9723 23511
rect 24409 23477 24443 23511
rect 34345 23477 34379 23511
rect 28549 23273 28583 23307
rect 5733 23137 5767 23171
rect 6009 23137 6043 23171
rect 10793 23137 10827 23171
rect 17509 23137 17543 23171
rect 25973 23137 26007 23171
rect 29837 23137 29871 23171
rect 1685 23069 1719 23103
rect 10517 23069 10551 23103
rect 15485 23069 15519 23103
rect 19441 23069 19475 23103
rect 21005 23069 21039 23103
rect 26157 23069 26191 23103
rect 28181 23069 28215 23103
rect 28365 23069 28399 23103
rect 1961 23001 1995 23035
rect 15761 23001 15795 23035
rect 19717 23001 19751 23035
rect 29929 23001 29963 23035
rect 30849 23001 30883 23035
rect 3433 22933 3467 22967
rect 7481 22933 7515 22967
rect 12265 22933 12299 22967
rect 21097 22933 21131 22967
rect 26617 22933 26651 22967
rect 3341 22729 3375 22763
rect 25789 22729 25823 22763
rect 28733 22729 28767 22763
rect 31125 22729 31159 22763
rect 1869 22661 1903 22695
rect 9597 22661 9631 22695
rect 15301 22661 15335 22695
rect 21189 22661 21223 22695
rect 22201 22661 22235 22695
rect 26525 22661 26559 22695
rect 27353 22661 27387 22695
rect 28273 22661 28307 22695
rect 13277 22593 13311 22627
rect 17877 22593 17911 22627
rect 18521 22593 18555 22627
rect 19441 22593 19475 22627
rect 21097 22593 21131 22627
rect 25973 22593 26007 22627
rect 26433 22593 26467 22627
rect 28917 22593 28951 22627
rect 31309 22593 31343 22627
rect 34437 22593 34471 22627
rect 38025 22593 38059 22627
rect 1593 22525 1627 22559
rect 4261 22525 4295 22559
rect 4537 22525 4571 22559
rect 9321 22525 9355 22559
rect 13553 22525 13587 22559
rect 18797 22525 18831 22559
rect 19625 22525 19659 22559
rect 22109 22525 22143 22559
rect 27261 22525 27295 22559
rect 11069 22457 11103 22491
rect 22661 22457 22695 22491
rect 34253 22457 34287 22491
rect 38209 22457 38243 22491
rect 6009 22389 6043 22423
rect 17969 22389 18003 22423
rect 5352 22185 5386 22219
rect 9400 22185 9434 22219
rect 12160 22185 12194 22219
rect 26157 22185 26191 22219
rect 5089 22049 5123 22083
rect 6837 22049 6871 22083
rect 11897 22049 11931 22083
rect 13645 22049 13679 22083
rect 21373 22049 21407 22083
rect 29837 22049 29871 22083
rect 9137 21981 9171 22015
rect 18429 21981 18463 22015
rect 19441 21981 19475 22015
rect 20085 21981 20119 22015
rect 22569 21981 22603 22015
rect 23213 21981 23247 22015
rect 23857 21981 23891 22015
rect 26341 21981 26375 22015
rect 29745 21981 29779 22015
rect 1685 21913 1719 21947
rect 1869 21913 1903 21947
rect 18705 21913 18739 21947
rect 20361 21913 20395 21947
rect 21097 21913 21131 21947
rect 21189 21913 21223 21947
rect 23305 21913 23339 21947
rect 24685 21913 24719 21947
rect 24777 21913 24811 21947
rect 25697 21913 25731 21947
rect 10885 21845 10919 21879
rect 19533 21845 19567 21879
rect 22661 21845 22695 21879
rect 23949 21845 23983 21879
rect 21281 21641 21315 21675
rect 24041 21641 24075 21675
rect 31493 21641 31527 21675
rect 5089 21573 5123 21607
rect 7757 21573 7791 21607
rect 18337 21505 18371 21539
rect 18981 21505 19015 21539
rect 19901 21505 19935 21539
rect 22017 21505 22051 21539
rect 23305 21505 23339 21539
rect 23949 21505 23983 21539
rect 24593 21505 24627 21539
rect 28089 21505 28123 21539
rect 29193 21505 29227 21539
rect 31677 21505 31711 21539
rect 38025 21505 38059 21539
rect 5825 21437 5859 21471
rect 7481 21437 7515 21471
rect 14473 21437 14507 21471
rect 19165 21437 19199 21471
rect 20637 21437 20671 21471
rect 22293 21437 22327 21471
rect 28273 21437 28307 21471
rect 16221 21369 16255 21403
rect 28457 21369 28491 21403
rect 9229 21301 9263 21335
rect 14736 21301 14770 21335
rect 18429 21301 18463 21335
rect 23397 21301 23431 21335
rect 24685 21301 24719 21335
rect 29285 21301 29319 21335
rect 38209 21301 38243 21335
rect 5352 21097 5386 21131
rect 21281 21097 21315 21131
rect 28365 21097 28399 21131
rect 29101 21097 29135 21131
rect 16681 21029 16715 21063
rect 5089 20961 5123 20995
rect 6837 20961 6871 20995
rect 9137 20961 9171 20995
rect 9413 20961 9447 20995
rect 20545 20961 20579 20995
rect 25881 20961 25915 20995
rect 30021 20961 30055 20995
rect 31033 20961 31067 20995
rect 14933 20893 14967 20927
rect 18521 20893 18555 20927
rect 21189 20893 21223 20927
rect 28273 20893 28307 20927
rect 29009 20893 29043 20927
rect 29837 20893 29871 20927
rect 30941 20893 30975 20927
rect 31769 20893 31803 20927
rect 37473 20893 37507 20927
rect 37749 20893 37783 20927
rect 1685 20825 1719 20859
rect 15209 20825 15243 20859
rect 19717 20825 19751 20859
rect 19809 20825 19843 20859
rect 25973 20825 26007 20859
rect 26893 20825 26927 20859
rect 30481 20825 30515 20859
rect 1777 20757 1811 20791
rect 10885 20757 10919 20791
rect 18613 20757 18647 20791
rect 31585 20757 31619 20791
rect 22109 20553 22143 20587
rect 25789 20553 25823 20587
rect 27997 20553 28031 20587
rect 30481 20553 30515 20587
rect 8217 20485 8251 20519
rect 9045 20485 9079 20519
rect 13737 20485 13771 20519
rect 1777 20417 1811 20451
rect 11713 20417 11747 20451
rect 20361 20417 20395 20451
rect 22017 20417 22051 20451
rect 25697 20417 25731 20451
rect 27261 20417 27295 20451
rect 27897 20417 27931 20451
rect 28641 20417 28675 20451
rect 30665 20417 30699 20451
rect 31309 20417 31343 20451
rect 31769 20417 31803 20451
rect 2697 20349 2731 20383
rect 2973 20349 3007 20383
rect 12449 20349 12483 20383
rect 14565 20349 14599 20383
rect 20637 20349 20671 20383
rect 31125 20349 31159 20383
rect 28825 20281 28859 20315
rect 1593 20213 1627 20247
rect 4445 20213 4479 20247
rect 27353 20213 27387 20247
rect 3433 19941 3467 19975
rect 1961 19873 1995 19907
rect 5917 19873 5951 19907
rect 11621 19873 11655 19907
rect 13369 19873 13403 19907
rect 20545 19873 20579 19907
rect 27445 19873 27479 19907
rect 27813 19873 27847 19907
rect 31309 19873 31343 19907
rect 1685 19805 1719 19839
rect 9321 19805 9355 19839
rect 15117 19805 15151 19839
rect 22109 19805 22143 19839
rect 6193 19737 6227 19771
rect 9597 19737 9631 19771
rect 11897 19737 11931 19771
rect 15393 19737 15427 19771
rect 20637 19737 20671 19771
rect 21557 19737 21591 19771
rect 22569 19737 22603 19771
rect 27537 19737 27571 19771
rect 7665 19669 7699 19703
rect 11069 19669 11103 19703
rect 16865 19669 16899 19703
rect 3341 19465 3375 19499
rect 11161 19465 11195 19499
rect 11805 19465 11839 19499
rect 23673 19465 23707 19499
rect 30941 19465 30975 19499
rect 38117 19465 38151 19499
rect 9689 19397 9723 19431
rect 22201 19397 22235 19431
rect 4261 19329 4295 19363
rect 6561 19329 6595 19363
rect 9413 19329 9447 19363
rect 11713 19329 11747 19363
rect 14565 19329 14599 19363
rect 19901 19329 19935 19363
rect 23581 19329 23615 19363
rect 30849 19329 30883 19363
rect 32597 19329 32631 19363
rect 32689 19329 32723 19363
rect 38301 19329 38335 19363
rect 1593 19261 1627 19295
rect 1869 19261 1903 19295
rect 4537 19261 4571 19295
rect 14841 19261 14875 19295
rect 22109 19261 22143 19295
rect 22385 19261 22419 19295
rect 6009 19125 6043 19159
rect 6824 19125 6858 19159
rect 8309 19125 8343 19159
rect 16313 19125 16347 19159
rect 19993 19125 20027 19159
rect 6193 18921 6227 18955
rect 22293 18921 22327 18955
rect 8585 18853 8619 18887
rect 23029 18853 23063 18887
rect 1869 18785 1903 18819
rect 3341 18785 3375 18819
rect 6837 18785 6871 18819
rect 11989 18785 12023 18819
rect 12265 18785 12299 18819
rect 1593 18717 1627 18751
rect 4445 18717 4479 18751
rect 9597 18717 9631 18751
rect 15393 18717 15427 18751
rect 17417 18717 17451 18751
rect 22201 18717 22235 18751
rect 22937 18717 22971 18751
rect 30297 18717 30331 18751
rect 4721 18649 4755 18683
rect 7113 18649 7147 18683
rect 9873 18649 9907 18683
rect 15669 18649 15703 18683
rect 19533 18649 19567 18683
rect 19625 18649 19659 18683
rect 20545 18649 20579 18683
rect 21097 18649 21131 18683
rect 11345 18581 11379 18615
rect 13737 18581 13771 18615
rect 21189 18581 21223 18615
rect 30389 18581 30423 18615
rect 9965 18377 9999 18411
rect 29745 18377 29779 18411
rect 33149 18377 33183 18411
rect 1685 18309 1719 18343
rect 19901 18309 19935 18343
rect 19993 18309 20027 18343
rect 23857 18309 23891 18343
rect 8217 18241 8251 18275
rect 16865 18241 16899 18275
rect 29653 18241 29687 18275
rect 33333 18241 33367 18275
rect 38025 18241 38059 18275
rect 2605 18173 2639 18207
rect 2881 18173 2915 18207
rect 4629 18173 4663 18207
rect 8493 18173 8527 18207
rect 12909 18173 12943 18207
rect 13185 18173 13219 18207
rect 14933 18173 14967 18207
rect 17141 18173 17175 18207
rect 18613 18173 18647 18207
rect 20269 18173 20303 18207
rect 23765 18173 23799 18207
rect 24041 18173 24075 18207
rect 1777 18037 1811 18071
rect 38209 18037 38243 18071
rect 9229 17833 9263 17867
rect 10333 17833 10367 17867
rect 11516 17833 11550 17867
rect 1593 17697 1627 17731
rect 6101 17697 6135 17731
rect 11253 17697 11287 17731
rect 15117 17697 15151 17731
rect 15393 17697 15427 17731
rect 19809 17697 19843 17731
rect 20821 17697 20855 17731
rect 9137 17629 9171 17663
rect 10241 17629 10275 17663
rect 21557 17629 21591 17663
rect 24593 17629 24627 17663
rect 25513 17629 25547 17663
rect 26341 17629 26375 17663
rect 27813 17629 27847 17663
rect 29009 17629 29043 17663
rect 30205 17629 30239 17663
rect 1869 17561 1903 17595
rect 6377 17561 6411 17595
rect 17141 17561 17175 17595
rect 19901 17561 19935 17595
rect 21649 17561 21683 17595
rect 22293 17561 22327 17595
rect 22385 17561 22419 17595
rect 23305 17561 23339 17595
rect 30389 17561 30423 17595
rect 3341 17493 3375 17527
rect 7849 17493 7883 17527
rect 13001 17493 13035 17527
rect 24685 17493 24719 17527
rect 25329 17493 25363 17527
rect 26157 17493 26191 17527
rect 27905 17493 27939 17527
rect 29101 17493 29135 17527
rect 16957 17289 16991 17323
rect 21005 17289 21039 17323
rect 29929 17221 29963 17255
rect 30849 17221 30883 17255
rect 1685 17153 1719 17187
rect 2513 17153 2547 17187
rect 14105 17153 14139 17187
rect 14197 17153 14231 17187
rect 16865 17153 16899 17187
rect 17785 17153 17819 17187
rect 20913 17153 20947 17187
rect 24685 17153 24719 17187
rect 27353 17153 27387 17187
rect 28089 17153 28123 17187
rect 25329 17085 25363 17119
rect 25973 17085 26007 17119
rect 26157 17085 26191 17119
rect 27905 17085 27939 17119
rect 29837 17085 29871 17119
rect 1869 17017 1903 17051
rect 2329 16949 2363 16983
rect 17877 16949 17911 16983
rect 24777 16949 24811 16983
rect 26341 16949 26375 16983
rect 27169 16949 27203 16983
rect 28549 16949 28583 16983
rect 2789 16745 2823 16779
rect 9781 16677 9815 16711
rect 1961 16609 1995 16643
rect 2329 16609 2363 16643
rect 22385 16609 22419 16643
rect 29929 16609 29963 16643
rect 2881 16541 2915 16575
rect 4169 16541 4203 16575
rect 5549 16541 5583 16575
rect 6745 16541 6779 16575
rect 7389 16541 7423 16575
rect 7481 16541 7515 16575
rect 8125 16541 8159 16575
rect 10885 16541 10919 16575
rect 11529 16541 11563 16575
rect 12173 16541 12207 16575
rect 12265 16541 12299 16575
rect 13553 16541 13587 16575
rect 14289 16541 14323 16575
rect 14381 16541 14415 16575
rect 20085 16541 20119 16575
rect 21189 16541 21223 16575
rect 22569 16541 22603 16575
rect 23489 16541 23523 16575
rect 24593 16541 24627 16575
rect 25421 16541 25455 16575
rect 26249 16541 26283 16575
rect 27813 16541 27847 16575
rect 29745 16541 29779 16575
rect 30389 16541 30423 16575
rect 38025 16541 38059 16575
rect 2237 16473 2271 16507
rect 6837 16473 6871 16507
rect 8217 16473 8251 16507
rect 9229 16473 9263 16507
rect 9330 16473 9364 16507
rect 11621 16473 11655 16507
rect 20177 16473 20211 16507
rect 23029 16473 23063 16507
rect 2973 16405 3007 16439
rect 3985 16405 4019 16439
rect 5641 16405 5675 16439
rect 10977 16405 11011 16439
rect 13645 16405 13679 16439
rect 21281 16405 21315 16439
rect 23581 16405 23615 16439
rect 24685 16405 24719 16439
rect 25237 16405 25271 16439
rect 26065 16405 26099 16439
rect 27905 16405 27939 16439
rect 38209 16405 38243 16439
rect 5273 16201 5307 16235
rect 5917 16201 5951 16235
rect 7757 16201 7791 16235
rect 10425 16201 10459 16235
rect 16957 16201 16991 16235
rect 23121 16201 23155 16235
rect 25605 16201 25639 16235
rect 30113 16201 30147 16235
rect 3065 16133 3099 16167
rect 4537 16133 4571 16167
rect 7297 16133 7331 16167
rect 9045 16133 9079 16167
rect 18245 16133 18279 16167
rect 19165 16133 19199 16167
rect 27353 16133 27387 16167
rect 1593 16065 1627 16099
rect 4445 16065 4479 16099
rect 5181 16065 5215 16099
rect 5825 16065 5859 16099
rect 6561 16065 6595 16099
rect 7205 16065 7239 16099
rect 7665 16065 7699 16099
rect 8493 16065 8527 16099
rect 9689 16065 9723 16099
rect 10333 16065 10367 16099
rect 16865 16065 16899 16099
rect 20085 16065 20119 16099
rect 23029 16065 23063 16099
rect 25789 16065 25823 16099
rect 29009 16065 29043 16099
rect 30021 16065 30055 16099
rect 38025 16065 38059 16099
rect 2973 15997 3007 16031
rect 3617 15997 3651 16031
rect 8217 15997 8251 16031
rect 9137 15997 9171 16031
rect 18153 15997 18187 16031
rect 20269 15997 20303 16031
rect 27261 15997 27295 16031
rect 27905 15997 27939 16031
rect 28825 15929 28859 15963
rect 1777 15861 1811 15895
rect 6653 15861 6687 15895
rect 9781 15861 9815 15895
rect 20729 15861 20763 15895
rect 38209 15861 38243 15895
rect 3341 15657 3375 15691
rect 4077 15657 4111 15691
rect 4813 15657 4847 15691
rect 6745 15657 6779 15691
rect 7849 15657 7883 15691
rect 9229 15657 9263 15691
rect 10609 15657 10643 15691
rect 14565 15657 14599 15691
rect 15485 15657 15519 15691
rect 16773 15657 16807 15691
rect 18061 15657 18095 15691
rect 23581 15657 23615 15691
rect 5457 15589 5491 15623
rect 2145 15521 2179 15555
rect 2421 15521 2455 15555
rect 6101 15521 6135 15555
rect 12725 15521 12759 15555
rect 16129 15521 16163 15555
rect 20545 15521 20579 15555
rect 27629 15521 27663 15555
rect 3249 15453 3283 15487
rect 3985 15453 4019 15487
rect 4721 15453 4755 15487
rect 5365 15453 5399 15487
rect 6009 15453 6043 15487
rect 6653 15453 6687 15487
rect 7757 15453 7791 15487
rect 8401 15453 8435 15487
rect 9137 15453 9171 15487
rect 10517 15453 10551 15487
rect 11989 15453 12023 15487
rect 14473 15453 14507 15487
rect 15393 15453 15427 15487
rect 16029 15447 16063 15481
rect 16681 15453 16715 15487
rect 17969 15453 18003 15487
rect 23489 15453 23523 15487
rect 2237 15385 2271 15419
rect 12817 15385 12851 15419
rect 13737 15385 13771 15419
rect 19809 15385 19843 15419
rect 20637 15385 20671 15419
rect 21189 15385 21223 15419
rect 27353 15385 27387 15419
rect 27445 15385 27479 15419
rect 8493 15317 8527 15351
rect 12081 15317 12115 15351
rect 19901 15317 19935 15351
rect 4813 15113 4847 15147
rect 17141 15113 17175 15147
rect 24869 15113 24903 15147
rect 26525 15113 26559 15147
rect 27721 15113 27755 15147
rect 35173 15113 35207 15147
rect 1961 15045 1995 15079
rect 4169 15045 4203 15079
rect 6745 15045 6779 15079
rect 7665 15045 7699 15079
rect 8217 15045 8251 15079
rect 8861 15045 8895 15079
rect 11989 15045 12023 15079
rect 13461 15045 13495 15079
rect 15117 15045 15151 15079
rect 20913 15045 20947 15079
rect 23397 15045 23431 15079
rect 23489 15045 23523 15079
rect 24041 15045 24075 15079
rect 4077 14977 4111 15011
rect 4721 14977 4755 15011
rect 5365 14977 5399 15011
rect 8125 14977 8159 15011
rect 8769 14977 8803 15011
rect 9781 14977 9815 15011
rect 13369 14977 13403 15011
rect 17049 14977 17083 15011
rect 18797 14977 18831 15011
rect 18889 14977 18923 15011
rect 24777 14977 24811 15011
rect 26433 14977 26467 15011
rect 27445 14977 27479 15011
rect 29377 14977 29411 15011
rect 29837 14977 29871 15011
rect 35357 14977 35391 15011
rect 38025 14977 38059 15011
rect 1869 14909 1903 14943
rect 2973 14909 3007 14943
rect 3157 14909 3191 14943
rect 6653 14909 6687 14943
rect 11897 14909 11931 14943
rect 12909 14909 12943 14943
rect 14473 14909 14507 14943
rect 14657 14909 14691 14943
rect 20821 14909 20855 14943
rect 29929 14909 29963 14943
rect 2421 14841 2455 14875
rect 21373 14841 21407 14875
rect 3617 14773 3651 14807
rect 5457 14773 5491 14807
rect 9873 14773 9907 14807
rect 29193 14773 29227 14807
rect 37841 14773 37875 14807
rect 5549 14569 5583 14603
rect 3341 14501 3375 14535
rect 9321 14501 9355 14535
rect 2513 14433 2547 14467
rect 4077 14433 4111 14467
rect 7113 14433 7147 14467
rect 9965 14433 9999 14467
rect 10609 14433 10643 14467
rect 14565 14433 14599 14467
rect 16313 14433 16347 14467
rect 19533 14433 19567 14467
rect 23397 14433 23431 14467
rect 23673 14433 23707 14467
rect 24685 14433 24719 14467
rect 30573 14433 30607 14467
rect 3249 14365 3283 14399
rect 3985 14365 4019 14399
rect 4905 14365 4939 14399
rect 5089 14365 5123 14399
rect 7665 14365 7699 14399
rect 9229 14365 9263 14399
rect 13553 14365 13587 14399
rect 20177 14365 20211 14399
rect 29009 14365 29043 14399
rect 31953 14365 31987 14399
rect 38025 14365 38059 14399
rect 2145 14297 2179 14331
rect 2237 14297 2271 14331
rect 6101 14297 6135 14331
rect 6193 14297 6227 14331
rect 10057 14297 10091 14331
rect 11897 14297 11931 14331
rect 11989 14297 12023 14331
rect 12909 14297 12943 14331
rect 14657 14297 14691 14331
rect 15209 14297 15243 14331
rect 16037 14297 16071 14331
rect 16129 14297 16163 14331
rect 19625 14297 19659 14331
rect 23489 14297 23523 14331
rect 24777 14297 24811 14331
rect 25697 14297 25731 14331
rect 30297 14297 30331 14331
rect 30389 14297 30423 14331
rect 7757 14229 7791 14263
rect 13645 14229 13679 14263
rect 28825 14229 28859 14263
rect 31769 14229 31803 14263
rect 38209 14229 38243 14263
rect 2053 14025 2087 14059
rect 2973 14025 3007 14059
rect 5181 14025 5215 14059
rect 6653 14025 6687 14059
rect 21005 14025 21039 14059
rect 24041 14025 24075 14059
rect 30849 14025 30883 14059
rect 3709 13957 3743 13991
rect 4629 13957 4663 13991
rect 7665 13957 7699 13991
rect 9229 13957 9263 13991
rect 10609 13957 10643 13991
rect 11897 13957 11931 13991
rect 13921 13957 13955 13991
rect 17601 13957 17635 13991
rect 18337 13957 18371 13991
rect 19257 13957 19291 13991
rect 19901 13957 19935 13991
rect 25973 13957 26007 13991
rect 26525 13957 26559 13991
rect 28917 13957 28951 13991
rect 1869 13889 1903 13923
rect 2881 13889 2915 13923
rect 5089 13889 5123 13923
rect 6561 13889 6595 13923
rect 14473 13889 14507 13923
rect 16865 13889 16899 13923
rect 17509 13889 17543 13923
rect 20913 13889 20947 13923
rect 22017 13889 22051 13923
rect 23949 13889 23983 13923
rect 28457 13889 28491 13923
rect 30757 13889 30791 13923
rect 3617 13821 3651 13855
rect 7573 13821 7607 13855
rect 7941 13821 7975 13855
rect 9137 13821 9171 13855
rect 9413 13821 9447 13855
rect 10517 13821 10551 13855
rect 11161 13821 11195 13855
rect 11805 13821 11839 13855
rect 12081 13821 12115 13855
rect 13829 13821 13863 13855
rect 16957 13821 16991 13855
rect 18245 13821 18279 13855
rect 19809 13821 19843 13855
rect 20453 13821 20487 13855
rect 25881 13821 25915 13855
rect 28273 13821 28307 13855
rect 22109 13753 22143 13787
rect 2605 13481 2639 13515
rect 3341 13481 3375 13515
rect 4077 13481 4111 13515
rect 4721 13481 4755 13515
rect 5733 13481 5767 13515
rect 8217 13481 8251 13515
rect 10793 13481 10827 13515
rect 22109 13481 22143 13515
rect 25973 13481 26007 13515
rect 7573 13413 7607 13447
rect 1869 13345 1903 13379
rect 21465 13345 21499 13379
rect 1685 13277 1719 13311
rect 2513 13277 2547 13311
rect 3249 13277 3283 13311
rect 3985 13277 4019 13311
rect 4629 13277 4663 13311
rect 5641 13277 5675 13311
rect 7481 13277 7515 13311
rect 8125 13277 8159 13311
rect 9505 13277 9539 13311
rect 10701 13277 10735 13311
rect 21373 13277 21407 13311
rect 22017 13277 22051 13311
rect 23397 13277 23431 13311
rect 25881 13277 25915 13311
rect 26525 13277 26559 13311
rect 31401 13277 31435 13311
rect 38025 13277 38059 13311
rect 14749 13209 14783 13243
rect 14841 13209 14875 13243
rect 15761 13209 15795 13243
rect 16313 13209 16347 13243
rect 16405 13209 16439 13243
rect 17325 13209 17359 13243
rect 18245 13209 18279 13243
rect 18337 13209 18371 13243
rect 18889 13209 18923 13243
rect 25237 13209 25271 13243
rect 9321 13141 9355 13175
rect 23489 13141 23523 13175
rect 25329 13141 25363 13175
rect 26617 13141 26651 13175
rect 31493 13141 31527 13175
rect 38209 13141 38243 13175
rect 2881 12937 2915 12971
rect 3525 12937 3559 12971
rect 4169 12937 4203 12971
rect 5089 12937 5123 12971
rect 14841 12937 14875 12971
rect 15577 12937 15611 12971
rect 16865 12937 16899 12971
rect 18889 12937 18923 12971
rect 29193 12937 29227 12971
rect 32321 12937 32355 12971
rect 1777 12869 1811 12903
rect 7205 12869 7239 12903
rect 7757 12869 7791 12903
rect 17785 12869 17819 12903
rect 23765 12869 23799 12903
rect 2789 12801 2823 12835
rect 3433 12801 3467 12835
rect 4077 12801 4111 12835
rect 4997 12801 5031 12835
rect 15025 12801 15059 12835
rect 15485 12801 15519 12835
rect 17049 12801 17083 12835
rect 18797 12801 18831 12835
rect 20361 12801 20395 12835
rect 22109 12801 22143 12835
rect 22753 12801 22787 12835
rect 29101 12801 29135 12835
rect 32505 12801 32539 12835
rect 38301 12801 38335 12835
rect 1685 12733 1719 12767
rect 7113 12733 7147 12767
rect 17693 12733 17727 12767
rect 23673 12733 23707 12767
rect 23949 12733 23983 12767
rect 2237 12665 2271 12699
rect 18245 12665 18279 12699
rect 22845 12665 22879 12699
rect 38117 12665 38151 12699
rect 20453 12597 20487 12631
rect 22201 12597 22235 12631
rect 2421 12393 2455 12427
rect 3065 12393 3099 12427
rect 7021 12393 7055 12427
rect 15945 12393 15979 12427
rect 1777 12325 1811 12359
rect 5641 12325 5675 12359
rect 14933 12325 14967 12359
rect 5089 12257 5123 12291
rect 12541 12257 12575 12291
rect 14381 12257 14415 12291
rect 19993 12257 20027 12291
rect 21005 12257 21039 12291
rect 22661 12257 22695 12291
rect 24685 12257 24719 12291
rect 25329 12257 25363 12291
rect 27169 12257 27203 12291
rect 1593 12189 1627 12223
rect 2329 12189 2363 12223
rect 2973 12189 3007 12223
rect 5549 12189 5583 12223
rect 6929 12189 6963 12223
rect 11621 12189 11655 12223
rect 12449 12189 12483 12223
rect 13093 12189 13127 12223
rect 16129 12189 16163 12223
rect 23765 12189 23799 12223
rect 4077 12121 4111 12155
rect 4169 12121 4203 12155
rect 14473 12121 14507 12155
rect 20085 12121 20119 12155
rect 22753 12121 22787 12155
rect 23305 12121 23339 12155
rect 24777 12121 24811 12155
rect 26525 12121 26559 12155
rect 26617 12121 26651 12155
rect 11713 12053 11747 12087
rect 13185 12053 13219 12087
rect 23857 12053 23891 12087
rect 4353 11849 4387 11883
rect 5641 11849 5675 11883
rect 7941 11849 7975 11883
rect 14105 11849 14139 11883
rect 14749 11849 14783 11883
rect 16865 11849 16899 11883
rect 27537 11849 27571 11883
rect 1961 11781 1995 11815
rect 2697 11781 2731 11815
rect 6745 11781 6779 11815
rect 7297 11781 7331 11815
rect 8769 11781 8803 11815
rect 9689 11781 9723 11815
rect 1869 11713 1903 11747
rect 4537 11713 4571 11747
rect 5549 11713 5583 11747
rect 8125 11713 8159 11747
rect 14013 11713 14047 11747
rect 14657 11713 14691 11747
rect 17049 11713 17083 11747
rect 22017 11713 22051 11747
rect 27445 11713 27479 11747
rect 2605 11645 2639 11679
rect 3709 11645 3743 11679
rect 6653 11645 6687 11679
rect 8677 11645 8711 11679
rect 10701 11645 10735 11679
rect 25605 11645 25639 11679
rect 28181 11645 28215 11679
rect 28365 11645 28399 11679
rect 3157 11577 3191 11611
rect 28549 11577 28583 11611
rect 22109 11509 22143 11543
rect 1685 11305 1719 11339
rect 11897 11305 11931 11339
rect 22661 11305 22695 11339
rect 26433 11305 26467 11339
rect 27445 11305 27479 11339
rect 38117 11305 38151 11339
rect 6653 11237 6687 11271
rect 14933 11237 14967 11271
rect 15945 11237 15979 11271
rect 3341 11169 3375 11203
rect 4813 11169 4847 11203
rect 5181 11169 5215 11203
rect 10701 11169 10735 11203
rect 11161 11169 11195 11203
rect 14381 11169 14415 11203
rect 22017 11169 22051 11203
rect 22201 11169 22235 11203
rect 24685 11169 24719 11203
rect 25789 11169 25823 11203
rect 28181 11169 28215 11203
rect 1593 11101 1627 11135
rect 6561 11101 6595 11135
rect 7205 11101 7239 11135
rect 8585 11101 8619 11135
rect 9321 11101 9355 11135
rect 9965 11101 9999 11135
rect 10057 11101 10091 11135
rect 11805 11101 11839 11135
rect 15761 11101 15795 11135
rect 25973 11101 26007 11135
rect 27353 11101 27387 11135
rect 38301 11101 38335 11135
rect 2329 11033 2363 11067
rect 2421 11033 2455 11067
rect 4905 11033 4939 11067
rect 7297 11033 7331 11067
rect 7941 11033 7975 11067
rect 8033 11033 8067 11067
rect 9413 11033 9447 11067
rect 10793 11033 10827 11067
rect 14473 11033 14507 11067
rect 17233 11033 17267 11067
rect 17325 11033 17359 11067
rect 18245 11033 18279 11067
rect 20545 11033 20579 11067
rect 20637 11033 20671 11067
rect 21557 11033 21591 11067
rect 24777 11033 24811 11067
rect 25329 11033 25363 11067
rect 2881 10761 2915 10795
rect 4445 10761 4479 10795
rect 5089 10761 5123 10795
rect 14657 10761 14691 10795
rect 17693 10761 17727 10795
rect 23305 10761 23339 10795
rect 23949 10761 23983 10795
rect 27353 10761 27387 10795
rect 28181 10761 28215 10795
rect 1869 10693 1903 10727
rect 3617 10693 3651 10727
rect 6653 10693 6687 10727
rect 15301 10693 15335 10727
rect 19165 10693 19199 10727
rect 26065 10693 26099 10727
rect 3525 10625 3559 10659
rect 4353 10625 4387 10659
rect 4997 10625 5031 10659
rect 5641 10625 5675 10659
rect 6561 10625 6595 10659
rect 11713 10625 11747 10659
rect 14565 10625 14599 10659
rect 15209 10625 15243 10659
rect 17601 10625 17635 10659
rect 18429 10625 18463 10659
rect 20729 10625 20763 10659
rect 22017 10625 22051 10659
rect 22661 10625 22695 10659
rect 23489 10625 23523 10659
rect 24133 10625 24167 10659
rect 24777 10625 24811 10659
rect 25421 10625 25455 10659
rect 27537 10625 27571 10659
rect 28365 10625 28399 10659
rect 1777 10557 1811 10591
rect 2421 10557 2455 10591
rect 19073 10557 19107 10591
rect 19441 10557 19475 10591
rect 25973 10557 26007 10591
rect 26617 10557 26651 10591
rect 24593 10489 24627 10523
rect 5733 10421 5767 10455
rect 11805 10421 11839 10455
rect 18245 10421 18279 10455
rect 20821 10421 20855 10455
rect 22109 10421 22143 10455
rect 22753 10421 22787 10455
rect 25237 10421 25271 10455
rect 2145 10217 2179 10251
rect 2789 10217 2823 10251
rect 18245 10217 18279 10251
rect 20085 10217 20119 10251
rect 23673 10217 23707 10251
rect 25237 10217 25271 10251
rect 14749 10081 14783 10115
rect 16221 10081 16255 10115
rect 17785 10081 17819 10115
rect 19441 10081 19475 10115
rect 19625 10081 19659 10115
rect 22477 10081 22511 10115
rect 37749 10081 37783 10115
rect 2053 10013 2087 10047
rect 2697 10013 2731 10047
rect 4169 10013 4203 10047
rect 5825 10013 5859 10047
rect 17601 10013 17635 10047
rect 18889 10013 18923 10047
rect 21373 10013 21407 10047
rect 23857 10013 23891 10047
rect 25421 10013 25455 10047
rect 37473 10013 37507 10047
rect 14841 9945 14875 9979
rect 15761 9945 15795 9979
rect 22569 9945 22603 9979
rect 23121 9945 23155 9979
rect 3985 9877 4019 9911
rect 5917 9877 5951 9911
rect 18705 9877 18739 9911
rect 21465 9877 21499 9911
rect 25881 9877 25915 9911
rect 1777 9673 1811 9707
rect 18705 9673 18739 9707
rect 2421 9605 2455 9639
rect 3157 9605 3191 9639
rect 3801 9605 3835 9639
rect 17049 9605 17083 9639
rect 17141 9605 17175 9639
rect 17693 9605 17727 9639
rect 19533 9605 19567 9639
rect 20729 9605 20763 9639
rect 30297 9605 30331 9639
rect 1685 9537 1719 9571
rect 2329 9537 2363 9571
rect 3065 9537 3099 9571
rect 3709 9537 3743 9571
rect 7113 9537 7147 9571
rect 14197 9537 14231 9571
rect 18613 9537 18647 9571
rect 20085 9537 20119 9571
rect 25237 9537 25271 9571
rect 25697 9537 25731 9571
rect 26341 9537 26375 9571
rect 27169 9537 27203 9571
rect 30205 9537 30239 9571
rect 7205 9469 7239 9503
rect 15301 9469 15335 9503
rect 15485 9469 15519 9503
rect 19441 9469 19475 9503
rect 20637 9469 20671 9503
rect 21281 9469 21315 9503
rect 25881 9469 25915 9503
rect 27353 9469 27387 9503
rect 14289 9333 14323 9367
rect 15945 9333 15979 9367
rect 25053 9333 25087 9367
rect 27537 9333 27571 9367
rect 2605 9129 2639 9163
rect 17877 9129 17911 9163
rect 19809 9129 19843 9163
rect 25973 9129 26007 9163
rect 26525 9129 26559 9163
rect 2053 9061 2087 9095
rect 3249 9061 3283 9095
rect 14657 9061 14691 9095
rect 11529 8993 11563 9027
rect 14289 8993 14323 9027
rect 15945 8993 15979 9027
rect 18797 8993 18831 9027
rect 19625 8993 19659 9027
rect 23121 8993 23155 9027
rect 23489 8993 23523 9027
rect 2513 8925 2547 8959
rect 3157 8925 3191 8959
rect 14473 8925 14507 8959
rect 17785 8925 17819 8959
rect 18705 8925 18739 8959
rect 19441 8925 19475 8959
rect 22385 8925 22419 8959
rect 25881 8925 25915 8959
rect 26709 8925 26743 8959
rect 36001 8925 36035 8959
rect 1869 8857 1903 8891
rect 11253 8857 11287 8891
rect 11345 8857 11379 8891
rect 15761 8857 15795 8891
rect 23213 8857 23247 8891
rect 22477 8789 22511 8823
rect 36093 8789 36127 8823
rect 1777 8585 1811 8619
rect 15393 8585 15427 8619
rect 27261 8585 27295 8619
rect 38117 8585 38151 8619
rect 2421 8517 2455 8551
rect 1593 8449 1627 8483
rect 2329 8449 2363 8483
rect 12081 8449 12115 8483
rect 13185 8449 13219 8483
rect 14657 8449 14691 8483
rect 15577 8449 15611 8483
rect 16221 8449 16255 8483
rect 20545 8449 20579 8483
rect 27169 8449 27203 8483
rect 36461 8449 36495 8483
rect 38301 8449 38335 8483
rect 3065 8381 3099 8415
rect 12265 8381 12299 8415
rect 13277 8381 13311 8415
rect 14749 8313 14783 8347
rect 16037 8313 16071 8347
rect 20361 8313 20395 8347
rect 36277 8313 36311 8347
rect 12449 8245 12483 8279
rect 19533 8041 19567 8075
rect 15301 7973 15335 8007
rect 2145 7905 2179 7939
rect 3157 7905 3191 7939
rect 12541 7905 12575 7939
rect 14749 7905 14783 7939
rect 25881 7905 25915 7939
rect 27445 7905 27479 7939
rect 3985 7837 4019 7871
rect 10241 7837 10275 7871
rect 11897 7837 11931 7871
rect 12081 7837 12115 7871
rect 16589 7837 16623 7871
rect 19441 7837 19475 7871
rect 23489 7837 23523 7871
rect 27353 7837 27387 7871
rect 38301 7837 38335 7871
rect 2237 7769 2271 7803
rect 14841 7769 14875 7803
rect 21557 7769 21591 7803
rect 21649 7769 21683 7803
rect 22569 7769 22603 7803
rect 25973 7769 26007 7803
rect 26893 7769 26927 7803
rect 4077 7701 4111 7735
rect 10333 7701 10367 7735
rect 13001 7701 13035 7735
rect 16405 7701 16439 7735
rect 23581 7701 23615 7735
rect 38117 7701 38151 7735
rect 1593 7497 1627 7531
rect 13553 7497 13587 7531
rect 14749 7497 14783 7531
rect 22109 7497 22143 7531
rect 2973 7429 3007 7463
rect 3065 7429 3099 7463
rect 3985 7429 4019 7463
rect 11897 7429 11931 7463
rect 18337 7429 18371 7463
rect 19257 7429 19291 7463
rect 19901 7429 19935 7463
rect 23121 7429 23155 7463
rect 1777 7361 1811 7395
rect 2237 7361 2271 7395
rect 6561 7361 6595 7395
rect 11161 7361 11195 7395
rect 12909 7361 12943 7395
rect 14657 7361 14691 7395
rect 22017 7361 22051 7395
rect 11805 7293 11839 7327
rect 12173 7293 12207 7327
rect 13093 7293 13127 7327
rect 17417 7293 17451 7327
rect 18245 7293 18279 7327
rect 19809 7293 19843 7327
rect 20085 7293 20119 7327
rect 23029 7293 23063 7327
rect 23581 7225 23615 7259
rect 2329 7157 2363 7191
rect 6653 7157 6687 7191
rect 10977 7157 11011 7191
rect 11529 6953 11563 6987
rect 23489 6953 23523 6987
rect 12449 6817 12483 6851
rect 17325 6817 17359 6851
rect 17969 6817 18003 6851
rect 1777 6749 1811 6783
rect 3249 6749 3283 6783
rect 6837 6749 6871 6783
rect 11713 6749 11747 6783
rect 12357 6749 12391 6783
rect 15393 6749 15427 6783
rect 15577 6749 15611 6783
rect 17509 6749 17543 6783
rect 19809 6749 19843 6783
rect 23029 6749 23063 6783
rect 23673 6749 23707 6783
rect 16037 6681 16071 6715
rect 1593 6613 1627 6647
rect 3065 6613 3099 6647
rect 6653 6613 6687 6647
rect 19901 6613 19935 6647
rect 22845 6613 22879 6647
rect 1961 6409 1995 6443
rect 11897 6409 11931 6443
rect 13185 6409 13219 6443
rect 13829 6409 13863 6443
rect 15669 6409 15703 6443
rect 17601 6409 17635 6443
rect 18521 6409 18555 6443
rect 25973 6409 26007 6443
rect 1869 6341 1903 6375
rect 6745 6273 6779 6307
rect 11805 6273 11839 6307
rect 13369 6273 13403 6307
rect 14013 6273 14047 6307
rect 15577 6273 15611 6307
rect 17509 6273 17543 6307
rect 18429 6273 18463 6307
rect 25237 6273 25271 6307
rect 25881 6273 25915 6307
rect 38301 6273 38335 6307
rect 6561 6069 6595 6103
rect 25329 6069 25363 6103
rect 38117 6069 38151 6103
rect 14381 5865 14415 5899
rect 27721 5865 27755 5899
rect 2053 5797 2087 5831
rect 2513 5661 2547 5695
rect 14289 5661 14323 5695
rect 25697 5661 25731 5695
rect 27629 5661 27663 5695
rect 1869 5593 1903 5627
rect 2605 5593 2639 5627
rect 25513 5525 25547 5559
rect 1593 5321 1627 5355
rect 17785 5253 17819 5287
rect 1777 5185 1811 5219
rect 29929 5185 29963 5219
rect 38025 5185 38059 5219
rect 17693 5117 17727 5151
rect 18705 5117 18739 5151
rect 30021 4981 30055 5015
rect 38209 4981 38243 5015
rect 38117 4777 38151 4811
rect 1593 4573 1627 4607
rect 38301 4573 38335 4607
rect 1777 4437 1811 4471
rect 38117 4165 38151 4199
rect 1777 4097 1811 4131
rect 6837 4097 6871 4131
rect 18613 4097 18647 4131
rect 20545 4097 20579 4131
rect 36369 4097 36403 4131
rect 18705 4029 18739 4063
rect 1593 3961 1627 3995
rect 38301 3961 38335 3995
rect 6929 3893 6963 3927
rect 20637 3893 20671 3927
rect 36185 3893 36219 3927
rect 1869 3485 1903 3519
rect 2237 3485 2271 3519
rect 21925 3485 21959 3519
rect 32781 3485 32815 3519
rect 38025 3485 38059 3519
rect 37381 3417 37415 3451
rect 1685 3349 1719 3383
rect 21741 3349 21775 3383
rect 32597 3349 32631 3383
rect 37473 3349 37507 3383
rect 38209 3349 38243 3383
rect 3065 3145 3099 3179
rect 9781 3145 9815 3179
rect 36829 3145 36863 3179
rect 1593 3009 1627 3043
rect 2329 3009 2363 3043
rect 3249 3009 3283 3043
rect 6745 3009 6779 3043
rect 9965 3009 9999 3043
rect 13185 3009 13219 3043
rect 14381 3009 14415 3043
rect 17233 3009 17267 3043
rect 36737 3009 36771 3043
rect 37473 2941 37507 2975
rect 37749 2941 37783 2975
rect 2513 2873 2547 2907
rect 14565 2873 14599 2907
rect 1777 2805 1811 2839
rect 6561 2805 6595 2839
rect 13001 2805 13035 2839
rect 17049 2805 17083 2839
rect 7297 2601 7331 2635
rect 11713 2601 11747 2635
rect 13001 2601 13035 2635
rect 16865 2601 16899 2635
rect 17509 2601 17543 2635
rect 19441 2601 19475 2635
rect 20729 2601 20763 2635
rect 22017 2601 22051 2635
rect 24593 2601 24627 2635
rect 27169 2601 27203 2635
rect 28457 2601 28491 2635
rect 32321 2601 32355 2635
rect 10977 2533 11011 2567
rect 30481 2533 30515 2567
rect 33241 2533 33275 2567
rect 4261 2465 4295 2499
rect 9413 2465 9447 2499
rect 37749 2465 37783 2499
rect 2053 2397 2087 2431
rect 2881 2397 2915 2431
rect 3433 2397 3467 2431
rect 3985 2397 4019 2431
rect 5273 2397 5307 2431
rect 6561 2397 6595 2431
rect 7481 2397 7515 2431
rect 9137 2397 9171 2431
rect 11161 2397 11195 2431
rect 11897 2397 11931 2431
rect 13185 2397 13219 2431
rect 14933 2397 14967 2431
rect 17049 2397 17083 2431
rect 17693 2397 17727 2431
rect 18153 2397 18187 2431
rect 19625 2397 19659 2431
rect 20913 2397 20947 2431
rect 22201 2397 22235 2431
rect 22661 2397 22695 2431
rect 24777 2397 24811 2431
rect 25237 2397 25271 2431
rect 25973 2397 26007 2431
rect 27353 2397 27387 2431
rect 28641 2397 28675 2431
rect 29745 2397 29779 2431
rect 30665 2397 30699 2431
rect 32505 2397 32539 2431
rect 33701 2397 33735 2431
rect 34897 2397 34931 2431
rect 36185 2397 36219 2431
rect 37473 2397 37507 2431
rect 33057 2329 33091 2363
rect 2237 2261 2271 2295
rect 3249 2261 3283 2295
rect 5457 2261 5491 2295
rect 6745 2261 6779 2295
rect 15117 2261 15151 2295
rect 18337 2261 18371 2295
rect 22845 2261 22879 2295
rect 25421 2261 25455 2295
rect 26157 2261 26191 2295
rect 29929 2261 29963 2295
rect 33885 2261 33919 2295
rect 35081 2261 35115 2295
rect 36369 2261 36403 2295
<< metal1 >>
rect 17218 37612 17224 37664
rect 17276 37652 17282 37664
rect 21358 37652 21364 37664
rect 17276 37624 21364 37652
rect 17276 37612 17282 37624
rect 21358 37612 21364 37624
rect 21416 37612 21422 37664
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 5902 37408 5908 37460
rect 5960 37448 5966 37460
rect 24026 37448 24032 37460
rect 5960 37420 24032 37448
rect 5960 37408 5966 37420
rect 24026 37408 24032 37420
rect 24084 37408 24090 37460
rect 3973 37383 4031 37389
rect 3973 37349 3985 37383
rect 4019 37380 4031 37383
rect 6914 37380 6920 37392
rect 4019 37352 6920 37380
rect 4019 37349 4031 37352
rect 3973 37343 4031 37349
rect 6914 37340 6920 37352
rect 6972 37340 6978 37392
rect 8754 37340 8760 37392
rect 8812 37380 8818 37392
rect 17218 37380 17224 37392
rect 8812 37352 17224 37380
rect 8812 37340 8818 37352
rect 17218 37340 17224 37352
rect 17276 37340 17282 37392
rect 17310 37340 17316 37392
rect 17368 37380 17374 37392
rect 19426 37380 19432 37392
rect 17368 37352 19432 37380
rect 17368 37340 17374 37352
rect 19426 37340 19432 37352
rect 19484 37340 19490 37392
rect 21082 37340 21088 37392
rect 21140 37380 21146 37392
rect 25317 37383 25375 37389
rect 25317 37380 25329 37383
rect 21140 37352 25329 37380
rect 21140 37340 21146 37352
rect 25317 37349 25329 37352
rect 25363 37349 25375 37383
rect 25317 37343 25375 37349
rect 1578 37312 1584 37324
rect 1539 37284 1584 37312
rect 1578 37272 1584 37284
rect 1636 37272 1642 37324
rect 11974 37312 11980 37324
rect 8220 37284 8524 37312
rect 1857 37247 1915 37253
rect 1857 37213 1869 37247
rect 1903 37213 1915 37247
rect 2866 37244 2872 37256
rect 2827 37216 2872 37244
rect 1857 37207 1915 37213
rect 1872 37176 1900 37207
rect 2866 37204 2872 37216
rect 2924 37204 2930 37256
rect 3234 37204 3240 37256
rect 3292 37244 3298 37256
rect 4157 37247 4215 37253
rect 4157 37244 4169 37247
rect 3292 37216 4169 37244
rect 3292 37204 3298 37216
rect 4157 37213 4169 37216
rect 4203 37213 4215 37247
rect 4157 37207 4215 37213
rect 4614 37204 4620 37256
rect 4672 37244 4678 37256
rect 4801 37247 4859 37253
rect 4801 37244 4813 37247
rect 4672 37216 4813 37244
rect 4672 37204 4678 37216
rect 4801 37213 4813 37216
rect 4847 37213 4859 37247
rect 4801 37207 4859 37213
rect 5810 37204 5816 37256
rect 5868 37244 5874 37256
rect 5997 37247 6055 37253
rect 5997 37244 6009 37247
rect 5868 37216 6009 37244
rect 5868 37204 5874 37216
rect 5997 37213 6009 37216
rect 6043 37213 6055 37247
rect 5997 37207 6055 37213
rect 6454 37204 6460 37256
rect 6512 37244 6518 37256
rect 6733 37247 6791 37253
rect 6733 37244 6745 37247
rect 6512 37216 6745 37244
rect 6512 37204 6518 37216
rect 6733 37213 6745 37216
rect 6779 37213 6791 37247
rect 6733 37207 6791 37213
rect 7561 37247 7619 37253
rect 7561 37213 7573 37247
rect 7607 37244 7619 37247
rect 8220 37244 8248 37284
rect 7607 37216 8248 37244
rect 8297 37247 8355 37253
rect 7607 37213 7619 37216
rect 7561 37207 7619 37213
rect 8297 37213 8309 37247
rect 8343 37244 8355 37247
rect 8386 37244 8392 37256
rect 8343 37216 8392 37244
rect 8343 37213 8355 37216
rect 8297 37207 8355 37213
rect 8386 37204 8392 37216
rect 8444 37204 8450 37256
rect 8496 37244 8524 37284
rect 9692 37284 10088 37312
rect 11935 37284 11980 37312
rect 9692 37244 9720 37284
rect 10060 37256 10088 37284
rect 11974 37272 11980 37284
rect 12032 37272 12038 37324
rect 22005 37315 22063 37321
rect 22005 37312 22017 37315
rect 14292 37284 21220 37312
rect 8496 37216 9720 37244
rect 9769 37247 9827 37253
rect 9769 37213 9781 37247
rect 9815 37244 9827 37247
rect 9950 37244 9956 37256
rect 9815 37216 9956 37244
rect 9815 37213 9827 37216
rect 9769 37207 9827 37213
rect 9950 37204 9956 37216
rect 10008 37204 10014 37256
rect 10042 37204 10048 37256
rect 10100 37204 10106 37256
rect 11149 37247 11207 37253
rect 11149 37213 11161 37247
rect 11195 37244 11207 37247
rect 12250 37244 12256 37256
rect 11195 37216 12256 37244
rect 11195 37213 11207 37216
rect 11149 37207 11207 37213
rect 12250 37204 12256 37216
rect 12308 37204 12314 37256
rect 13081 37247 13139 37253
rect 13081 37213 13093 37247
rect 13127 37213 13139 37247
rect 13081 37207 13139 37213
rect 13725 37247 13783 37253
rect 13725 37213 13737 37247
rect 13771 37244 13783 37247
rect 14090 37244 14096 37256
rect 13771 37216 14096 37244
rect 13771 37213 13783 37216
rect 13725 37207 13783 37213
rect 4706 37176 4712 37188
rect 1872 37148 4712 37176
rect 4706 37136 4712 37148
rect 4764 37136 4770 37188
rect 10870 37176 10876 37188
rect 5828 37148 10876 37176
rect 2774 37068 2780 37120
rect 2832 37108 2838 37120
rect 3053 37111 3111 37117
rect 3053 37108 3065 37111
rect 2832 37080 3065 37108
rect 2832 37068 2838 37080
rect 3053 37077 3065 37080
rect 3099 37077 3111 37111
rect 3053 37071 3111 37077
rect 4614 37068 4620 37120
rect 4672 37108 4678 37120
rect 5828 37117 5856 37148
rect 10870 37136 10876 37148
rect 10928 37136 10934 37188
rect 11054 37136 11060 37188
rect 11112 37176 11118 37188
rect 11793 37179 11851 37185
rect 11793 37176 11805 37179
rect 11112 37148 11805 37176
rect 11112 37136 11118 37148
rect 11793 37145 11805 37148
rect 11839 37145 11851 37179
rect 13096 37176 13124 37207
rect 14090 37204 14096 37216
rect 14148 37204 14154 37256
rect 14292 37253 14320 37284
rect 14277 37247 14335 37253
rect 14277 37213 14289 37247
rect 14323 37213 14335 37247
rect 14277 37207 14335 37213
rect 15194 37204 15200 37256
rect 15252 37244 15258 37256
rect 15381 37247 15439 37253
rect 15381 37244 15393 37247
rect 15252 37216 15393 37244
rect 15252 37204 15258 37216
rect 15381 37213 15393 37216
rect 15427 37213 15439 37247
rect 15381 37207 15439 37213
rect 15470 37204 15476 37256
rect 15528 37204 15534 37256
rect 16025 37247 16083 37253
rect 16025 37213 16037 37247
rect 16071 37213 16083 37247
rect 16025 37207 16083 37213
rect 15488 37176 15516 37204
rect 13096 37148 15516 37176
rect 16040 37176 16068 37207
rect 16850 37204 16856 37256
rect 16908 37244 16914 37256
rect 17310 37244 17316 37256
rect 16908 37216 17316 37244
rect 16908 37204 16914 37216
rect 17310 37204 17316 37216
rect 17368 37204 17374 37256
rect 17494 37244 17500 37256
rect 17455 37216 17500 37244
rect 17494 37204 17500 37216
rect 17552 37204 17558 37256
rect 18598 37204 18604 37256
rect 18656 37244 18662 37256
rect 18693 37247 18751 37253
rect 18693 37244 18705 37247
rect 18656 37216 18705 37244
rect 18656 37204 18662 37216
rect 18693 37213 18705 37216
rect 18739 37213 18751 37247
rect 18693 37207 18751 37213
rect 18782 37204 18788 37256
rect 18840 37244 18846 37256
rect 18840 37216 18885 37244
rect 18840 37204 18846 37216
rect 19426 37204 19432 37256
rect 19484 37244 19490 37256
rect 20070 37244 20076 37256
rect 19484 37216 19529 37244
rect 20031 37216 20076 37244
rect 19484 37204 19490 37216
rect 20070 37204 20076 37216
rect 20128 37204 20134 37256
rect 21082 37176 21088 37188
rect 16040 37148 18644 37176
rect 11793 37139 11851 37145
rect 5813 37111 5871 37117
rect 4672 37080 4717 37108
rect 4672 37068 4678 37080
rect 5813 37077 5825 37111
rect 5859 37077 5871 37111
rect 6546 37108 6552 37120
rect 6507 37080 6552 37108
rect 5813 37071 5871 37077
rect 6546 37068 6552 37080
rect 6604 37068 6610 37120
rect 7742 37108 7748 37120
rect 7703 37080 7748 37108
rect 7742 37068 7748 37080
rect 7800 37068 7806 37120
rect 8481 37111 8539 37117
rect 8481 37077 8493 37111
rect 8527 37108 8539 37111
rect 9030 37108 9036 37120
rect 8527 37080 9036 37108
rect 8527 37077 8539 37080
rect 8481 37071 8539 37077
rect 9030 37068 9036 37080
rect 9088 37068 9094 37120
rect 9674 37068 9680 37120
rect 9732 37108 9738 37120
rect 9953 37111 10011 37117
rect 9953 37108 9965 37111
rect 9732 37080 9965 37108
rect 9732 37068 9738 37080
rect 9953 37077 9965 37080
rect 9999 37077 10011 37111
rect 9953 37071 10011 37077
rect 10965 37111 11023 37117
rect 10965 37077 10977 37111
rect 11011 37108 11023 37111
rect 12802 37108 12808 37120
rect 11011 37080 12808 37108
rect 11011 37077 11023 37080
rect 10965 37071 11023 37077
rect 12802 37068 12808 37080
rect 12860 37068 12866 37120
rect 12897 37111 12955 37117
rect 12897 37077 12909 37111
rect 12943 37108 12955 37111
rect 13446 37108 13452 37120
rect 12943 37080 13452 37108
rect 12943 37077 12955 37080
rect 12897 37071 12955 37077
rect 13446 37068 13452 37080
rect 13504 37068 13510 37120
rect 13541 37111 13599 37117
rect 13541 37077 13553 37111
rect 13587 37108 13599 37111
rect 13722 37108 13728 37120
rect 13587 37080 13728 37108
rect 13587 37077 13599 37080
rect 13541 37071 13599 37077
rect 13722 37068 13728 37080
rect 13780 37068 13786 37120
rect 13814 37068 13820 37120
rect 13872 37108 13878 37120
rect 14461 37111 14519 37117
rect 14461 37108 14473 37111
rect 13872 37080 14473 37108
rect 13872 37068 13878 37080
rect 14461 37077 14473 37080
rect 14507 37077 14519 37111
rect 14461 37071 14519 37077
rect 15286 37068 15292 37120
rect 15344 37108 15350 37120
rect 15473 37111 15531 37117
rect 15473 37108 15485 37111
rect 15344 37080 15485 37108
rect 15344 37068 15350 37080
rect 15473 37077 15485 37080
rect 15519 37077 15531 37111
rect 15473 37071 15531 37077
rect 16209 37111 16267 37117
rect 16209 37077 16221 37111
rect 16255 37108 16267 37111
rect 16758 37108 16764 37120
rect 16255 37080 16764 37108
rect 16255 37077 16267 37080
rect 16209 37071 16267 37077
rect 16758 37068 16764 37080
rect 16816 37068 16822 37120
rect 16942 37108 16948 37120
rect 16903 37080 16948 37108
rect 16942 37068 16948 37080
rect 17000 37068 17006 37120
rect 17402 37068 17408 37120
rect 17460 37108 17466 37120
rect 17681 37111 17739 37117
rect 17681 37108 17693 37111
rect 17460 37080 17693 37108
rect 17460 37068 17466 37080
rect 17681 37077 17693 37080
rect 17727 37077 17739 37111
rect 18616 37108 18644 37148
rect 18800 37148 21088 37176
rect 18800 37108 18828 37148
rect 21082 37136 21088 37148
rect 21140 37136 21146 37188
rect 18616 37080 18828 37108
rect 17681 37071 17739 37077
rect 19334 37068 19340 37120
rect 19392 37108 19398 37120
rect 19521 37111 19579 37117
rect 19521 37108 19533 37111
rect 19392 37080 19533 37108
rect 19392 37068 19398 37080
rect 19521 37077 19533 37080
rect 19567 37077 19579 37111
rect 19521 37071 19579 37077
rect 19978 37068 19984 37120
rect 20036 37108 20042 37120
rect 21192 37117 21220 37284
rect 21284 37284 22017 37312
rect 21284 37256 21312 37284
rect 22005 37281 22017 37284
rect 22051 37281 22063 37315
rect 22005 37275 22063 37281
rect 23569 37315 23627 37321
rect 23569 37281 23581 37315
rect 23615 37312 23627 37315
rect 23658 37312 23664 37324
rect 23615 37284 23664 37312
rect 23615 37281 23627 37284
rect 23569 37275 23627 37281
rect 23658 37272 23664 37284
rect 23716 37272 23722 37324
rect 25130 37272 25136 37324
rect 25188 37312 25194 37324
rect 25188 37284 26004 37312
rect 25188 37272 25194 37284
rect 21266 37204 21272 37256
rect 21324 37204 21330 37256
rect 21361 37247 21419 37253
rect 21361 37213 21373 37247
rect 21407 37246 21419 37247
rect 21450 37246 21456 37256
rect 21407 37218 21456 37246
rect 21407 37213 21419 37218
rect 21361 37207 21419 37213
rect 21450 37204 21456 37218
rect 21508 37204 21514 37256
rect 22281 37247 22339 37253
rect 22281 37213 22293 37247
rect 22327 37244 22339 37247
rect 22830 37244 22836 37256
rect 22327 37216 22836 37244
rect 22327 37213 22339 37216
rect 22281 37207 22339 37213
rect 22830 37204 22836 37216
rect 22888 37204 22894 37256
rect 23198 37204 23204 37256
rect 23256 37244 23262 37256
rect 23385 37247 23443 37253
rect 23385 37244 23397 37247
rect 23256 37216 23397 37244
rect 23256 37204 23262 37216
rect 23385 37213 23397 37216
rect 23431 37213 23443 37247
rect 23385 37207 23443 37213
rect 23750 37204 23756 37256
rect 23808 37244 23814 37256
rect 24581 37247 24639 37253
rect 24581 37244 24593 37247
rect 23808 37216 24593 37244
rect 23808 37204 23814 37216
rect 24581 37213 24593 37216
rect 24627 37213 24639 37247
rect 24581 37207 24639 37213
rect 25501 37247 25559 37253
rect 25501 37213 25513 37247
rect 25547 37244 25559 37247
rect 25866 37244 25872 37256
rect 25547 37216 25872 37244
rect 25547 37213 25559 37216
rect 25501 37207 25559 37213
rect 25866 37204 25872 37216
rect 25924 37204 25930 37256
rect 25976 37244 26004 37284
rect 27264 37284 27936 37312
rect 27264 37244 27292 37284
rect 25976 37216 27292 37244
rect 27341 37247 27399 37253
rect 27341 37213 27353 37247
rect 27387 37244 27399 37247
rect 27430 37244 27436 37256
rect 27387 37216 27436 37244
rect 27387 37213 27399 37216
rect 27341 37207 27399 37213
rect 27430 37204 27436 37216
rect 27488 37204 27494 37256
rect 27798 37244 27804 37256
rect 27759 37216 27804 37244
rect 27798 37204 27804 37216
rect 27856 37204 27862 37256
rect 27908 37244 27936 37284
rect 28350 37272 28356 37324
rect 28408 37312 28414 37324
rect 28408 37284 29040 37312
rect 28408 37272 28414 37284
rect 28721 37247 28779 37253
rect 28721 37244 28733 37247
rect 27908 37216 28733 37244
rect 28721 37213 28733 37216
rect 28767 37213 28779 37247
rect 29012 37244 29040 37284
rect 29638 37272 29644 37324
rect 29696 37312 29702 37324
rect 29696 37284 30236 37312
rect 29696 37272 29702 37284
rect 29917 37247 29975 37253
rect 29917 37244 29929 37247
rect 29012 37216 29929 37244
rect 28721 37207 28779 37213
rect 29917 37213 29929 37216
rect 29963 37213 29975 37247
rect 30208 37244 30236 37284
rect 34146 37272 34152 37324
rect 34204 37312 34210 37324
rect 34885 37315 34943 37321
rect 34885 37312 34897 37315
rect 34204 37284 34897 37312
rect 34204 37272 34210 37284
rect 34885 37281 34897 37284
rect 34931 37281 34943 37315
rect 34885 37275 34943 37281
rect 37918 37272 37924 37324
rect 37976 37312 37982 37324
rect 38289 37315 38347 37321
rect 38289 37312 38301 37315
rect 37976 37284 38301 37312
rect 37976 37272 37982 37284
rect 38289 37281 38301 37284
rect 38335 37281 38347 37315
rect 38289 37275 38347 37281
rect 30561 37247 30619 37253
rect 30561 37244 30573 37247
rect 30208 37216 30573 37244
rect 29917 37207 29975 37213
rect 30561 37213 30573 37216
rect 30607 37213 30619 37247
rect 30561 37207 30619 37213
rect 30926 37204 30932 37256
rect 30984 37244 30990 37256
rect 31205 37247 31263 37253
rect 31205 37244 31217 37247
rect 30984 37216 31217 37244
rect 30984 37204 30990 37216
rect 31205 37213 31217 37216
rect 31251 37213 31263 37247
rect 31205 37207 31263 37213
rect 32309 37247 32367 37253
rect 32309 37213 32321 37247
rect 32355 37213 32367 37247
rect 32309 37207 32367 37213
rect 32324 37176 32352 37207
rect 32858 37204 32864 37256
rect 32916 37244 32922 37256
rect 33229 37247 33287 37253
rect 33229 37244 33241 37247
rect 32916 37216 33241 37244
rect 32916 37204 32922 37216
rect 33229 37213 33241 37216
rect 33275 37213 33287 37247
rect 33229 37207 33287 37213
rect 35161 37247 35219 37253
rect 35161 37213 35173 37247
rect 35207 37244 35219 37247
rect 36170 37244 36176 37256
rect 35207 37216 35894 37244
rect 36131 37216 36176 37244
rect 35207 37213 35219 37216
rect 35161 37207 35219 37213
rect 27172 37148 32352 37176
rect 35866 37176 35894 37216
rect 36170 37204 36176 37216
rect 36228 37204 36234 37256
rect 38102 37244 38108 37256
rect 38063 37216 38108 37244
rect 38102 37204 38108 37216
rect 38160 37204 38166 37256
rect 36814 37176 36820 37188
rect 35866 37148 36820 37176
rect 20257 37111 20315 37117
rect 20257 37108 20269 37111
rect 20036 37080 20269 37108
rect 20036 37068 20042 37080
rect 20257 37077 20269 37080
rect 20303 37077 20315 37111
rect 20257 37071 20315 37077
rect 21177 37111 21235 37117
rect 21177 37077 21189 37111
rect 21223 37077 21235 37111
rect 21177 37071 21235 37077
rect 21450 37068 21456 37120
rect 21508 37108 21514 37120
rect 21910 37108 21916 37120
rect 21508 37080 21916 37108
rect 21508 37068 21514 37080
rect 21910 37068 21916 37080
rect 21968 37068 21974 37120
rect 22002 37068 22008 37120
rect 22060 37108 22066 37120
rect 24394 37108 24400 37120
rect 22060 37080 24400 37108
rect 22060 37068 22066 37080
rect 24394 37068 24400 37080
rect 24452 37068 24458 37120
rect 24486 37068 24492 37120
rect 24544 37108 24550 37120
rect 24765 37111 24823 37117
rect 24765 37108 24777 37111
rect 24544 37080 24777 37108
rect 24544 37068 24550 37080
rect 24765 37077 24777 37080
rect 24811 37077 24823 37111
rect 24765 37071 24823 37077
rect 25498 37068 25504 37120
rect 25556 37108 25562 37120
rect 27172 37117 27200 37148
rect 36814 37136 36820 37148
rect 36872 37136 36878 37188
rect 25961 37111 26019 37117
rect 25961 37108 25973 37111
rect 25556 37080 25973 37108
rect 25556 37068 25562 37080
rect 25961 37077 25973 37080
rect 26007 37077 26019 37111
rect 25961 37071 26019 37077
rect 27157 37111 27215 37117
rect 27157 37077 27169 37111
rect 27203 37077 27215 37111
rect 27157 37071 27215 37077
rect 27706 37068 27712 37120
rect 27764 37108 27770 37120
rect 27985 37111 28043 37117
rect 27985 37108 27997 37111
rect 27764 37080 27997 37108
rect 27764 37068 27770 37080
rect 27985 37077 27997 37080
rect 28031 37077 28043 37111
rect 28534 37108 28540 37120
rect 28495 37080 28540 37108
rect 27985 37071 28043 37077
rect 28534 37068 28540 37080
rect 28592 37068 28598 37120
rect 28902 37068 28908 37120
rect 28960 37108 28966 37120
rect 29733 37111 29791 37117
rect 29733 37108 29745 37111
rect 28960 37080 29745 37108
rect 28960 37068 28966 37080
rect 29733 37077 29745 37080
rect 29779 37077 29791 37111
rect 29733 37071 29791 37077
rect 29822 37068 29828 37120
rect 29880 37108 29886 37120
rect 30377 37111 30435 37117
rect 30377 37108 30389 37111
rect 29880 37080 30389 37108
rect 29880 37068 29886 37080
rect 30377 37077 30389 37080
rect 30423 37077 30435 37111
rect 31018 37108 31024 37120
rect 30979 37080 31024 37108
rect 30377 37071 30435 37077
rect 31018 37068 31024 37080
rect 31076 37068 31082 37120
rect 32214 37068 32220 37120
rect 32272 37108 32278 37120
rect 32493 37111 32551 37117
rect 32493 37108 32505 37111
rect 32272 37080 32505 37108
rect 32272 37068 32278 37080
rect 32493 37077 32505 37080
rect 32539 37077 32551 37111
rect 33042 37108 33048 37120
rect 33003 37080 33048 37108
rect 32493 37071 32551 37077
rect 33042 37068 33048 37080
rect 33100 37068 33106 37120
rect 35894 37068 35900 37120
rect 35952 37108 35958 37120
rect 36357 37111 36415 37117
rect 36357 37108 36369 37111
rect 35952 37080 36369 37108
rect 35952 37068 35958 37080
rect 36357 37077 36369 37080
rect 36403 37077 36415 37111
rect 36357 37071 36415 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 1762 36904 1768 36916
rect 1723 36876 1768 36904
rect 1762 36864 1768 36876
rect 1820 36864 1826 36916
rect 2317 36907 2375 36913
rect 2317 36873 2329 36907
rect 2363 36873 2375 36907
rect 2317 36867 2375 36873
rect 14 36796 20 36848
rect 72 36836 78 36848
rect 2332 36836 2360 36867
rect 6546 36864 6552 36916
rect 6604 36904 6610 36916
rect 6604 36876 13584 36904
rect 6604 36864 6610 36876
rect 72 36808 1716 36836
rect 2332 36808 4292 36836
rect 72 36796 78 36808
rect 1578 36768 1584 36780
rect 1539 36740 1584 36768
rect 1578 36728 1584 36740
rect 1636 36728 1642 36780
rect 1688 36768 1716 36808
rect 2501 36771 2559 36777
rect 2501 36768 2513 36771
rect 1688 36740 2513 36768
rect 2501 36737 2513 36740
rect 2547 36737 2559 36771
rect 2958 36768 2964 36780
rect 2919 36740 2964 36768
rect 2501 36731 2559 36737
rect 2958 36728 2964 36740
rect 3016 36728 3022 36780
rect 3789 36771 3847 36777
rect 3789 36737 3801 36771
rect 3835 36768 3847 36771
rect 3970 36768 3976 36780
rect 3835 36740 3976 36768
rect 3835 36737 3847 36740
rect 3789 36731 3847 36737
rect 3970 36728 3976 36740
rect 4028 36728 4034 36780
rect 4264 36777 4292 36808
rect 7926 36796 7932 36848
rect 7984 36836 7990 36848
rect 8665 36839 8723 36845
rect 8665 36836 8677 36839
rect 7984 36808 8677 36836
rect 7984 36796 7990 36808
rect 8665 36805 8677 36808
rect 8711 36805 8723 36839
rect 8665 36799 8723 36805
rect 10229 36839 10287 36845
rect 10229 36805 10241 36839
rect 10275 36836 10287 36839
rect 13354 36836 13360 36848
rect 10275 36808 13360 36836
rect 10275 36805 10287 36808
rect 10229 36799 10287 36805
rect 13354 36796 13360 36808
rect 13412 36796 13418 36848
rect 4249 36771 4307 36777
rect 4249 36737 4261 36771
rect 4295 36737 4307 36771
rect 4249 36731 4307 36737
rect 6733 36771 6791 36777
rect 6733 36737 6745 36771
rect 6779 36768 6791 36771
rect 8294 36768 8300 36780
rect 6779 36740 8300 36768
rect 6779 36737 6791 36740
rect 6733 36731 6791 36737
rect 8294 36728 8300 36740
rect 8352 36728 8358 36780
rect 9674 36728 9680 36780
rect 9732 36768 9738 36780
rect 10137 36771 10195 36777
rect 10137 36768 10149 36771
rect 9732 36740 10149 36768
rect 9732 36728 9738 36740
rect 10137 36737 10149 36740
rect 10183 36737 10195 36771
rect 10965 36771 11023 36777
rect 10965 36768 10977 36771
rect 10137 36731 10195 36737
rect 10244 36740 10977 36768
rect 4798 36660 4804 36712
rect 4856 36700 4862 36712
rect 4893 36703 4951 36709
rect 4893 36700 4905 36703
rect 4856 36672 4905 36700
rect 4856 36660 4862 36672
rect 4893 36669 4905 36672
rect 4939 36669 4951 36703
rect 8573 36703 8631 36709
rect 8573 36700 8585 36703
rect 4893 36663 4951 36669
rect 8128 36672 8585 36700
rect 4341 36635 4399 36641
rect 4341 36601 4353 36635
rect 4387 36632 4399 36635
rect 8128 36632 8156 36672
rect 8573 36669 8585 36672
rect 8619 36669 8631 36703
rect 8573 36663 8631 36669
rect 8754 36660 8760 36712
rect 8812 36700 8818 36712
rect 8849 36703 8907 36709
rect 8849 36700 8861 36703
rect 8812 36672 8861 36700
rect 8812 36660 8818 36672
rect 8849 36669 8861 36672
rect 8895 36669 8907 36703
rect 8849 36663 8907 36669
rect 4387 36604 8156 36632
rect 4387 36601 4399 36604
rect 4341 36595 4399 36601
rect 3050 36564 3056 36576
rect 3011 36536 3056 36564
rect 3050 36524 3056 36536
rect 3108 36524 3114 36576
rect 3605 36567 3663 36573
rect 3605 36533 3617 36567
rect 3651 36564 3663 36567
rect 4890 36564 4896 36576
rect 3651 36536 4896 36564
rect 3651 36533 3663 36536
rect 3605 36527 3663 36533
rect 4890 36524 4896 36536
rect 4948 36524 4954 36576
rect 6454 36524 6460 36576
rect 6512 36564 6518 36576
rect 6825 36567 6883 36573
rect 6825 36564 6837 36567
rect 6512 36536 6837 36564
rect 6512 36524 6518 36536
rect 6825 36533 6837 36536
rect 6871 36533 6883 36567
rect 6825 36527 6883 36533
rect 6914 36524 6920 36576
rect 6972 36564 6978 36576
rect 10244 36564 10272 36740
rect 10965 36737 10977 36740
rect 11011 36737 11023 36771
rect 10965 36731 11023 36737
rect 12253 36771 12311 36777
rect 12253 36737 12265 36771
rect 12299 36737 12311 36771
rect 12253 36731 12311 36737
rect 10870 36660 10876 36712
rect 10928 36700 10934 36712
rect 12268 36700 12296 36731
rect 12342 36728 12348 36780
rect 12400 36768 12406 36780
rect 13556 36777 13584 36876
rect 13630 36864 13636 36916
rect 13688 36904 13694 36916
rect 13688 36876 18460 36904
rect 13688 36864 13694 36876
rect 13722 36796 13728 36848
rect 13780 36836 13786 36848
rect 15378 36836 15384 36848
rect 13780 36808 15384 36836
rect 13780 36796 13786 36808
rect 15378 36796 15384 36808
rect 15436 36796 15442 36848
rect 15565 36839 15623 36845
rect 15565 36805 15577 36839
rect 15611 36836 15623 36839
rect 18432 36836 18460 36876
rect 18506 36864 18512 36916
rect 18564 36904 18570 36916
rect 21726 36904 21732 36916
rect 18564 36876 21732 36904
rect 18564 36864 18570 36876
rect 21726 36864 21732 36876
rect 21784 36864 21790 36916
rect 21818 36864 21824 36916
rect 21876 36904 21882 36916
rect 22002 36904 22008 36916
rect 21876 36876 22008 36904
rect 21876 36864 21882 36876
rect 22002 36864 22008 36876
rect 22060 36864 22066 36916
rect 22094 36864 22100 36916
rect 22152 36904 22158 36916
rect 22189 36907 22247 36913
rect 22189 36904 22201 36907
rect 22152 36876 22201 36904
rect 22152 36864 22158 36876
rect 22189 36873 22201 36876
rect 22235 36873 22247 36907
rect 22189 36867 22247 36873
rect 26145 36907 26203 36913
rect 26145 36873 26157 36907
rect 26191 36904 26203 36907
rect 27798 36904 27804 36916
rect 26191 36876 27804 36904
rect 26191 36873 26203 36876
rect 26145 36867 26203 36873
rect 27798 36864 27804 36876
rect 27856 36864 27862 36916
rect 28718 36864 28724 36916
rect 28776 36904 28782 36916
rect 31018 36904 31024 36916
rect 28776 36876 31024 36904
rect 28776 36864 28782 36876
rect 31018 36864 31024 36876
rect 31076 36864 31082 36916
rect 35713 36907 35771 36913
rect 35713 36873 35725 36907
rect 35759 36904 35771 36907
rect 36817 36907 36875 36913
rect 35759 36876 35894 36904
rect 35759 36873 35771 36876
rect 35713 36867 35771 36873
rect 22738 36836 22744 36848
rect 15611 36808 17618 36836
rect 18432 36808 22744 36836
rect 15611 36805 15623 36808
rect 15565 36799 15623 36805
rect 22738 36796 22744 36808
rect 22796 36796 22802 36848
rect 25130 36836 25136 36848
rect 22848 36808 23428 36836
rect 25091 36808 25136 36836
rect 12897 36771 12955 36777
rect 12897 36768 12909 36771
rect 12400 36740 12909 36768
rect 12400 36728 12406 36740
rect 12897 36737 12909 36740
rect 12943 36737 12955 36771
rect 12897 36731 12955 36737
rect 13541 36771 13599 36777
rect 13541 36737 13553 36771
rect 13587 36737 13599 36771
rect 14182 36768 14188 36780
rect 14143 36740 14188 36768
rect 13541 36731 13599 36737
rect 14182 36728 14188 36740
rect 14240 36728 14246 36780
rect 14829 36771 14887 36777
rect 14829 36737 14841 36771
rect 14875 36768 14887 36771
rect 15194 36768 15200 36780
rect 14875 36740 15200 36768
rect 14875 36737 14887 36740
rect 14829 36731 14887 36737
rect 15194 36728 15200 36740
rect 15252 36728 15258 36780
rect 15473 36771 15531 36777
rect 15473 36737 15485 36771
rect 15519 36768 15531 36771
rect 16117 36771 16175 36777
rect 16117 36768 16129 36771
rect 15519 36740 16129 36768
rect 15519 36737 15531 36740
rect 15473 36731 15531 36737
rect 16117 36737 16129 36740
rect 16163 36768 16175 36771
rect 16758 36768 16764 36780
rect 16163 36740 16764 36768
rect 16163 36737 16175 36740
rect 16117 36731 16175 36737
rect 16758 36728 16764 36740
rect 16816 36728 16822 36780
rect 19334 36728 19340 36780
rect 19392 36768 19398 36780
rect 19392 36740 19437 36768
rect 19392 36728 19398 36740
rect 19518 36728 19524 36780
rect 19576 36768 19582 36780
rect 20349 36771 20407 36777
rect 20349 36768 20361 36771
rect 19576 36740 20361 36768
rect 19576 36728 19582 36740
rect 20349 36737 20361 36740
rect 20395 36768 20407 36771
rect 20993 36771 21051 36777
rect 20993 36768 21005 36771
rect 20395 36740 21005 36768
rect 20395 36737 20407 36740
rect 20349 36731 20407 36737
rect 20993 36737 21005 36740
rect 21039 36768 21051 36771
rect 21082 36768 21088 36780
rect 21039 36740 21088 36768
rect 21039 36737 21051 36740
rect 20993 36731 21051 36737
rect 21082 36728 21088 36740
rect 21140 36768 21146 36780
rect 21450 36768 21456 36780
rect 21140 36740 21456 36768
rect 21140 36728 21146 36740
rect 21450 36728 21456 36740
rect 21508 36728 21514 36780
rect 21542 36728 21548 36780
rect 21600 36768 21606 36780
rect 22005 36771 22063 36777
rect 22005 36768 22017 36771
rect 21600 36740 22017 36768
rect 21600 36728 21606 36740
rect 22005 36737 22017 36740
rect 22051 36737 22063 36771
rect 22005 36731 22063 36737
rect 22094 36728 22100 36780
rect 22152 36768 22158 36780
rect 22848 36768 22876 36808
rect 22152 36740 22876 36768
rect 22152 36728 22158 36740
rect 22922 36728 22928 36780
rect 22980 36768 22986 36780
rect 23400 36777 23428 36808
rect 25130 36796 25136 36808
rect 25188 36796 25194 36848
rect 25222 36796 25228 36848
rect 25280 36836 25286 36848
rect 27430 36836 27436 36848
rect 25280 36808 27436 36836
rect 25280 36796 25286 36808
rect 27430 36796 27436 36808
rect 27488 36796 27494 36848
rect 27525 36839 27583 36845
rect 27525 36805 27537 36839
rect 27571 36836 27583 36839
rect 28810 36836 28816 36848
rect 27571 36808 28816 36836
rect 27571 36805 27583 36808
rect 27525 36799 27583 36805
rect 28810 36796 28816 36808
rect 28868 36796 28874 36848
rect 35866 36836 35894 36876
rect 36817 36873 36829 36907
rect 36863 36904 36875 36907
rect 39298 36904 39304 36916
rect 36863 36876 39304 36904
rect 36863 36873 36875 36876
rect 36817 36867 36875 36873
rect 39298 36864 39304 36876
rect 39356 36864 39362 36916
rect 38105 36839 38163 36845
rect 35866 36808 36676 36836
rect 23385 36771 23443 36777
rect 22980 36740 23025 36768
rect 22980 36728 22986 36740
rect 23385 36737 23397 36771
rect 23431 36768 23443 36771
rect 24029 36771 24087 36777
rect 24029 36768 24041 36771
rect 23431 36740 24041 36768
rect 23431 36737 23443 36740
rect 23385 36731 23443 36737
rect 24029 36737 24041 36740
rect 24075 36737 24087 36771
rect 24029 36731 24087 36737
rect 26329 36771 26387 36777
rect 26329 36737 26341 36771
rect 26375 36768 26387 36771
rect 26970 36768 26976 36780
rect 26375 36740 26976 36768
rect 26375 36737 26387 36740
rect 26329 36731 26387 36737
rect 26970 36728 26976 36740
rect 27028 36728 27034 36780
rect 28626 36728 28632 36780
rect 28684 36768 28690 36780
rect 36648 36777 36676 36808
rect 38105 36805 38117 36839
rect 38151 36836 38163 36839
rect 38654 36836 38660 36848
rect 38151 36808 38660 36836
rect 38151 36805 38163 36808
rect 38105 36799 38163 36805
rect 38654 36796 38660 36808
rect 38712 36796 38718 36848
rect 29089 36771 29147 36777
rect 29089 36768 29101 36771
rect 28684 36740 29101 36768
rect 28684 36728 28690 36740
rect 29089 36737 29101 36740
rect 29135 36737 29147 36771
rect 29089 36731 29147 36737
rect 29549 36771 29607 36777
rect 29549 36737 29561 36771
rect 29595 36737 29607 36771
rect 29549 36731 29607 36737
rect 35069 36771 35127 36777
rect 35069 36737 35081 36771
rect 35115 36737 35127 36771
rect 35069 36731 35127 36737
rect 35161 36771 35219 36777
rect 35161 36737 35173 36771
rect 35207 36768 35219 36771
rect 35897 36771 35955 36777
rect 35897 36768 35909 36771
rect 35207 36740 35909 36768
rect 35207 36737 35219 36740
rect 35161 36731 35219 36737
rect 35897 36737 35909 36740
rect 35943 36737 35955 36771
rect 35897 36731 35955 36737
rect 36633 36771 36691 36777
rect 36633 36737 36645 36771
rect 36679 36737 36691 36771
rect 36633 36731 36691 36737
rect 14550 36700 14556 36712
rect 10928 36672 12296 36700
rect 12820 36672 14556 36700
rect 10928 36660 10934 36672
rect 12345 36635 12403 36641
rect 12345 36601 12357 36635
rect 12391 36632 12403 36635
rect 12710 36632 12716 36644
rect 12391 36604 12716 36632
rect 12391 36601 12403 36604
rect 12345 36595 12403 36601
rect 12710 36592 12716 36604
rect 12768 36592 12774 36644
rect 6972 36536 10272 36564
rect 11057 36567 11115 36573
rect 6972 36524 6978 36536
rect 11057 36533 11069 36567
rect 11103 36564 11115 36567
rect 12820 36564 12848 36672
rect 14550 36660 14556 36672
rect 14608 36660 14614 36712
rect 16482 36660 16488 36712
rect 16540 36700 16546 36712
rect 16853 36703 16911 36709
rect 16853 36700 16865 36703
rect 16540 36672 16865 36700
rect 16540 36660 16546 36672
rect 16853 36669 16865 36672
rect 16899 36669 16911 36703
rect 17586 36700 17592 36712
rect 16853 36663 16911 36669
rect 16960 36672 17592 36700
rect 14458 36592 14464 36644
rect 14516 36632 14522 36644
rect 16960 36632 16988 36672
rect 17586 36660 17592 36672
rect 17644 36660 17650 36712
rect 17678 36660 17684 36712
rect 17736 36700 17742 36712
rect 19429 36703 19487 36709
rect 19429 36700 19441 36703
rect 17736 36672 19441 36700
rect 17736 36660 17742 36672
rect 19429 36669 19441 36672
rect 19475 36669 19487 36703
rect 19429 36663 19487 36669
rect 20898 36660 20904 36712
rect 20956 36700 20962 36712
rect 24121 36703 24179 36709
rect 24121 36700 24133 36703
rect 20956 36672 24133 36700
rect 20956 36660 20962 36672
rect 24121 36669 24133 36672
rect 24167 36669 24179 36703
rect 25038 36700 25044 36712
rect 24999 36672 25044 36700
rect 24121 36663 24179 36669
rect 25038 36660 25044 36672
rect 25096 36660 25102 36712
rect 25222 36660 25228 36712
rect 25280 36700 25286 36712
rect 25317 36703 25375 36709
rect 25317 36700 25329 36703
rect 25280 36672 25329 36700
rect 25280 36660 25286 36672
rect 25317 36669 25329 36672
rect 25363 36700 25375 36703
rect 27433 36703 27491 36709
rect 25363 36672 27384 36700
rect 25363 36669 25375 36672
rect 25317 36663 25375 36669
rect 14516 36604 16988 36632
rect 14516 36592 14522 36604
rect 20714 36592 20720 36644
rect 20772 36632 20778 36644
rect 22741 36635 22799 36641
rect 22741 36632 22753 36635
rect 20772 36604 22753 36632
rect 20772 36592 20778 36604
rect 22741 36601 22753 36604
rect 22787 36601 22799 36635
rect 22741 36595 22799 36601
rect 25130 36592 25136 36644
rect 25188 36632 25194 36644
rect 27246 36632 27252 36644
rect 25188 36604 27252 36632
rect 25188 36592 25194 36604
rect 27246 36592 27252 36604
rect 27304 36592 27310 36644
rect 27356 36632 27384 36672
rect 27433 36669 27445 36703
rect 27479 36700 27491 36703
rect 27522 36700 27528 36712
rect 27479 36672 27528 36700
rect 27479 36669 27491 36672
rect 27433 36663 27491 36669
rect 27522 36660 27528 36672
rect 27580 36700 27586 36712
rect 28350 36700 28356 36712
rect 27580 36672 28212 36700
rect 28311 36672 28356 36700
rect 27580 36660 27586 36672
rect 27982 36632 27988 36644
rect 27356 36604 27988 36632
rect 27982 36592 27988 36604
rect 28040 36592 28046 36644
rect 12986 36564 12992 36576
rect 11103 36536 12848 36564
rect 12947 36536 12992 36564
rect 11103 36533 11115 36536
rect 11057 36527 11115 36533
rect 12986 36524 12992 36536
rect 13044 36524 13050 36576
rect 13630 36564 13636 36576
rect 13591 36536 13636 36564
rect 13630 36524 13636 36536
rect 13688 36524 13694 36576
rect 14277 36567 14335 36573
rect 14277 36533 14289 36567
rect 14323 36564 14335 36567
rect 14826 36564 14832 36576
rect 14323 36536 14832 36564
rect 14323 36533 14335 36536
rect 14277 36527 14335 36533
rect 14826 36524 14832 36536
rect 14884 36524 14890 36576
rect 14918 36524 14924 36576
rect 14976 36564 14982 36576
rect 16206 36564 16212 36576
rect 14976 36536 15021 36564
rect 16167 36536 16212 36564
rect 14976 36524 14982 36536
rect 16206 36524 16212 36536
rect 16264 36524 16270 36576
rect 17126 36573 17132 36576
rect 17116 36567 17132 36573
rect 17116 36533 17128 36567
rect 17116 36527 17132 36533
rect 17126 36524 17132 36527
rect 17184 36524 17190 36576
rect 18598 36564 18604 36576
rect 18559 36536 18604 36564
rect 18598 36524 18604 36536
rect 18656 36524 18662 36576
rect 20438 36564 20444 36576
rect 20399 36536 20444 36564
rect 20438 36524 20444 36536
rect 20496 36524 20502 36576
rect 20990 36524 20996 36576
rect 21048 36564 21054 36576
rect 21085 36567 21143 36573
rect 21085 36564 21097 36567
rect 21048 36536 21097 36564
rect 21048 36524 21054 36536
rect 21085 36533 21097 36536
rect 21131 36533 21143 36567
rect 21085 36527 21143 36533
rect 21174 36524 21180 36576
rect 21232 36564 21238 36576
rect 22462 36564 22468 36576
rect 21232 36536 22468 36564
rect 21232 36524 21238 36536
rect 22462 36524 22468 36536
rect 22520 36524 22526 36576
rect 23014 36524 23020 36576
rect 23072 36564 23078 36576
rect 23477 36567 23535 36573
rect 23477 36564 23489 36567
rect 23072 36536 23489 36564
rect 23072 36524 23078 36536
rect 23477 36533 23489 36536
rect 23523 36533 23535 36567
rect 28184 36564 28212 36672
rect 28350 36660 28356 36672
rect 28408 36660 28414 36712
rect 29564 36700 29592 36731
rect 28920 36672 29592 36700
rect 28920 36641 28948 36672
rect 28905 36635 28963 36641
rect 28905 36601 28917 36635
rect 28951 36601 28963 36635
rect 28905 36595 28963 36601
rect 29730 36592 29736 36644
rect 29788 36632 29794 36644
rect 35084 36632 35112 36731
rect 29788 36604 35112 36632
rect 29788 36592 29794 36604
rect 29641 36567 29699 36573
rect 29641 36564 29653 36567
rect 28184 36536 29653 36564
rect 23477 36527 23535 36533
rect 29641 36533 29653 36536
rect 29687 36533 29699 36567
rect 38194 36564 38200 36576
rect 38155 36536 38200 36564
rect 29641 36527 29699 36533
rect 38194 36524 38200 36536
rect 38252 36524 38258 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 1581 36363 1639 36369
rect 1581 36329 1593 36363
rect 1627 36360 1639 36363
rect 2958 36360 2964 36372
rect 1627 36332 2964 36360
rect 1627 36329 1639 36332
rect 1581 36323 1639 36329
rect 2958 36320 2964 36332
rect 3016 36320 3022 36372
rect 3970 36360 3976 36372
rect 3931 36332 3976 36360
rect 3970 36320 3976 36332
rect 4028 36320 4034 36372
rect 4614 36320 4620 36372
rect 4672 36360 4678 36372
rect 7926 36360 7932 36372
rect 4672 36332 7788 36360
rect 7887 36332 7932 36360
rect 4672 36320 4678 36332
rect 3050 36252 3056 36304
rect 3108 36292 3114 36304
rect 3108 36264 6408 36292
rect 3108 36252 3114 36264
rect 4798 36224 4804 36236
rect 4759 36196 4804 36224
rect 4798 36184 4804 36196
rect 4856 36184 4862 36236
rect 5813 36227 5871 36233
rect 5813 36193 5825 36227
rect 5859 36224 5871 36227
rect 5902 36224 5908 36236
rect 5859 36196 5908 36224
rect 5859 36193 5871 36196
rect 5813 36187 5871 36193
rect 5902 36184 5908 36196
rect 5960 36184 5966 36236
rect 6380 36233 6408 36264
rect 6365 36227 6423 36233
rect 6365 36193 6377 36227
rect 6411 36193 6423 36227
rect 7760 36224 7788 36332
rect 7926 36320 7932 36332
rect 7984 36320 7990 36372
rect 8478 36320 8484 36372
rect 8536 36360 8542 36372
rect 12342 36360 12348 36372
rect 8536 36332 12348 36360
rect 8536 36320 8542 36332
rect 12342 36320 12348 36332
rect 12400 36320 12406 36372
rect 12710 36320 12716 36372
rect 12768 36360 12774 36372
rect 14734 36360 14740 36372
rect 12768 36332 14740 36360
rect 12768 36320 12774 36332
rect 14734 36320 14740 36332
rect 14792 36320 14798 36372
rect 14826 36320 14832 36372
rect 14884 36360 14890 36372
rect 22922 36360 22928 36372
rect 14884 36332 22928 36360
rect 14884 36320 14890 36332
rect 22922 36320 22928 36332
rect 22980 36320 22986 36372
rect 24394 36320 24400 36372
rect 24452 36360 24458 36372
rect 24452 36332 25820 36360
rect 24452 36320 24458 36332
rect 17494 36252 17500 36304
rect 17552 36292 17558 36304
rect 21174 36292 21180 36304
rect 17552 36264 21180 36292
rect 17552 36252 17558 36264
rect 21174 36252 21180 36264
rect 21232 36252 21238 36304
rect 21634 36252 21640 36304
rect 21692 36292 21698 36304
rect 25792 36292 25820 36332
rect 25866 36320 25872 36372
rect 25924 36360 25930 36372
rect 26697 36363 26755 36369
rect 26697 36360 26709 36363
rect 25924 36332 26709 36360
rect 25924 36320 25930 36332
rect 26697 36329 26709 36332
rect 26743 36329 26755 36363
rect 26697 36323 26755 36329
rect 27430 36320 27436 36372
rect 27488 36360 27494 36372
rect 27488 36332 31754 36360
rect 27488 36320 27494 36332
rect 31726 36292 31754 36332
rect 37182 36320 37188 36372
rect 37240 36360 37246 36372
rect 37461 36363 37519 36369
rect 37461 36360 37473 36363
rect 37240 36332 37473 36360
rect 37240 36320 37246 36332
rect 37461 36329 37473 36332
rect 37507 36329 37519 36363
rect 37461 36323 37519 36329
rect 33042 36292 33048 36304
rect 21692 36264 25636 36292
rect 25792 36264 28672 36292
rect 31726 36264 33048 36292
rect 21692 36252 21698 36264
rect 11977 36227 12035 36233
rect 7760 36196 9536 36224
rect 6365 36187 6423 36193
rect 1302 36116 1308 36168
rect 1360 36156 1366 36168
rect 1765 36159 1823 36165
rect 1765 36156 1777 36159
rect 1360 36128 1777 36156
rect 1360 36116 1366 36128
rect 1765 36125 1777 36128
rect 1811 36125 1823 36159
rect 1765 36119 1823 36125
rect 2869 36159 2927 36165
rect 2869 36125 2881 36159
rect 2915 36125 2927 36159
rect 4154 36156 4160 36168
rect 4115 36128 4160 36156
rect 2869 36119 2927 36125
rect 2682 36020 2688 36032
rect 2643 35992 2688 36020
rect 2682 35980 2688 35992
rect 2740 35980 2746 36032
rect 2884 36020 2912 36119
rect 4154 36116 4160 36128
rect 4212 36116 4218 36168
rect 7837 36159 7895 36165
rect 5644 36128 6040 36156
rect 4890 36088 4896 36100
rect 4851 36060 4896 36088
rect 4890 36048 4896 36060
rect 4948 36048 4954 36100
rect 4982 36048 4988 36100
rect 5040 36088 5046 36100
rect 5644 36088 5672 36128
rect 5040 36060 5672 36088
rect 5040 36048 5046 36060
rect 5902 36020 5908 36032
rect 2884 35992 5908 36020
rect 5902 35980 5908 35992
rect 5960 35980 5966 36032
rect 6012 36020 6040 36128
rect 7837 36125 7849 36159
rect 7883 36125 7895 36159
rect 7837 36119 7895 36125
rect 6454 36048 6460 36100
rect 6512 36088 6518 36100
rect 7374 36088 7380 36100
rect 6512 36060 6557 36088
rect 7335 36060 7380 36088
rect 6512 36048 6518 36060
rect 7374 36048 7380 36060
rect 7432 36048 7438 36100
rect 7852 36020 7880 36119
rect 8294 36048 8300 36100
rect 8352 36088 8358 36100
rect 9398 36088 9404 36100
rect 8352 36060 9404 36088
rect 8352 36048 8358 36060
rect 9398 36048 9404 36060
rect 9456 36048 9462 36100
rect 6012 35992 7880 36020
rect 9125 36023 9183 36029
rect 9125 35989 9137 36023
rect 9171 36020 9183 36023
rect 9214 36020 9220 36032
rect 9171 35992 9220 36020
rect 9171 35989 9183 35992
rect 9125 35983 9183 35989
rect 9214 35980 9220 35992
rect 9272 35980 9278 36032
rect 9508 36020 9536 36196
rect 11977 36193 11989 36227
rect 12023 36224 12035 36227
rect 14458 36224 14464 36236
rect 12023 36196 14464 36224
rect 12023 36193 12035 36196
rect 11977 36187 12035 36193
rect 14458 36184 14464 36196
rect 14516 36184 14522 36236
rect 15841 36227 15899 36233
rect 15841 36193 15853 36227
rect 15887 36224 15899 36227
rect 16482 36224 16488 36236
rect 15887 36196 16488 36224
rect 15887 36193 15899 36196
rect 15841 36187 15899 36193
rect 16482 36184 16488 36196
rect 16540 36184 16546 36236
rect 16758 36184 16764 36236
rect 16816 36224 16822 36236
rect 20438 36224 20444 36236
rect 16816 36196 20444 36224
rect 16816 36184 16822 36196
rect 20438 36184 20444 36196
rect 20496 36184 20502 36236
rect 22554 36224 22560 36236
rect 21192 36196 22560 36224
rect 11698 36156 11704 36168
rect 11659 36128 11704 36156
rect 11698 36116 11704 36128
rect 11756 36116 11762 36168
rect 14366 36156 14372 36168
rect 13110 36128 14372 36156
rect 14366 36116 14372 36128
rect 14424 36116 14430 36168
rect 14553 36159 14611 36165
rect 14553 36125 14565 36159
rect 14599 36156 14611 36159
rect 15010 36156 15016 36168
rect 14599 36128 15016 36156
rect 14599 36125 14611 36128
rect 14553 36119 14611 36125
rect 15010 36116 15016 36128
rect 15068 36116 15074 36168
rect 15194 36156 15200 36168
rect 15107 36128 15200 36156
rect 15194 36116 15200 36128
rect 15252 36156 15258 36168
rect 15252 36128 15884 36156
rect 15252 36116 15258 36128
rect 13722 36088 13728 36100
rect 13683 36060 13728 36088
rect 13722 36048 13728 36060
rect 13780 36048 13786 36100
rect 14645 36091 14703 36097
rect 14645 36057 14657 36091
rect 14691 36088 14703 36091
rect 15856 36088 15884 36128
rect 18506 36116 18512 36168
rect 18564 36156 18570 36168
rect 18693 36159 18751 36165
rect 18693 36156 18705 36159
rect 18564 36128 18705 36156
rect 18564 36116 18570 36128
rect 18693 36125 18705 36128
rect 18739 36156 18751 36159
rect 19889 36159 19947 36165
rect 19889 36156 19901 36159
rect 18739 36128 19901 36156
rect 18739 36125 18751 36128
rect 18693 36119 18751 36125
rect 19889 36125 19901 36128
rect 19935 36156 19947 36159
rect 20162 36156 20168 36168
rect 19935 36128 20168 36156
rect 19935 36125 19947 36128
rect 19889 36119 19947 36125
rect 20162 36116 20168 36128
rect 20220 36116 20226 36168
rect 20625 36159 20683 36165
rect 20625 36125 20637 36159
rect 20671 36156 20683 36159
rect 21082 36156 21088 36168
rect 20671 36128 21088 36156
rect 20671 36125 20683 36128
rect 20625 36119 20683 36125
rect 21082 36116 21088 36128
rect 21140 36116 21146 36168
rect 16022 36088 16028 36100
rect 14691 36060 15608 36088
rect 15856 36060 16028 36088
rect 14691 36057 14703 36060
rect 14645 36051 14703 36057
rect 13906 36020 13912 36032
rect 9508 35992 13912 36020
rect 13906 35980 13912 35992
rect 13964 35980 13970 36032
rect 14090 35980 14096 36032
rect 14148 36020 14154 36032
rect 15194 36020 15200 36032
rect 14148 35992 15200 36020
rect 14148 35980 14154 35992
rect 15194 35980 15200 35992
rect 15252 35980 15258 36032
rect 15289 36023 15347 36029
rect 15289 35989 15301 36023
rect 15335 36020 15347 36023
rect 15378 36020 15384 36032
rect 15335 35992 15384 36020
rect 15335 35989 15347 35992
rect 15289 35983 15347 35989
rect 15378 35980 15384 35992
rect 15436 35980 15442 36032
rect 15580 36020 15608 36060
rect 16022 36048 16028 36060
rect 16080 36048 16086 36100
rect 16114 36048 16120 36100
rect 16172 36088 16178 36100
rect 16172 36060 16217 36088
rect 16316 36060 16606 36088
rect 16172 36048 16178 36060
rect 16316 36020 16344 36060
rect 15580 35992 16344 36020
rect 16850 35980 16856 36032
rect 16908 36020 16914 36032
rect 17589 36023 17647 36029
rect 17589 36020 17601 36023
rect 16908 35992 17601 36020
rect 16908 35980 16914 35992
rect 17589 35989 17601 35992
rect 17635 35989 17647 36023
rect 17589 35983 17647 35989
rect 17954 35980 17960 36032
rect 18012 36020 18018 36032
rect 18785 36023 18843 36029
rect 18785 36020 18797 36023
rect 18012 35992 18797 36020
rect 18012 35980 18018 35992
rect 18785 35989 18797 35992
rect 18831 35989 18843 36023
rect 19978 36020 19984 36032
rect 19939 35992 19984 36020
rect 18785 35983 18843 35989
rect 19978 35980 19984 35992
rect 20036 35980 20042 36032
rect 20714 36020 20720 36032
rect 20675 35992 20720 36020
rect 20714 35980 20720 35992
rect 20772 35980 20778 36032
rect 21192 36020 21220 36196
rect 22554 36184 22560 36196
rect 22612 36184 22618 36236
rect 22738 36184 22744 36236
rect 22796 36224 22802 36236
rect 25498 36224 25504 36236
rect 22796 36196 24624 36224
rect 25459 36196 25504 36224
rect 22796 36184 22802 36196
rect 24596 36165 24624 36196
rect 25498 36184 25504 36196
rect 25556 36184 25562 36236
rect 25608 36224 25636 36264
rect 25777 36227 25835 36233
rect 25777 36224 25789 36227
rect 25608 36196 25789 36224
rect 25777 36193 25789 36196
rect 25823 36224 25835 36227
rect 27522 36224 27528 36236
rect 25823 36196 26648 36224
rect 27483 36196 27528 36224
rect 25823 36193 25835 36196
rect 25777 36187 25835 36193
rect 26620 36165 26648 36196
rect 27522 36184 27528 36196
rect 27580 36184 27586 36236
rect 27614 36184 27620 36236
rect 27672 36224 27678 36236
rect 27672 36196 28580 36224
rect 27672 36184 27678 36196
rect 24581 36159 24639 36165
rect 24581 36125 24593 36159
rect 24627 36125 24639 36159
rect 24581 36119 24639 36125
rect 26605 36159 26663 36165
rect 26605 36125 26617 36159
rect 26651 36125 26663 36159
rect 26605 36119 26663 36125
rect 21358 36088 21364 36100
rect 21319 36060 21364 36088
rect 21358 36048 21364 36060
rect 21416 36048 21422 36100
rect 21453 36091 21511 36097
rect 21453 36057 21465 36091
rect 21499 36057 21511 36091
rect 21453 36051 21511 36057
rect 21468 36020 21496 36051
rect 21634 36048 21640 36100
rect 21692 36088 21698 36100
rect 22005 36091 22063 36097
rect 22005 36088 22017 36091
rect 21692 36060 22017 36088
rect 21692 36048 21698 36060
rect 22005 36057 22017 36060
rect 22051 36057 22063 36091
rect 22005 36051 22063 36057
rect 22278 36048 22284 36100
rect 22336 36088 22342 36100
rect 22557 36091 22615 36097
rect 22557 36088 22569 36091
rect 22336 36060 22569 36088
rect 22336 36048 22342 36060
rect 22557 36057 22569 36060
rect 22603 36057 22615 36091
rect 22557 36051 22615 36057
rect 22649 36091 22707 36097
rect 22649 36057 22661 36091
rect 22695 36057 22707 36091
rect 22649 36051 22707 36057
rect 23569 36091 23627 36097
rect 23569 36057 23581 36091
rect 23615 36088 23627 36091
rect 25590 36088 25596 36100
rect 23615 36060 25452 36088
rect 25551 36060 25596 36088
rect 23615 36057 23627 36060
rect 23569 36051 23627 36057
rect 21192 35992 21496 36020
rect 21726 35980 21732 36032
rect 21784 36020 21790 36032
rect 22664 36020 22692 36051
rect 21784 35992 22692 36020
rect 21784 35980 21790 35992
rect 23474 35980 23480 36032
rect 23532 36020 23538 36032
rect 24673 36023 24731 36029
rect 24673 36020 24685 36023
rect 23532 35992 24685 36020
rect 23532 35980 23538 35992
rect 24673 35989 24685 35992
rect 24719 35989 24731 36023
rect 25424 36020 25452 36060
rect 25590 36048 25596 36060
rect 25648 36048 25654 36100
rect 27617 36091 27675 36097
rect 27617 36057 27629 36091
rect 27663 36088 27675 36091
rect 27663 36060 27936 36088
rect 27663 36057 27675 36060
rect 27617 36051 27675 36057
rect 26786 36020 26792 36032
rect 25424 35992 26792 36020
rect 24673 35983 24731 35989
rect 26786 35980 26792 35992
rect 26844 35980 26850 36032
rect 26970 35980 26976 36032
rect 27028 36020 27034 36032
rect 27522 36020 27528 36032
rect 27028 35992 27528 36020
rect 27028 35980 27034 35992
rect 27522 35980 27528 35992
rect 27580 35980 27586 36032
rect 27908 36020 27936 36060
rect 27982 36048 27988 36100
rect 28040 36088 28046 36100
rect 28169 36091 28227 36097
rect 28169 36088 28181 36091
rect 28040 36060 28181 36088
rect 28040 36048 28046 36060
rect 28169 36057 28181 36060
rect 28215 36057 28227 36091
rect 28552 36088 28580 36196
rect 28644 36165 28672 36264
rect 33042 36252 33048 36264
rect 33100 36252 33106 36304
rect 38194 36292 38200 36304
rect 35866 36264 38200 36292
rect 35866 36224 35894 36264
rect 38194 36252 38200 36264
rect 38252 36252 38258 36304
rect 31726 36196 35894 36224
rect 28629 36159 28687 36165
rect 28629 36125 28641 36159
rect 28675 36125 28687 36159
rect 28629 36119 28687 36125
rect 31726 36088 31754 36196
rect 36078 36116 36084 36168
rect 36136 36156 36142 36168
rect 36357 36159 36415 36165
rect 36357 36156 36369 36159
rect 36136 36128 36369 36156
rect 36136 36116 36142 36128
rect 36357 36125 36369 36128
rect 36403 36125 36415 36159
rect 37274 36156 37280 36168
rect 37235 36128 37280 36156
rect 36357 36119 36415 36125
rect 37274 36116 37280 36128
rect 37332 36116 37338 36168
rect 38013 36159 38071 36165
rect 38013 36125 38025 36159
rect 38059 36125 38071 36159
rect 38013 36119 38071 36125
rect 28552 36060 31754 36088
rect 28169 36051 28227 36057
rect 36538 36048 36544 36100
rect 36596 36088 36602 36100
rect 38028 36088 38056 36119
rect 36596 36060 38056 36088
rect 36596 36048 36602 36060
rect 28721 36023 28779 36029
rect 28721 36020 28733 36023
rect 27908 35992 28733 36020
rect 28721 35989 28733 35992
rect 28767 35989 28779 36023
rect 28721 35983 28779 35989
rect 34514 35980 34520 36032
rect 34572 36020 34578 36032
rect 36173 36023 36231 36029
rect 36173 36020 36185 36023
rect 34572 35992 36185 36020
rect 34572 35980 34578 35992
rect 36173 35989 36185 35992
rect 36219 35989 36231 36023
rect 38194 36020 38200 36032
rect 38155 35992 38200 36020
rect 36173 35983 36231 35989
rect 38194 35980 38200 35992
rect 38252 35980 38258 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 3329 35819 3387 35825
rect 3329 35785 3341 35819
rect 3375 35785 3387 35819
rect 5902 35816 5908 35828
rect 5863 35788 5908 35816
rect 3329 35779 3387 35785
rect 3234 35748 3240 35760
rect 3082 35720 3240 35748
rect 3234 35708 3240 35720
rect 3292 35708 3298 35760
rect 3344 35748 3372 35779
rect 5902 35776 5908 35788
rect 5960 35776 5966 35828
rect 7208 35788 11284 35816
rect 7208 35757 7236 35788
rect 7193 35751 7251 35757
rect 7193 35748 7205 35751
rect 3344 35720 7205 35748
rect 7193 35717 7205 35720
rect 7239 35717 7251 35751
rect 9398 35748 9404 35760
rect 9359 35720 9404 35748
rect 7193 35711 7251 35717
rect 9398 35708 9404 35720
rect 9456 35708 9462 35760
rect 5813 35683 5871 35689
rect 5813 35649 5825 35683
rect 5859 35680 5871 35683
rect 6822 35680 6828 35692
rect 5859 35652 6828 35680
rect 5859 35649 5871 35652
rect 5813 35643 5871 35649
rect 6822 35640 6828 35652
rect 6880 35640 6886 35692
rect 1578 35612 1584 35624
rect 1539 35584 1584 35612
rect 1578 35572 1584 35584
rect 1636 35572 1642 35624
rect 1857 35615 1915 35621
rect 1857 35581 1869 35615
rect 1903 35612 1915 35615
rect 4154 35612 4160 35624
rect 1903 35584 4160 35612
rect 1903 35581 1915 35584
rect 1857 35575 1915 35581
rect 4154 35572 4160 35584
rect 4212 35572 4218 35624
rect 4614 35572 4620 35624
rect 4672 35612 4678 35624
rect 5442 35612 5448 35624
rect 4672 35584 5448 35612
rect 4672 35572 4678 35584
rect 5442 35572 5448 35584
rect 5500 35612 5506 35624
rect 6917 35615 6975 35621
rect 6917 35612 6929 35615
rect 5500 35584 6929 35612
rect 5500 35572 5506 35584
rect 6917 35581 6929 35584
rect 6963 35581 6975 35615
rect 6917 35575 6975 35581
rect 8312 35544 8340 35666
rect 10502 35640 10508 35692
rect 10560 35640 10566 35692
rect 9122 35612 9128 35624
rect 9083 35584 9128 35612
rect 9122 35572 9128 35584
rect 9180 35572 9186 35624
rect 9398 35572 9404 35624
rect 9456 35612 9462 35624
rect 9456 35584 10824 35612
rect 9456 35572 9462 35584
rect 10796 35544 10824 35584
rect 10870 35572 10876 35624
rect 10928 35612 10934 35624
rect 11149 35615 11207 35621
rect 11149 35612 11161 35615
rect 10928 35584 11161 35612
rect 10928 35572 10934 35584
rect 11149 35581 11161 35584
rect 11195 35581 11207 35615
rect 11256 35612 11284 35788
rect 12434 35776 12440 35828
rect 12492 35816 12498 35828
rect 13722 35816 13728 35828
rect 12492 35788 13728 35816
rect 12492 35776 12498 35788
rect 13722 35776 13728 35788
rect 13780 35776 13786 35828
rect 13998 35816 14004 35828
rect 13959 35788 14004 35816
rect 13998 35776 14004 35788
rect 14056 35776 14062 35828
rect 15194 35776 15200 35828
rect 15252 35816 15258 35828
rect 18690 35816 18696 35828
rect 15252 35788 18696 35816
rect 15252 35776 15258 35788
rect 18690 35776 18696 35788
rect 18748 35776 18754 35828
rect 22002 35776 22008 35828
rect 22060 35816 22066 35828
rect 22060 35788 25544 35816
rect 22060 35776 22066 35788
rect 11330 35708 11336 35760
rect 11388 35748 11394 35760
rect 15102 35748 15108 35760
rect 11388 35720 15108 35748
rect 11388 35708 11394 35720
rect 15102 35708 15108 35720
rect 15160 35708 15166 35760
rect 16298 35708 16304 35760
rect 16356 35748 16362 35760
rect 17218 35748 17224 35760
rect 16356 35720 17224 35748
rect 16356 35708 16362 35720
rect 17218 35708 17224 35720
rect 17276 35708 17282 35760
rect 17402 35708 17408 35760
rect 17460 35748 17466 35760
rect 17460 35720 17618 35748
rect 17460 35708 17466 35720
rect 19794 35708 19800 35760
rect 19852 35748 19858 35760
rect 20346 35748 20352 35760
rect 19852 35720 20352 35748
rect 19852 35708 19858 35720
rect 20346 35708 20352 35720
rect 20404 35708 20410 35760
rect 20806 35748 20812 35760
rect 20767 35720 20812 35748
rect 20806 35708 20812 35720
rect 20864 35708 20870 35760
rect 20901 35751 20959 35757
rect 20901 35717 20913 35751
rect 20947 35748 20959 35751
rect 22186 35748 22192 35760
rect 20947 35720 22192 35748
rect 20947 35717 20959 35720
rect 20901 35711 20959 35717
rect 22186 35708 22192 35720
rect 22244 35708 22250 35760
rect 22646 35708 22652 35760
rect 22704 35748 22710 35760
rect 23201 35751 23259 35757
rect 23201 35748 23213 35751
rect 22704 35720 23213 35748
rect 22704 35708 22710 35720
rect 23201 35717 23213 35720
rect 23247 35717 23259 35751
rect 23201 35711 23259 35717
rect 23293 35751 23351 35757
rect 23293 35717 23305 35751
rect 23339 35748 23351 35751
rect 25130 35748 25136 35760
rect 23339 35720 25136 35748
rect 23339 35717 23351 35720
rect 23293 35711 23351 35717
rect 25130 35708 25136 35720
rect 25188 35708 25194 35760
rect 25406 35748 25412 35760
rect 25367 35720 25412 35748
rect 25406 35708 25412 35720
rect 25464 35708 25470 35760
rect 25516 35748 25544 35788
rect 26418 35776 26424 35828
rect 26476 35816 26482 35828
rect 28626 35816 28632 35828
rect 26476 35788 28632 35816
rect 26476 35776 26482 35788
rect 28626 35776 28632 35788
rect 28684 35776 28690 35828
rect 28810 35816 28816 35828
rect 28771 35788 28816 35816
rect 28810 35776 28816 35788
rect 28868 35776 28874 35828
rect 27246 35748 27252 35760
rect 25516 35720 26556 35748
rect 27207 35720 27252 35748
rect 11422 35640 11428 35692
rect 11480 35680 11486 35692
rect 12437 35683 12495 35689
rect 12437 35680 12449 35683
rect 11480 35652 12449 35680
rect 11480 35640 11486 35652
rect 12437 35649 12449 35652
rect 12483 35649 12495 35683
rect 13906 35680 13912 35692
rect 13867 35652 13912 35680
rect 12437 35643 12495 35649
rect 13906 35640 13912 35652
rect 13964 35640 13970 35692
rect 14090 35612 14096 35624
rect 11256 35584 14096 35612
rect 11149 35575 11207 35581
rect 14090 35572 14096 35584
rect 14148 35572 14154 35624
rect 14553 35615 14611 35621
rect 14553 35581 14565 35615
rect 14599 35581 14611 35615
rect 14826 35612 14832 35624
rect 14787 35584 14832 35612
rect 14553 35575 14611 35581
rect 12434 35544 12440 35556
rect 8312 35516 9260 35544
rect 10796 35516 12440 35544
rect 4154 35436 4160 35488
rect 4212 35476 4218 35488
rect 7006 35476 7012 35488
rect 4212 35448 7012 35476
rect 4212 35436 4218 35448
rect 7006 35436 7012 35448
rect 7064 35476 7070 35488
rect 8202 35476 8208 35488
rect 7064 35448 8208 35476
rect 7064 35436 7070 35448
rect 8202 35436 8208 35448
rect 8260 35436 8266 35488
rect 8662 35476 8668 35488
rect 8623 35448 8668 35476
rect 8662 35436 8668 35448
rect 8720 35436 8726 35488
rect 9232 35476 9260 35516
rect 12434 35504 12440 35516
rect 12492 35504 12498 35556
rect 12529 35547 12587 35553
rect 12529 35513 12541 35547
rect 12575 35544 12587 35547
rect 14458 35544 14464 35556
rect 12575 35516 14464 35544
rect 12575 35513 12587 35516
rect 12529 35507 12587 35513
rect 14458 35504 14464 35516
rect 14516 35504 14522 35556
rect 13446 35476 13452 35488
rect 9232 35448 13452 35476
rect 13446 35436 13452 35448
rect 13504 35436 13510 35488
rect 14568 35476 14596 35575
rect 14826 35572 14832 35584
rect 14884 35572 14890 35624
rect 15194 35572 15200 35624
rect 15252 35612 15258 35624
rect 15948 35612 15976 35666
rect 16482 35640 16488 35692
rect 16540 35680 16546 35692
rect 16853 35683 16911 35689
rect 16853 35680 16865 35683
rect 16540 35652 16865 35680
rect 16540 35640 16546 35652
rect 16853 35649 16865 35652
rect 16899 35649 16911 35683
rect 16853 35643 16911 35649
rect 18690 35640 18696 35692
rect 18748 35680 18754 35692
rect 19245 35683 19303 35689
rect 19245 35680 19257 35683
rect 18748 35652 19257 35680
rect 18748 35640 18754 35652
rect 19245 35649 19257 35652
rect 19291 35649 19303 35683
rect 19245 35643 19303 35649
rect 19889 35683 19947 35689
rect 19889 35649 19901 35683
rect 19935 35680 19947 35683
rect 20162 35680 20168 35692
rect 19935 35652 20168 35680
rect 19935 35649 19947 35652
rect 19889 35643 19947 35649
rect 20162 35640 20168 35652
rect 20220 35680 20226 35692
rect 20530 35680 20536 35692
rect 20220 35652 20536 35680
rect 20220 35640 20226 35652
rect 20530 35640 20536 35652
rect 20588 35640 20594 35692
rect 21453 35683 21511 35689
rect 21453 35649 21465 35683
rect 21499 35680 21511 35683
rect 21634 35680 21640 35692
rect 21499 35652 21640 35680
rect 21499 35649 21511 35652
rect 21453 35643 21511 35649
rect 21634 35640 21640 35652
rect 21692 35640 21698 35692
rect 21818 35640 21824 35692
rect 21876 35680 21882 35692
rect 22465 35683 22523 35689
rect 22465 35680 22477 35683
rect 21876 35652 22477 35680
rect 21876 35640 21882 35652
rect 22465 35649 22477 35652
rect 22511 35649 22523 35683
rect 22465 35643 22523 35649
rect 24305 35683 24363 35689
rect 24305 35649 24317 35683
rect 24351 35649 24363 35683
rect 24305 35643 24363 35649
rect 26421 35683 26479 35689
rect 26421 35649 26433 35683
rect 26467 35649 26479 35683
rect 26528 35680 26556 35720
rect 27246 35708 27252 35720
rect 27304 35708 27310 35760
rect 28902 35748 28908 35760
rect 28000 35720 28908 35748
rect 27157 35683 27215 35689
rect 27157 35680 27169 35683
rect 26528 35652 27169 35680
rect 26421 35643 26479 35649
rect 27157 35649 27169 35652
rect 27203 35649 27215 35683
rect 27157 35643 27215 35649
rect 17126 35612 17132 35624
rect 15252 35584 15884 35612
rect 15948 35584 16988 35612
rect 17087 35584 17132 35612
rect 15252 35572 15258 35584
rect 15194 35476 15200 35488
rect 14568 35448 15200 35476
rect 15194 35436 15200 35448
rect 15252 35436 15258 35488
rect 15856 35476 15884 35584
rect 16298 35544 16304 35556
rect 16259 35516 16304 35544
rect 16298 35504 16304 35516
rect 16356 35504 16362 35556
rect 16666 35476 16672 35488
rect 15856 35448 16672 35476
rect 16666 35436 16672 35448
rect 16724 35436 16730 35488
rect 16960 35476 16988 35584
rect 17126 35572 17132 35584
rect 17184 35572 17190 35624
rect 17218 35572 17224 35624
rect 17276 35612 17282 35624
rect 17276 35584 23244 35612
rect 17276 35572 17282 35584
rect 20898 35544 20904 35556
rect 18524 35516 20904 35544
rect 18524 35476 18552 35516
rect 20898 35504 20904 35516
rect 20956 35504 20962 35556
rect 21266 35504 21272 35556
rect 21324 35544 21330 35556
rect 23216 35544 23244 35584
rect 23290 35572 23296 35624
rect 23348 35612 23354 35624
rect 23477 35615 23535 35621
rect 23477 35612 23489 35615
rect 23348 35584 23489 35612
rect 23348 35572 23354 35584
rect 23477 35581 23489 35584
rect 23523 35581 23535 35615
rect 24320 35612 24348 35643
rect 23477 35575 23535 35581
rect 23584 35584 24348 35612
rect 25317 35615 25375 35621
rect 23584 35544 23612 35584
rect 25317 35581 25329 35615
rect 25363 35581 25375 35615
rect 25593 35615 25651 35621
rect 25593 35612 25605 35615
rect 25317 35575 25375 35581
rect 25516 35584 25605 35612
rect 25332 35544 25360 35575
rect 21324 35516 23060 35544
rect 23216 35516 23612 35544
rect 24320 35516 25360 35544
rect 21324 35504 21330 35516
rect 16960 35448 18552 35476
rect 18601 35479 18659 35485
rect 18601 35445 18613 35479
rect 18647 35476 18659 35479
rect 18874 35476 18880 35488
rect 18647 35448 18880 35476
rect 18647 35445 18659 35448
rect 18601 35439 18659 35445
rect 18874 35436 18880 35448
rect 18932 35436 18938 35488
rect 19334 35476 19340 35488
rect 19295 35448 19340 35476
rect 19334 35436 19340 35448
rect 19392 35436 19398 35488
rect 19981 35479 20039 35485
rect 19981 35445 19993 35479
rect 20027 35476 20039 35479
rect 20346 35476 20352 35488
rect 20027 35448 20352 35476
rect 20027 35445 20039 35448
rect 19981 35439 20039 35445
rect 20346 35436 20352 35448
rect 20404 35436 20410 35488
rect 22370 35436 22376 35488
rect 22428 35476 22434 35488
rect 22557 35479 22615 35485
rect 22557 35476 22569 35479
rect 22428 35448 22569 35476
rect 22428 35436 22434 35448
rect 22557 35445 22569 35448
rect 22603 35445 22615 35479
rect 23032 35476 23060 35516
rect 24320 35476 24348 35516
rect 23032 35448 24348 35476
rect 24397 35479 24455 35485
rect 22557 35439 22615 35445
rect 24397 35445 24409 35479
rect 24443 35476 24455 35479
rect 24762 35476 24768 35488
rect 24443 35448 24768 35476
rect 24443 35445 24455 35448
rect 24397 35439 24455 35445
rect 24762 35436 24768 35448
rect 24820 35436 24826 35488
rect 25222 35436 25228 35488
rect 25280 35476 25286 35488
rect 25516 35476 25544 35584
rect 25593 35581 25605 35584
rect 25639 35581 25651 35615
rect 26436 35612 26464 35643
rect 28000 35612 28028 35720
rect 28902 35708 28908 35720
rect 28960 35708 28966 35760
rect 28077 35683 28135 35689
rect 28077 35649 28089 35683
rect 28123 35649 28135 35683
rect 28077 35643 28135 35649
rect 26436 35584 28028 35612
rect 25593 35575 25651 35581
rect 25774 35504 25780 35556
rect 25832 35544 25838 35556
rect 28092 35544 28120 35643
rect 28442 35640 28448 35692
rect 28500 35680 28506 35692
rect 28721 35683 28779 35689
rect 28721 35680 28733 35683
rect 28500 35652 28733 35680
rect 28500 35640 28506 35652
rect 28721 35649 28733 35652
rect 28767 35649 28779 35683
rect 38010 35680 38016 35692
rect 37971 35652 38016 35680
rect 28721 35643 28779 35649
rect 38010 35640 38016 35652
rect 38068 35640 38074 35692
rect 25832 35516 28120 35544
rect 25832 35504 25838 35516
rect 25280 35448 25544 35476
rect 25280 35436 25286 35448
rect 26326 35436 26332 35488
rect 26384 35476 26390 35488
rect 26513 35479 26571 35485
rect 26513 35476 26525 35479
rect 26384 35448 26525 35476
rect 26384 35436 26390 35448
rect 26513 35445 26525 35448
rect 26559 35445 26571 35479
rect 26513 35439 26571 35445
rect 27338 35436 27344 35488
rect 27396 35476 27402 35488
rect 28169 35479 28227 35485
rect 28169 35476 28181 35479
rect 27396 35448 28181 35476
rect 27396 35436 27402 35448
rect 28169 35445 28181 35448
rect 28215 35445 28227 35479
rect 38194 35476 38200 35488
rect 38155 35448 38200 35476
rect 28169 35439 28227 35445
rect 38194 35436 38200 35448
rect 38252 35436 38258 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 1762 35272 1768 35284
rect 1723 35244 1768 35272
rect 1762 35232 1768 35244
rect 1820 35232 1826 35284
rect 6822 35232 6828 35284
rect 6880 35272 6886 35284
rect 6880 35244 9812 35272
rect 6880 35232 6886 35244
rect 9784 35213 9812 35244
rect 10502 35232 10508 35284
rect 10560 35272 10566 35284
rect 17402 35272 17408 35284
rect 10560 35244 17408 35272
rect 10560 35232 10566 35244
rect 17402 35232 17408 35244
rect 17460 35232 17466 35284
rect 17586 35232 17592 35284
rect 17644 35272 17650 35284
rect 18874 35272 18880 35284
rect 17644 35244 18880 35272
rect 17644 35232 17650 35244
rect 18874 35232 18880 35244
rect 18932 35272 18938 35284
rect 21174 35272 21180 35284
rect 18932 35244 21180 35272
rect 18932 35232 18938 35244
rect 21174 35232 21180 35244
rect 21232 35232 21238 35284
rect 24673 35275 24731 35281
rect 24673 35241 24685 35275
rect 24719 35272 24731 35275
rect 25590 35272 25596 35284
rect 24719 35244 25596 35272
rect 24719 35241 24731 35244
rect 24673 35235 24731 35241
rect 25590 35232 25596 35244
rect 25648 35232 25654 35284
rect 35069 35275 35127 35281
rect 35069 35241 35081 35275
rect 35115 35272 35127 35275
rect 36538 35272 36544 35284
rect 35115 35244 36544 35272
rect 35115 35241 35127 35244
rect 35069 35235 35127 35241
rect 36538 35232 36544 35244
rect 36596 35232 36602 35284
rect 9769 35207 9827 35213
rect 6012 35176 9352 35204
rect 4614 35136 4620 35148
rect 4575 35108 4620 35136
rect 4614 35096 4620 35108
rect 4672 35096 4678 35148
rect 1581 35071 1639 35077
rect 1581 35037 1593 35071
rect 1627 35068 1639 35071
rect 2682 35068 2688 35080
rect 1627 35040 2688 35068
rect 1627 35037 1639 35040
rect 1581 35031 1639 35037
rect 2682 35028 2688 35040
rect 2740 35028 2746 35080
rect 6012 35054 6040 35176
rect 6365 35139 6423 35145
rect 6365 35105 6377 35139
rect 6411 35136 6423 35139
rect 8478 35136 8484 35148
rect 6411 35108 8484 35136
rect 6411 35105 6423 35108
rect 6365 35099 6423 35105
rect 8478 35096 8484 35108
rect 8536 35096 8542 35148
rect 9214 35136 9220 35148
rect 9175 35108 9220 35136
rect 9214 35096 9220 35108
rect 9272 35096 9278 35148
rect 9324 35136 9352 35176
rect 9769 35173 9781 35207
rect 9815 35204 9827 35207
rect 9858 35204 9864 35216
rect 9815 35176 9864 35204
rect 9815 35173 9827 35176
rect 9769 35167 9827 35173
rect 9858 35164 9864 35176
rect 9916 35164 9922 35216
rect 11146 35164 11152 35216
rect 11204 35204 11210 35216
rect 14277 35207 14335 35213
rect 11204 35176 11836 35204
rect 11204 35164 11210 35176
rect 11606 35136 11612 35148
rect 9324 35108 11612 35136
rect 11606 35096 11612 35108
rect 11664 35096 11670 35148
rect 11808 35136 11836 35176
rect 14277 35173 14289 35207
rect 14323 35204 14335 35207
rect 15010 35204 15016 35216
rect 14323 35176 15016 35204
rect 14323 35173 14335 35176
rect 14277 35167 14335 35173
rect 15010 35164 15016 35176
rect 15068 35164 15074 35216
rect 17126 35164 17132 35216
rect 17184 35204 17190 35216
rect 18598 35204 18604 35216
rect 17184 35176 18604 35204
rect 17184 35164 17190 35176
rect 18598 35164 18604 35176
rect 18656 35164 18662 35216
rect 18690 35164 18696 35216
rect 18748 35204 18754 35216
rect 19886 35204 19892 35216
rect 18748 35176 19892 35204
rect 18748 35164 18754 35176
rect 19886 35164 19892 35176
rect 19944 35164 19950 35216
rect 22554 35164 22560 35216
rect 22612 35204 22618 35216
rect 23382 35204 23388 35216
rect 22612 35176 23388 35204
rect 22612 35164 22618 35176
rect 23382 35164 23388 35176
rect 23440 35164 23446 35216
rect 24486 35164 24492 35216
rect 24544 35204 24550 35216
rect 24544 35176 25084 35204
rect 24544 35164 24550 35176
rect 11977 35139 12035 35145
rect 11977 35136 11989 35139
rect 11808 35108 11989 35136
rect 11977 35105 11989 35108
rect 12023 35105 12035 35139
rect 11977 35099 12035 35105
rect 15194 35096 15200 35148
rect 15252 35136 15258 35148
rect 15749 35139 15807 35145
rect 15749 35136 15761 35139
rect 15252 35108 15761 35136
rect 15252 35096 15258 35108
rect 15749 35105 15761 35108
rect 15795 35136 15807 35139
rect 16482 35136 16488 35148
rect 15795 35108 16488 35136
rect 15795 35105 15807 35108
rect 15749 35099 15807 35105
rect 16482 35096 16488 35108
rect 16540 35096 16546 35148
rect 16666 35096 16672 35148
rect 16724 35136 16730 35148
rect 16724 35108 17264 35136
rect 16724 35096 16730 35108
rect 8570 35068 8576 35080
rect 8531 35040 8576 35068
rect 8570 35028 8576 35040
rect 8628 35028 8634 35080
rect 11698 35068 11704 35080
rect 11659 35040 11704 35068
rect 11698 35028 11704 35040
rect 11756 35028 11762 35080
rect 14274 35028 14280 35080
rect 14332 35068 14338 35080
rect 14461 35071 14519 35077
rect 14461 35068 14473 35071
rect 14332 35040 14473 35068
rect 14332 35028 14338 35040
rect 14461 35037 14473 35040
rect 14507 35037 14519 35071
rect 17236 35068 17264 35108
rect 17310 35096 17316 35148
rect 17368 35136 17374 35148
rect 19702 35136 19708 35148
rect 17368 35108 19708 35136
rect 17368 35096 17374 35108
rect 19702 35096 19708 35108
rect 19760 35096 19766 35148
rect 20438 35096 20444 35148
rect 20496 35136 20502 35148
rect 25056 35136 25084 35176
rect 25130 35164 25136 35216
rect 25188 35204 25194 35216
rect 25409 35207 25467 35213
rect 25409 35204 25421 35207
rect 25188 35176 25421 35204
rect 25188 35164 25194 35176
rect 25409 35173 25421 35176
rect 25455 35173 25467 35207
rect 25409 35167 25467 35173
rect 25792 35176 26648 35204
rect 25792 35136 25820 35176
rect 26326 35136 26332 35148
rect 20496 35108 24624 35136
rect 25056 35108 25820 35136
rect 26287 35108 26332 35136
rect 20496 35096 20502 35108
rect 18693 35071 18751 35077
rect 18693 35068 18705 35071
rect 17236 35040 18705 35068
rect 14461 35031 14519 35037
rect 18693 35037 18705 35040
rect 18739 35068 18751 35071
rect 19794 35068 19800 35080
rect 18739 35040 19800 35068
rect 18739 35037 18751 35040
rect 18693 35031 18751 35037
rect 19794 35028 19800 35040
rect 19852 35028 19858 35080
rect 19886 35028 19892 35080
rect 19944 35068 19950 35080
rect 19944 35040 19989 35068
rect 19944 35028 19950 35040
rect 20162 35028 20168 35080
rect 20220 35068 20226 35080
rect 24596 35077 24624 35108
rect 26326 35096 26332 35108
rect 26384 35096 26390 35148
rect 26620 35145 26648 35176
rect 26605 35139 26663 35145
rect 26605 35105 26617 35139
rect 26651 35105 26663 35139
rect 26605 35099 26663 35105
rect 26786 35096 26792 35148
rect 26844 35136 26850 35148
rect 27062 35136 27068 35148
rect 26844 35108 27068 35136
rect 26844 35096 26850 35108
rect 27062 35096 27068 35108
rect 27120 35136 27126 35148
rect 28445 35139 28503 35145
rect 28445 35136 28457 35139
rect 27120 35108 28457 35136
rect 27120 35096 27126 35108
rect 28445 35105 28457 35108
rect 28491 35136 28503 35139
rect 29730 35136 29736 35148
rect 28491 35108 29736 35136
rect 28491 35105 28503 35108
rect 28445 35099 28503 35105
rect 29730 35096 29736 35108
rect 29788 35096 29794 35148
rect 20533 35071 20591 35077
rect 20533 35068 20545 35071
rect 20220 35040 20545 35068
rect 20220 35028 20226 35040
rect 20533 35037 20545 35040
rect 20579 35068 20591 35071
rect 21177 35071 21235 35077
rect 21177 35068 21189 35071
rect 20579 35040 21189 35068
rect 20579 35037 20591 35040
rect 20533 35031 20591 35037
rect 21177 35037 21189 35040
rect 21223 35068 21235 35071
rect 21821 35071 21879 35077
rect 21821 35068 21833 35071
rect 21223 35040 21833 35068
rect 21223 35037 21235 35040
rect 21177 35031 21235 35037
rect 21821 35037 21833 35040
rect 21867 35037 21879 35071
rect 21821 35031 21879 35037
rect 24581 35071 24639 35077
rect 24581 35037 24593 35071
rect 24627 35037 24639 35071
rect 25314 35068 25320 35080
rect 25275 35040 25320 35068
rect 24581 35031 24639 35037
rect 25314 35028 25320 35040
rect 25372 35028 25378 35080
rect 35253 35071 35311 35077
rect 35253 35037 35265 35071
rect 35299 35037 35311 35071
rect 35253 35031 35311 35037
rect 4890 35000 4896 35012
rect 4851 34972 4896 35000
rect 4890 34960 4896 34972
rect 4948 34960 4954 35012
rect 9306 35000 9312 35012
rect 9267 34972 9312 35000
rect 9306 34960 9312 34972
rect 9364 34960 9370 35012
rect 9858 34960 9864 35012
rect 9916 35000 9922 35012
rect 13538 35000 13544 35012
rect 9916 34972 12204 35000
rect 13202 34972 13544 35000
rect 9916 34960 9922 34972
rect 8389 34935 8447 34941
rect 8389 34901 8401 34935
rect 8435 34932 8447 34935
rect 8938 34932 8944 34944
rect 8435 34904 8944 34932
rect 8435 34901 8447 34904
rect 8389 34895 8447 34901
rect 8938 34892 8944 34904
rect 8996 34892 9002 34944
rect 9214 34892 9220 34944
rect 9272 34932 9278 34944
rect 12066 34932 12072 34944
rect 9272 34904 12072 34932
rect 9272 34892 9278 34904
rect 12066 34892 12072 34904
rect 12124 34892 12130 34944
rect 12176 34932 12204 34972
rect 13538 34960 13544 34972
rect 13596 34960 13602 35012
rect 13630 34960 13636 35012
rect 13688 35000 13694 35012
rect 13725 35003 13783 35009
rect 13725 35000 13737 35003
rect 13688 34972 13737 35000
rect 13688 34960 13694 34972
rect 13725 34969 13737 34972
rect 13771 34969 13783 35003
rect 15930 35000 15936 35012
rect 13725 34963 13783 34969
rect 14200 34972 15936 35000
rect 14200 34932 14228 34972
rect 15930 34960 15936 34972
rect 15988 34960 15994 35012
rect 16025 35003 16083 35009
rect 16025 34969 16037 35003
rect 16071 35000 16083 35003
rect 16114 35000 16120 35012
rect 16071 34972 16120 35000
rect 16071 34969 16083 34972
rect 16025 34963 16083 34969
rect 16114 34960 16120 34972
rect 16172 34960 16178 35012
rect 17678 35000 17684 35012
rect 17250 34972 17684 35000
rect 17678 34960 17684 34972
rect 17736 34960 17742 35012
rect 17770 34960 17776 35012
rect 17828 35000 17834 35012
rect 20070 35000 20076 35012
rect 17828 34972 17873 35000
rect 18248 34972 20076 35000
rect 17828 34960 17834 34972
rect 12176 34904 14228 34932
rect 14458 34892 14464 34944
rect 14516 34932 14522 34944
rect 18248 34932 18276 34972
rect 20070 34960 20076 34972
rect 20128 34960 20134 35012
rect 22554 34960 22560 35012
rect 22612 35000 22618 35012
rect 23017 35003 23075 35009
rect 23017 35000 23029 35003
rect 22612 34972 23029 35000
rect 22612 34960 22618 34972
rect 23017 34969 23029 34972
rect 23063 34969 23075 35003
rect 23017 34963 23075 34969
rect 23106 34960 23112 35012
rect 23164 35000 23170 35012
rect 24026 35000 24032 35012
rect 23164 34972 23209 35000
rect 23987 34972 24032 35000
rect 23164 34960 23170 34972
rect 24026 34960 24032 34972
rect 24084 34960 24090 35012
rect 26418 35000 26424 35012
rect 26379 34972 26424 35000
rect 26418 34960 26424 34972
rect 26476 34960 26482 35012
rect 28166 35000 28172 35012
rect 28127 34972 28172 35000
rect 28166 34960 28172 34972
rect 28224 34960 28230 35012
rect 28258 34960 28264 35012
rect 28316 35000 28322 35012
rect 28316 34972 28361 35000
rect 28316 34960 28322 34972
rect 14516 34904 18276 34932
rect 14516 34892 14522 34904
rect 18322 34892 18328 34944
rect 18380 34932 18386 34944
rect 18785 34935 18843 34941
rect 18785 34932 18797 34935
rect 18380 34904 18797 34932
rect 18380 34892 18386 34904
rect 18785 34901 18797 34904
rect 18831 34901 18843 34935
rect 18785 34895 18843 34901
rect 18874 34892 18880 34944
rect 18932 34932 18938 34944
rect 19981 34935 20039 34941
rect 19981 34932 19993 34935
rect 18932 34904 19993 34932
rect 18932 34892 18938 34904
rect 19981 34901 19993 34904
rect 20027 34901 20039 34935
rect 20622 34932 20628 34944
rect 20583 34904 20628 34932
rect 19981 34895 20039 34901
rect 20622 34892 20628 34904
rect 20680 34892 20686 34944
rect 21266 34932 21272 34944
rect 21227 34904 21272 34932
rect 21266 34892 21272 34904
rect 21324 34892 21330 34944
rect 21910 34932 21916 34944
rect 21871 34904 21916 34932
rect 21910 34892 21916 34904
rect 21968 34892 21974 34944
rect 26510 34892 26516 34944
rect 26568 34932 26574 34944
rect 35268 34932 35296 35031
rect 37366 35028 37372 35080
rect 37424 35068 37430 35080
rect 37645 35071 37703 35077
rect 37645 35068 37657 35071
rect 37424 35040 37657 35068
rect 37424 35028 37430 35040
rect 37645 35037 37657 35040
rect 37691 35037 37703 35071
rect 37645 35031 37703 35037
rect 37458 34932 37464 34944
rect 26568 34904 35296 34932
rect 37419 34904 37464 34932
rect 26568 34892 26574 34904
rect 37458 34892 37464 34904
rect 37516 34892 37522 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1581 34731 1639 34737
rect 1581 34697 1593 34731
rect 1627 34728 1639 34731
rect 1627 34700 5580 34728
rect 1627 34697 1639 34700
rect 1581 34691 1639 34697
rect 1762 34592 1768 34604
rect 1723 34564 1768 34592
rect 1762 34552 1768 34564
rect 1820 34552 1826 34604
rect 5552 34601 5580 34700
rect 8570 34688 8576 34740
rect 8628 34728 8634 34740
rect 9585 34731 9643 34737
rect 9585 34728 9597 34731
rect 8628 34700 9597 34728
rect 8628 34688 8634 34700
rect 9585 34697 9597 34700
rect 9631 34697 9643 34731
rect 9585 34691 9643 34697
rect 12360 34700 13492 34728
rect 5629 34663 5687 34669
rect 5629 34629 5641 34663
rect 5675 34660 5687 34663
rect 12360 34660 12388 34700
rect 13354 34660 13360 34672
rect 5675 34632 12388 34660
rect 13202 34632 13360 34660
rect 5675 34629 5687 34632
rect 5629 34623 5687 34629
rect 13354 34620 13360 34632
rect 13412 34620 13418 34672
rect 5537 34595 5595 34601
rect 1578 34484 1584 34536
rect 1636 34524 1642 34536
rect 3237 34527 3295 34533
rect 3237 34524 3249 34527
rect 1636 34496 3249 34524
rect 1636 34484 1642 34496
rect 3237 34493 3249 34496
rect 3283 34493 3295 34527
rect 4632 34524 4660 34578
rect 5537 34561 5549 34595
rect 5583 34561 5595 34595
rect 5537 34555 5595 34561
rect 8662 34552 8668 34604
rect 8720 34592 8726 34604
rect 9769 34595 9827 34601
rect 9769 34592 9781 34595
rect 8720 34564 9781 34592
rect 8720 34552 8726 34564
rect 9769 34561 9781 34564
rect 9815 34592 9827 34595
rect 13464 34592 13492 34700
rect 13538 34688 13544 34740
rect 13596 34728 13602 34740
rect 19337 34731 19395 34737
rect 19337 34728 19349 34731
rect 13596 34700 19349 34728
rect 13596 34688 13602 34700
rect 19337 34697 19349 34700
rect 19383 34697 19395 34731
rect 19337 34691 19395 34697
rect 22094 34688 22100 34740
rect 22152 34728 22158 34740
rect 22152 34700 22324 34728
rect 22152 34688 22158 34700
rect 13722 34620 13728 34672
rect 13780 34660 13786 34672
rect 17678 34660 17684 34672
rect 13780 34632 17684 34660
rect 13780 34620 13786 34632
rect 17678 34620 17684 34632
rect 17736 34620 17742 34672
rect 18046 34620 18052 34672
rect 18104 34660 18110 34672
rect 18690 34660 18696 34672
rect 18104 34632 18696 34660
rect 18104 34620 18110 34632
rect 15562 34592 15568 34604
rect 9815 34564 11560 34592
rect 13464 34564 15568 34592
rect 9815 34561 9827 34564
rect 9769 34555 9827 34561
rect 11330 34524 11336 34536
rect 4632 34496 11336 34524
rect 3237 34487 3295 34493
rect 11330 34484 11336 34496
rect 11388 34484 11394 34536
rect 8202 34456 8208 34468
rect 4908 34428 8208 34456
rect 3500 34391 3558 34397
rect 3500 34357 3512 34391
rect 3546 34388 3558 34391
rect 4908 34388 4936 34428
rect 8202 34416 8208 34428
rect 8260 34416 8266 34468
rect 11532 34456 11560 34564
rect 15562 34552 15568 34564
rect 15620 34552 15626 34604
rect 17313 34595 17371 34601
rect 17313 34561 17325 34595
rect 17359 34561 17371 34595
rect 17313 34555 17371 34561
rect 11698 34524 11704 34536
rect 11659 34496 11704 34524
rect 11698 34484 11704 34496
rect 11756 34484 11762 34536
rect 11977 34527 12035 34533
rect 11977 34524 11989 34527
rect 11808 34496 11989 34524
rect 11808 34456 11836 34496
rect 11977 34493 11989 34496
rect 12023 34524 12035 34527
rect 13725 34527 13783 34533
rect 12023 34496 13584 34524
rect 12023 34493 12035 34496
rect 11977 34487 12035 34493
rect 11532 34428 11836 34456
rect 13556 34456 13584 34496
rect 13725 34493 13737 34527
rect 13771 34524 13783 34527
rect 13906 34524 13912 34536
rect 13771 34496 13912 34524
rect 13771 34493 13783 34496
rect 13725 34487 13783 34493
rect 13906 34484 13912 34496
rect 13964 34484 13970 34536
rect 17328 34524 17356 34555
rect 17402 34552 17408 34604
rect 17460 34592 17466 34604
rect 18616 34601 18644 34632
rect 18690 34620 18696 34632
rect 18748 34620 18754 34672
rect 18966 34620 18972 34672
rect 19024 34660 19030 34672
rect 20165 34663 20223 34669
rect 20165 34660 20177 34663
rect 19024 34632 20177 34660
rect 19024 34620 19030 34632
rect 20165 34629 20177 34632
rect 20211 34629 20223 34663
rect 20165 34623 20223 34629
rect 20254 34620 20260 34672
rect 20312 34660 20318 34672
rect 22296 34660 22324 34700
rect 23382 34688 23388 34740
rect 23440 34728 23446 34740
rect 24029 34731 24087 34737
rect 24029 34728 24041 34731
rect 23440 34700 24041 34728
rect 23440 34688 23446 34700
rect 24029 34697 24041 34700
rect 24075 34697 24087 34731
rect 25130 34728 25136 34740
rect 24029 34691 24087 34697
rect 24412 34700 25136 34728
rect 22465 34663 22523 34669
rect 22465 34660 22477 34663
rect 20312 34632 22094 34660
rect 22296 34632 22477 34660
rect 20312 34620 20318 34632
rect 17957 34595 18015 34601
rect 17460 34564 17505 34592
rect 17460 34552 17466 34564
rect 17957 34561 17969 34595
rect 18003 34592 18015 34595
rect 18601 34595 18659 34601
rect 18003 34564 18184 34592
rect 18003 34561 18015 34564
rect 17957 34555 18015 34561
rect 18156 34536 18184 34564
rect 18601 34561 18613 34595
rect 18647 34561 18659 34595
rect 19242 34592 19248 34604
rect 19203 34564 19248 34592
rect 18601 34555 18659 34561
rect 19242 34552 19248 34564
rect 19300 34552 19306 34604
rect 20073 34595 20131 34601
rect 20073 34561 20085 34595
rect 20119 34592 20131 34595
rect 20530 34592 20536 34604
rect 20119 34564 20536 34592
rect 20119 34561 20131 34564
rect 20073 34555 20131 34561
rect 20530 34552 20536 34564
rect 20588 34592 20594 34604
rect 20717 34595 20775 34601
rect 20717 34592 20729 34595
rect 20588 34564 20729 34592
rect 20588 34552 20594 34564
rect 20717 34561 20729 34564
rect 20763 34561 20775 34595
rect 22066 34592 22094 34632
rect 22465 34629 22477 34632
rect 22511 34629 22523 34663
rect 22465 34623 22523 34629
rect 22557 34663 22615 34669
rect 22557 34629 22569 34663
rect 22603 34660 22615 34663
rect 24412 34660 24440 34700
rect 25130 34688 25136 34700
rect 25188 34688 25194 34740
rect 26510 34728 26516 34740
rect 26471 34700 26516 34728
rect 26510 34688 26516 34700
rect 26568 34688 26574 34740
rect 28166 34688 28172 34740
rect 28224 34728 28230 34740
rect 28353 34731 28411 34737
rect 28353 34728 28365 34731
rect 28224 34700 28365 34728
rect 28224 34688 28230 34700
rect 28353 34697 28365 34700
rect 28399 34697 28411 34731
rect 28353 34691 28411 34697
rect 24673 34663 24731 34669
rect 24673 34660 24685 34663
rect 22603 34632 24440 34660
rect 24504 34632 24685 34660
rect 22603 34629 22615 34632
rect 22557 34623 22615 34629
rect 24504 34604 24532 34632
rect 24673 34629 24685 34632
rect 24719 34629 24731 34663
rect 24673 34623 24731 34629
rect 24762 34620 24768 34672
rect 24820 34660 24826 34672
rect 24820 34632 24865 34660
rect 24820 34620 24826 34632
rect 24946 34620 24952 34672
rect 25004 34660 25010 34672
rect 25317 34663 25375 34669
rect 25317 34660 25329 34663
rect 25004 34632 25329 34660
rect 25004 34620 25010 34632
rect 25317 34629 25329 34632
rect 25363 34660 25375 34663
rect 27338 34660 27344 34672
rect 25363 34632 26464 34660
rect 27299 34632 27344 34660
rect 25363 34629 25375 34632
rect 25317 34623 25375 34629
rect 22066 34590 22140 34592
rect 22278 34590 22284 34604
rect 22066 34564 22284 34590
rect 22112 34562 22284 34564
rect 20717 34555 20775 34561
rect 22278 34552 22284 34562
rect 22336 34552 22342 34604
rect 23934 34592 23940 34604
rect 23400 34564 23612 34592
rect 23895 34564 23940 34592
rect 17328 34496 17448 34524
rect 17310 34456 17316 34468
rect 13556 34428 17316 34456
rect 17310 34416 17316 34428
rect 17368 34416 17374 34468
rect 17420 34456 17448 34496
rect 17494 34484 17500 34536
rect 17552 34524 17558 34536
rect 18049 34527 18107 34533
rect 18049 34524 18061 34527
rect 17552 34496 18061 34524
rect 17552 34484 17558 34496
rect 18049 34493 18061 34496
rect 18095 34493 18107 34527
rect 18049 34487 18107 34493
rect 18138 34484 18144 34536
rect 18196 34524 18202 34536
rect 18690 34524 18696 34536
rect 18196 34496 18289 34524
rect 18651 34496 18696 34524
rect 18196 34484 18202 34496
rect 18690 34484 18696 34496
rect 18748 34484 18754 34536
rect 19334 34484 19340 34536
rect 19392 34524 19398 34536
rect 20809 34527 20867 34533
rect 20809 34524 20821 34527
rect 19392 34496 20821 34524
rect 19392 34484 19398 34496
rect 20809 34493 20821 34496
rect 20855 34493 20867 34527
rect 20809 34487 20867 34493
rect 20898 34484 20904 34536
rect 20956 34524 20962 34536
rect 23400 34524 23428 34564
rect 20956 34496 22140 34524
rect 20956 34484 20962 34496
rect 18156 34456 18184 34484
rect 19518 34456 19524 34468
rect 17420 34428 19524 34456
rect 19518 34416 19524 34428
rect 19576 34416 19582 34468
rect 20714 34416 20720 34468
rect 20772 34456 20778 34468
rect 21174 34456 21180 34468
rect 20772 34428 21180 34456
rect 20772 34416 20778 34428
rect 21174 34416 21180 34428
rect 21232 34416 21238 34468
rect 3546 34360 4936 34388
rect 3546 34357 3558 34360
rect 3500 34351 3558 34357
rect 4982 34348 4988 34400
rect 5040 34388 5046 34400
rect 5040 34360 5085 34388
rect 5040 34348 5046 34360
rect 6914 34348 6920 34400
rect 6972 34388 6978 34400
rect 11790 34388 11796 34400
rect 6972 34360 11796 34388
rect 6972 34348 6978 34360
rect 11790 34348 11796 34360
rect 11848 34348 11854 34400
rect 14366 34348 14372 34400
rect 14424 34388 14430 34400
rect 18138 34388 18144 34400
rect 14424 34360 18144 34388
rect 14424 34348 14430 34360
rect 18138 34348 18144 34360
rect 18196 34348 18202 34400
rect 18230 34348 18236 34400
rect 18288 34388 18294 34400
rect 21266 34388 21272 34400
rect 18288 34360 21272 34388
rect 18288 34348 18294 34360
rect 21266 34348 21272 34360
rect 21324 34388 21330 34400
rect 22002 34388 22008 34400
rect 21324 34360 22008 34388
rect 21324 34348 21330 34360
rect 22002 34348 22008 34360
rect 22060 34348 22066 34400
rect 22112 34388 22140 34496
rect 22388 34496 23428 34524
rect 23477 34527 23535 34533
rect 22388 34388 22416 34496
rect 23477 34493 23489 34527
rect 23523 34493 23535 34527
rect 23584 34524 23612 34564
rect 23934 34552 23940 34564
rect 23992 34552 23998 34604
rect 24486 34552 24492 34604
rect 24544 34552 24550 34604
rect 26436 34601 26464 34632
rect 27338 34620 27344 34632
rect 27396 34620 27402 34672
rect 26421 34595 26479 34601
rect 26421 34561 26433 34595
rect 26467 34561 26479 34595
rect 26421 34555 26479 34561
rect 36630 34552 36636 34604
rect 36688 34592 36694 34604
rect 38013 34595 38071 34601
rect 38013 34592 38025 34595
rect 36688 34564 38025 34592
rect 36688 34552 36694 34564
rect 38013 34561 38025 34564
rect 38059 34561 38071 34595
rect 38013 34555 38071 34561
rect 27249 34527 27307 34533
rect 27249 34524 27261 34527
rect 23584 34512 24716 34524
rect 24780 34512 27261 34524
rect 23584 34496 27261 34512
rect 23477 34487 23535 34493
rect 23382 34416 23388 34468
rect 23440 34456 23446 34468
rect 23492 34456 23520 34487
rect 24688 34484 24808 34496
rect 27249 34493 27261 34496
rect 27295 34493 27307 34527
rect 27890 34524 27896 34536
rect 27851 34496 27896 34524
rect 27249 34487 27307 34493
rect 27890 34484 27896 34496
rect 27948 34484 27954 34536
rect 28350 34456 28356 34468
rect 23440 34428 28356 34456
rect 23440 34416 23446 34428
rect 28350 34416 28356 34428
rect 28408 34416 28414 34468
rect 22112 34360 22416 34388
rect 24118 34348 24124 34400
rect 24176 34388 24182 34400
rect 28718 34388 28724 34400
rect 24176 34360 28724 34388
rect 24176 34348 24182 34360
rect 28718 34348 28724 34360
rect 28776 34348 28782 34400
rect 38194 34388 38200 34400
rect 38155 34360 38200 34388
rect 38194 34348 38200 34360
rect 38252 34348 38258 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 3234 34144 3240 34196
rect 3292 34184 3298 34196
rect 6914 34184 6920 34196
rect 3292 34156 6920 34184
rect 3292 34144 3298 34156
rect 6914 34144 6920 34156
rect 6972 34144 6978 34196
rect 7024 34156 12020 34184
rect 5442 34008 5448 34060
rect 5500 34048 5506 34060
rect 5629 34051 5687 34057
rect 5629 34048 5641 34051
rect 5500 34020 5641 34048
rect 5500 34008 5506 34020
rect 5629 34017 5641 34020
rect 5675 34017 5687 34051
rect 5629 34011 5687 34017
rect 1581 33983 1639 33989
rect 1581 33949 1593 33983
rect 1627 33980 1639 33983
rect 2406 33980 2412 33992
rect 1627 33952 2412 33980
rect 1627 33949 1639 33952
rect 1581 33943 1639 33949
rect 2406 33940 2412 33952
rect 2464 33940 2470 33992
rect 2498 33940 2504 33992
rect 2556 33980 2562 33992
rect 2556 33952 2601 33980
rect 7024 33966 7052 34156
rect 9122 34008 9128 34060
rect 9180 34048 9186 34060
rect 9401 34051 9459 34057
rect 9401 34048 9413 34051
rect 9180 34020 9413 34048
rect 9180 34008 9186 34020
rect 9401 34017 9413 34020
rect 9447 34017 9459 34051
rect 9674 34048 9680 34060
rect 9635 34020 9680 34048
rect 9401 34011 9459 34017
rect 9674 34008 9680 34020
rect 9732 34008 9738 34060
rect 11698 34008 11704 34060
rect 11756 34048 11762 34060
rect 11874 34051 11932 34057
rect 11874 34048 11886 34051
rect 11756 34020 11886 34048
rect 11756 34008 11762 34020
rect 11874 34017 11886 34020
rect 11920 34017 11932 34051
rect 11992 34048 12020 34156
rect 12158 34144 12164 34196
rect 12216 34184 12222 34196
rect 13722 34184 13728 34196
rect 12216 34156 13728 34184
rect 12216 34144 12222 34156
rect 13722 34144 13728 34156
rect 13780 34144 13786 34196
rect 15286 34144 15292 34196
rect 15344 34184 15350 34196
rect 16850 34184 16856 34196
rect 15344 34156 16856 34184
rect 15344 34144 15350 34156
rect 16850 34144 16856 34156
rect 16908 34144 16914 34196
rect 17126 34144 17132 34196
rect 17184 34184 17190 34196
rect 18230 34184 18236 34196
rect 17184 34156 18236 34184
rect 17184 34144 17190 34156
rect 18230 34144 18236 34156
rect 18288 34144 18294 34196
rect 18506 34144 18512 34196
rect 18564 34184 18570 34196
rect 18785 34187 18843 34193
rect 18785 34184 18797 34187
rect 18564 34156 18797 34184
rect 18564 34144 18570 34156
rect 18785 34153 18797 34156
rect 18831 34153 18843 34187
rect 18785 34147 18843 34153
rect 19058 34144 19064 34196
rect 19116 34184 19122 34196
rect 20254 34184 20260 34196
rect 19116 34156 20260 34184
rect 19116 34144 19122 34156
rect 20254 34144 20260 34156
rect 20312 34144 20318 34196
rect 22097 34187 22155 34193
rect 22097 34153 22109 34187
rect 22143 34184 22155 34187
rect 28258 34184 28264 34196
rect 22143 34156 28264 34184
rect 22143 34153 22155 34156
rect 22097 34147 22155 34153
rect 28258 34144 28264 34156
rect 28316 34144 28322 34196
rect 36630 34184 36636 34196
rect 36591 34156 36636 34184
rect 36630 34144 36636 34156
rect 36688 34144 36694 34196
rect 16574 34076 16580 34128
rect 16632 34116 16638 34128
rect 20622 34116 20628 34128
rect 16632 34088 20628 34116
rect 16632 34076 16638 34088
rect 20622 34076 20628 34088
rect 20680 34076 20686 34128
rect 22738 34076 22744 34128
rect 22796 34116 22802 34128
rect 23474 34116 23480 34128
rect 22796 34088 23480 34116
rect 22796 34076 22802 34088
rect 23474 34076 23480 34088
rect 23532 34116 23538 34128
rect 24026 34116 24032 34128
rect 23532 34088 24032 34116
rect 23532 34076 23538 34088
rect 24026 34076 24032 34088
rect 24084 34076 24090 34128
rect 27801 34119 27859 34125
rect 27801 34116 27813 34119
rect 24504 34088 27813 34116
rect 24504 34060 24532 34088
rect 27801 34085 27813 34088
rect 27847 34085 27859 34119
rect 27801 34079 27859 34085
rect 14918 34048 14924 34060
rect 11992 34020 14924 34048
rect 11874 34011 11932 34017
rect 14918 34008 14924 34020
rect 14976 34008 14982 34060
rect 15194 34008 15200 34060
rect 15252 34048 15258 34060
rect 15289 34051 15347 34057
rect 15289 34048 15301 34051
rect 15252 34020 15301 34048
rect 15252 34008 15258 34020
rect 15289 34017 15301 34020
rect 15335 34017 15347 34051
rect 15289 34011 15347 34017
rect 17126 34008 17132 34060
rect 17184 34048 17190 34060
rect 17313 34051 17371 34057
rect 17313 34048 17325 34051
rect 17184 34020 17325 34048
rect 17184 34008 17190 34020
rect 17313 34017 17325 34020
rect 17359 34017 17371 34051
rect 17313 34011 17371 34017
rect 17402 34008 17408 34060
rect 17460 34048 17466 34060
rect 23014 34048 23020 34060
rect 17460 34020 23020 34048
rect 17460 34008 17466 34020
rect 23014 34008 23020 34020
rect 23072 34008 23078 34060
rect 23385 34051 23443 34057
rect 23385 34017 23397 34051
rect 23431 34048 23443 34051
rect 24486 34048 24492 34060
rect 23431 34020 24492 34048
rect 23431 34017 23443 34020
rect 23385 34011 23443 34017
rect 24486 34008 24492 34020
rect 24544 34008 24550 34060
rect 27246 34048 27252 34060
rect 27207 34020 27252 34048
rect 27246 34008 27252 34020
rect 27304 34008 27310 34060
rect 2556 33940 2562 33952
rect 13262 33940 13268 33992
rect 13320 33940 13326 33992
rect 18046 33980 18052 33992
rect 18007 33952 18052 33980
rect 18046 33940 18052 33952
rect 18104 33940 18110 33992
rect 18138 33940 18144 33992
rect 18196 33980 18202 33992
rect 18693 33983 18751 33989
rect 18196 33952 18241 33980
rect 18196 33940 18202 33952
rect 18693 33949 18705 33983
rect 18739 33980 18751 33983
rect 19426 33980 19432 33992
rect 18739 33952 19432 33980
rect 18739 33949 18751 33952
rect 18693 33943 18751 33949
rect 19426 33940 19432 33952
rect 19484 33940 19490 33992
rect 19518 33940 19524 33992
rect 19576 33980 19582 33992
rect 20622 33980 20628 33992
rect 19576 33952 20628 33980
rect 19576 33940 19582 33952
rect 20622 33940 20628 33952
rect 20680 33940 20686 33992
rect 20809 33983 20867 33989
rect 20809 33949 20821 33983
rect 20855 33949 20867 33983
rect 20809 33943 20867 33949
rect 5902 33912 5908 33924
rect 5863 33884 5908 33912
rect 5902 33872 5908 33884
rect 5960 33872 5966 33924
rect 12161 33915 12219 33921
rect 10902 33884 12112 33912
rect 1762 33844 1768 33856
rect 1723 33816 1768 33844
rect 1762 33804 1768 33816
rect 1820 33804 1826 33856
rect 1854 33804 1860 33856
rect 1912 33844 1918 33856
rect 2317 33847 2375 33853
rect 2317 33844 2329 33847
rect 1912 33816 2329 33844
rect 1912 33804 1918 33816
rect 2317 33813 2329 33816
rect 2363 33813 2375 33847
rect 2317 33807 2375 33813
rect 7377 33847 7435 33853
rect 7377 33813 7389 33847
rect 7423 33844 7435 33847
rect 9582 33844 9588 33856
rect 7423 33816 9588 33844
rect 7423 33813 7435 33816
rect 7377 33807 7435 33813
rect 9582 33804 9588 33816
rect 9640 33804 9646 33856
rect 11146 33844 11152 33856
rect 11107 33816 11152 33844
rect 11146 33804 11152 33816
rect 11204 33804 11210 33856
rect 12084 33844 12112 33884
rect 12161 33881 12173 33915
rect 12207 33912 12219 33915
rect 12250 33912 12256 33924
rect 12207 33884 12256 33912
rect 12207 33881 12219 33884
rect 12161 33875 12219 33881
rect 12250 33872 12256 33884
rect 12308 33872 12314 33924
rect 15565 33915 15623 33921
rect 13464 33884 15424 33912
rect 13464 33844 13492 33884
rect 12084 33816 13492 33844
rect 13633 33847 13691 33853
rect 13633 33813 13645 33847
rect 13679 33844 13691 33847
rect 15286 33844 15292 33856
rect 13679 33816 15292 33844
rect 13679 33813 13691 33816
rect 13633 33807 13691 33813
rect 15286 33804 15292 33816
rect 15344 33804 15350 33856
rect 15396 33844 15424 33884
rect 15565 33881 15577 33915
rect 15611 33912 15623 33915
rect 15838 33912 15844 33924
rect 15611 33884 15844 33912
rect 15611 33881 15623 33884
rect 15565 33875 15623 33881
rect 15838 33872 15844 33884
rect 15896 33872 15902 33924
rect 16942 33912 16948 33924
rect 16790 33884 16948 33912
rect 16942 33872 16948 33884
rect 17000 33872 17006 33924
rect 17034 33872 17040 33924
rect 17092 33912 17098 33924
rect 19334 33912 19340 33924
rect 17092 33884 19340 33912
rect 17092 33872 17098 33884
rect 19334 33872 19340 33884
rect 19392 33872 19398 33924
rect 20824 33912 20852 33943
rect 21082 33940 21088 33992
rect 21140 33980 21146 33992
rect 22005 33983 22063 33989
rect 22005 33980 22017 33983
rect 21140 33952 22017 33980
rect 21140 33940 21146 33952
rect 22005 33949 22017 33952
rect 22051 33949 22063 33983
rect 22005 33943 22063 33949
rect 23566 33940 23572 33992
rect 23624 33980 23630 33992
rect 23624 33952 24256 33980
rect 23624 33940 23630 33952
rect 22738 33912 22744 33924
rect 19444 33884 20852 33912
rect 22699 33884 22744 33912
rect 16574 33844 16580 33856
rect 15396 33816 16580 33844
rect 16574 33804 16580 33816
rect 16632 33804 16638 33856
rect 19242 33804 19248 33856
rect 19300 33844 19306 33856
rect 19444 33844 19472 33884
rect 22738 33872 22744 33884
rect 22796 33872 22802 33924
rect 22833 33915 22891 33921
rect 22833 33881 22845 33915
rect 22879 33912 22891 33915
rect 24228 33912 24256 33952
rect 24302 33940 24308 33992
rect 24360 33980 24366 33992
rect 25225 33983 25283 33989
rect 25225 33980 25237 33983
rect 24360 33952 25237 33980
rect 24360 33940 24366 33952
rect 25225 33949 25237 33952
rect 25271 33949 25283 33983
rect 28350 33980 28356 33992
rect 28311 33952 28356 33980
rect 25225 33943 25283 33949
rect 28350 33940 28356 33952
rect 28408 33940 28414 33992
rect 36814 33980 36820 33992
rect 36775 33952 36820 33980
rect 36814 33940 36820 33952
rect 36872 33940 36878 33992
rect 27341 33915 27399 33921
rect 22879 33884 24072 33912
rect 24228 33884 27292 33912
rect 22879 33881 22891 33884
rect 22833 33875 22891 33881
rect 19300 33816 19472 33844
rect 19613 33847 19671 33853
rect 19300 33804 19306 33816
rect 19613 33813 19625 33847
rect 19659 33844 19671 33847
rect 19978 33844 19984 33856
rect 19659 33816 19984 33844
rect 19659 33813 19671 33816
rect 19613 33807 19671 33813
rect 19978 33804 19984 33816
rect 20036 33804 20042 33856
rect 20165 33847 20223 33853
rect 20165 33813 20177 33847
rect 20211 33844 20223 33847
rect 20438 33844 20444 33856
rect 20211 33816 20444 33844
rect 20211 33813 20223 33816
rect 20165 33807 20223 33813
rect 20438 33804 20444 33816
rect 20496 33804 20502 33856
rect 20898 33844 20904 33856
rect 20859 33816 20904 33844
rect 20898 33804 20904 33816
rect 20956 33804 20962 33856
rect 24044 33844 24072 33884
rect 25317 33847 25375 33853
rect 25317 33844 25329 33847
rect 24044 33816 25329 33844
rect 25317 33813 25329 33816
rect 25363 33813 25375 33847
rect 27264 33844 27292 33884
rect 27341 33881 27353 33915
rect 27387 33912 27399 33915
rect 27706 33912 27712 33924
rect 27387 33884 27712 33912
rect 27387 33881 27399 33884
rect 27341 33875 27399 33881
rect 27706 33872 27712 33884
rect 27764 33872 27770 33924
rect 29638 33912 29644 33924
rect 28276 33884 29644 33912
rect 28276 33844 28304 33884
rect 29638 33872 29644 33884
rect 29696 33872 29702 33924
rect 28442 33844 28448 33856
rect 27264 33816 28304 33844
rect 28403 33816 28448 33844
rect 25317 33807 25375 33813
rect 28442 33804 28448 33816
rect 28500 33804 28506 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 5442 33640 5448 33652
rect 2056 33612 5448 33640
rect 1578 33464 1584 33516
rect 1636 33504 1642 33516
rect 2056 33513 2084 33612
rect 4062 33572 4068 33584
rect 3542 33544 4068 33572
rect 4062 33532 4068 33544
rect 4120 33532 4126 33584
rect 4264 33513 4292 33612
rect 5442 33600 5448 33612
rect 5500 33600 5506 33652
rect 5902 33600 5908 33652
rect 5960 33640 5966 33652
rect 5997 33643 6055 33649
rect 5997 33640 6009 33643
rect 5960 33612 6009 33640
rect 5960 33600 5966 33612
rect 5997 33609 6009 33612
rect 6043 33609 6055 33643
rect 5997 33603 6055 33609
rect 7484 33612 9168 33640
rect 7484 33516 7512 33612
rect 9140 33584 9168 33612
rect 13262 33600 13268 33652
rect 13320 33640 13326 33652
rect 17034 33640 17040 33652
rect 13320 33612 17040 33640
rect 13320 33600 13326 33612
rect 17034 33600 17040 33612
rect 17092 33600 17098 33652
rect 23566 33640 23572 33652
rect 20548 33612 23572 33640
rect 9122 33532 9128 33584
rect 9180 33572 9186 33584
rect 10413 33575 10471 33581
rect 10413 33572 10425 33575
rect 9180 33544 10425 33572
rect 9180 33532 9186 33544
rect 10413 33541 10425 33544
rect 10459 33541 10471 33575
rect 10413 33535 10471 33541
rect 11146 33532 11152 33584
rect 11204 33572 11210 33584
rect 12989 33575 13047 33581
rect 11204 33544 12283 33572
rect 11204 33532 11210 33544
rect 2041 33507 2099 33513
rect 2041 33504 2053 33507
rect 1636 33476 2053 33504
rect 1636 33464 1642 33476
rect 2041 33473 2053 33476
rect 2087 33473 2099 33507
rect 2041 33467 2099 33473
rect 4249 33507 4307 33513
rect 4249 33473 4261 33507
rect 4295 33473 4307 33507
rect 7466 33504 7472 33516
rect 4249 33467 4307 33473
rect 2317 33439 2375 33445
rect 2317 33405 2329 33439
rect 2363 33436 2375 33439
rect 3789 33439 3847 33445
rect 2363 33408 3740 33436
rect 2363 33405 2375 33408
rect 2317 33399 2375 33405
rect 3712 33300 3740 33408
rect 3789 33405 3801 33439
rect 3835 33436 3847 33439
rect 4525 33439 4583 33445
rect 4525 33436 4537 33439
rect 3835 33408 4537 33436
rect 3835 33405 3847 33408
rect 3789 33399 3847 33405
rect 4525 33405 4537 33408
rect 4571 33436 4583 33439
rect 5258 33436 5264 33448
rect 4571 33408 5264 33436
rect 4571 33405 4583 33408
rect 4525 33399 4583 33405
rect 5258 33396 5264 33408
rect 5316 33396 5322 33448
rect 4982 33300 4988 33312
rect 3712 33272 4988 33300
rect 4982 33260 4988 33272
rect 5040 33260 5046 33312
rect 5644 33300 5672 33490
rect 7379 33476 7472 33504
rect 7466 33464 7472 33476
rect 7524 33464 7530 33516
rect 7745 33439 7803 33445
rect 7745 33405 7757 33439
rect 7791 33436 7803 33439
rect 8478 33436 8484 33448
rect 7791 33408 8484 33436
rect 7791 33405 7803 33408
rect 7745 33399 7803 33405
rect 8478 33396 8484 33408
rect 8536 33436 8542 33448
rect 8864 33436 8892 33490
rect 9030 33464 9036 33516
rect 9088 33504 9094 33516
rect 9490 33504 9496 33516
rect 9088 33476 9496 33504
rect 9088 33464 9094 33476
rect 9490 33464 9496 33476
rect 9548 33464 9554 33516
rect 9677 33507 9735 33513
rect 9677 33473 9689 33507
rect 9723 33504 9735 33507
rect 11974 33504 11980 33516
rect 9723 33476 11980 33504
rect 9723 33473 9735 33476
rect 9677 33467 9735 33473
rect 11974 33464 11980 33476
rect 12032 33464 12038 33516
rect 11606 33436 11612 33448
rect 8536 33408 8800 33436
rect 8864 33408 11612 33436
rect 8536 33396 8542 33408
rect 8772 33368 8800 33408
rect 11606 33396 11612 33408
rect 11664 33396 11670 33448
rect 9030 33368 9036 33380
rect 8772 33340 9036 33368
rect 9030 33328 9036 33340
rect 9088 33328 9094 33380
rect 11882 33368 11888 33380
rect 9140 33340 11888 33368
rect 9140 33300 9168 33340
rect 11882 33328 11888 33340
rect 11940 33328 11946 33380
rect 12255 33368 12283 33544
rect 12989 33541 13001 33575
rect 13035 33572 13047 33575
rect 13078 33572 13084 33584
rect 13035 33544 13084 33572
rect 13035 33541 13047 33544
rect 12989 33535 13047 33541
rect 13078 33532 13084 33544
rect 13136 33532 13142 33584
rect 17402 33572 17408 33584
rect 14214 33544 17408 33572
rect 17402 33532 17408 33544
rect 17460 33532 17466 33584
rect 18782 33572 18788 33584
rect 18354 33544 18788 33572
rect 18782 33532 18788 33544
rect 18840 33532 18846 33584
rect 20070 33572 20076 33584
rect 19168 33544 20076 33572
rect 19168 33516 19196 33544
rect 20070 33532 20076 33544
rect 20128 33532 20134 33584
rect 20438 33572 20444 33584
rect 20399 33544 20444 33572
rect 20438 33532 20444 33544
rect 20496 33532 20502 33584
rect 20548 33581 20576 33612
rect 23566 33600 23572 33612
rect 23624 33600 23630 33652
rect 23842 33640 23848 33652
rect 23803 33612 23848 33640
rect 23842 33600 23848 33612
rect 23900 33600 23906 33652
rect 25130 33640 25136 33652
rect 25091 33612 25136 33640
rect 25130 33600 25136 33612
rect 25188 33600 25194 33652
rect 25777 33643 25835 33649
rect 25777 33609 25789 33643
rect 25823 33640 25835 33643
rect 26418 33640 26424 33652
rect 25823 33612 26424 33640
rect 25823 33609 25835 33612
rect 25777 33603 25835 33609
rect 26418 33600 26424 33612
rect 26476 33600 26482 33652
rect 26528 33612 27476 33640
rect 20533 33575 20591 33581
rect 20533 33541 20545 33575
rect 20579 33541 20591 33575
rect 20533 33535 20591 33541
rect 22186 33532 22192 33584
rect 22244 33572 22250 33584
rect 22833 33575 22891 33581
rect 22833 33572 22845 33575
rect 22244 33544 22845 33572
rect 22244 33532 22250 33544
rect 22833 33541 22845 33544
rect 22879 33541 22891 33575
rect 22833 33535 22891 33541
rect 23753 33575 23811 33581
rect 23753 33541 23765 33575
rect 23799 33572 23811 33575
rect 24118 33572 24124 33584
rect 23799 33544 24124 33572
rect 23799 33541 23811 33544
rect 23753 33535 23811 33541
rect 24118 33532 24124 33544
rect 24176 33532 24182 33584
rect 26528 33572 26556 33612
rect 27338 33572 27344 33584
rect 24412 33544 26556 33572
rect 27299 33544 27344 33572
rect 15194 33464 15200 33516
rect 15252 33504 15258 33516
rect 16482 33504 16488 33516
rect 15252 33476 16488 33504
rect 15252 33464 15258 33476
rect 16482 33464 16488 33476
rect 16540 33504 16546 33516
rect 16853 33507 16911 33513
rect 16853 33504 16865 33507
rect 16540 33476 16865 33504
rect 16540 33464 16546 33476
rect 16853 33473 16865 33476
rect 16899 33473 16911 33507
rect 16853 33467 16911 33473
rect 19150 33464 19156 33516
rect 19208 33464 19214 33516
rect 19426 33464 19432 33516
rect 19484 33504 19490 33516
rect 19521 33507 19579 33513
rect 19521 33504 19533 33507
rect 19484 33476 19533 33504
rect 19484 33464 19490 33476
rect 19521 33473 19533 33476
rect 19567 33473 19579 33507
rect 22738 33504 22744 33516
rect 22699 33476 22744 33504
rect 19521 33467 19579 33473
rect 22738 33464 22744 33476
rect 22796 33464 22802 33516
rect 24412 33513 24440 33544
rect 27338 33532 27344 33544
rect 27396 33532 27402 33584
rect 27448 33572 27476 33612
rect 27706 33600 27712 33652
rect 27764 33640 27770 33652
rect 28445 33643 28503 33649
rect 28445 33640 28457 33643
rect 27764 33612 28457 33640
rect 27764 33600 27770 33612
rect 28445 33609 28457 33612
rect 28491 33609 28503 33643
rect 28445 33603 28503 33609
rect 28534 33572 28540 33584
rect 27448 33544 28540 33572
rect 28534 33532 28540 33544
rect 28592 33532 28598 33584
rect 29822 33572 29828 33584
rect 29012 33544 29828 33572
rect 24397 33507 24455 33513
rect 24397 33473 24409 33507
rect 24443 33473 24455 33507
rect 25038 33504 25044 33516
rect 24999 33476 25044 33504
rect 24397 33467 24455 33473
rect 25038 33464 25044 33476
rect 25096 33464 25102 33516
rect 25685 33507 25743 33513
rect 25685 33473 25697 33507
rect 25731 33504 25743 33507
rect 25958 33504 25964 33516
rect 25731 33476 25964 33504
rect 25731 33473 25743 33476
rect 25685 33467 25743 33473
rect 25958 33464 25964 33476
rect 26016 33464 26022 33516
rect 29012 33513 29040 33544
rect 29822 33532 29828 33544
rect 29880 33532 29886 33584
rect 28353 33507 28411 33513
rect 28353 33473 28365 33507
rect 28399 33473 28411 33507
rect 28353 33467 28411 33473
rect 28997 33507 29055 33513
rect 28997 33473 29009 33507
rect 29043 33473 29055 33507
rect 29638 33504 29644 33516
rect 29599 33476 29644 33504
rect 28997 33467 29055 33473
rect 12342 33396 12348 33448
rect 12400 33436 12406 33448
rect 12713 33439 12771 33445
rect 12713 33436 12725 33439
rect 12400 33408 12725 33436
rect 12400 33396 12406 33408
rect 12713 33405 12725 33408
rect 12759 33405 12771 33439
rect 12713 33399 12771 33405
rect 14737 33439 14795 33445
rect 14737 33405 14749 33439
rect 14783 33436 14795 33439
rect 15838 33436 15844 33448
rect 14783 33408 15844 33436
rect 14783 33405 14795 33408
rect 14737 33399 14795 33405
rect 15838 33396 15844 33408
rect 15896 33396 15902 33448
rect 17129 33439 17187 33445
rect 17129 33405 17141 33439
rect 17175 33436 17187 33439
rect 17586 33436 17592 33448
rect 17175 33408 17592 33436
rect 17175 33405 17187 33408
rect 17129 33399 17187 33405
rect 17586 33396 17592 33408
rect 17644 33396 17650 33448
rect 17678 33396 17684 33448
rect 17736 33436 17742 33448
rect 21453 33439 21511 33445
rect 17736 33408 21220 33436
rect 17736 33396 17742 33408
rect 21082 33368 21088 33380
rect 12255 33340 12848 33368
rect 5644 33272 9168 33300
rect 9217 33303 9275 33309
rect 9217 33269 9229 33303
rect 9263 33300 9275 33303
rect 12158 33300 12164 33312
rect 9263 33272 12164 33300
rect 9263 33269 9275 33272
rect 9217 33263 9275 33269
rect 12158 33260 12164 33272
rect 12216 33260 12222 33312
rect 12820 33300 12848 33340
rect 18156 33340 21088 33368
rect 18156 33300 18184 33340
rect 21082 33328 21088 33340
rect 21140 33328 21146 33380
rect 21192 33368 21220 33408
rect 21453 33405 21465 33439
rect 21499 33436 21511 33439
rect 27246 33436 27252 33448
rect 21499 33408 22324 33436
rect 27207 33408 27252 33436
rect 21499 33405 21511 33408
rect 21453 33399 21511 33405
rect 22296 33368 22324 33408
rect 27246 33396 27252 33408
rect 27304 33396 27310 33448
rect 27890 33436 27896 33448
rect 27851 33408 27896 33436
rect 27890 33396 27896 33408
rect 27948 33396 27954 33448
rect 26142 33368 26148 33380
rect 21192 33340 22094 33368
rect 22296 33340 26148 33368
rect 12820 33272 18184 33300
rect 18506 33260 18512 33312
rect 18564 33300 18570 33312
rect 18601 33303 18659 33309
rect 18601 33300 18613 33303
rect 18564 33272 18613 33300
rect 18564 33260 18570 33272
rect 18601 33269 18613 33272
rect 18647 33269 18659 33303
rect 18601 33263 18659 33269
rect 19334 33260 19340 33312
rect 19392 33300 19398 33312
rect 19613 33303 19671 33309
rect 19613 33300 19625 33303
rect 19392 33272 19625 33300
rect 19392 33260 19398 33272
rect 19613 33269 19625 33272
rect 19659 33269 19671 33303
rect 19613 33263 19671 33269
rect 19702 33260 19708 33312
rect 19760 33300 19766 33312
rect 21818 33300 21824 33312
rect 19760 33272 21824 33300
rect 19760 33260 19766 33272
rect 21818 33260 21824 33272
rect 21876 33260 21882 33312
rect 22066 33300 22094 33340
rect 26142 33328 26148 33340
rect 26200 33328 26206 33380
rect 26234 33328 26240 33380
rect 26292 33368 26298 33380
rect 28368 33368 28396 33467
rect 29638 33464 29644 33476
rect 29696 33464 29702 33516
rect 26292 33340 28396 33368
rect 26292 33328 26298 33340
rect 23474 33300 23480 33312
rect 22066 33272 23480 33300
rect 23474 33260 23480 33272
rect 23532 33260 23538 33312
rect 23934 33260 23940 33312
rect 23992 33300 23998 33312
rect 24489 33303 24547 33309
rect 24489 33300 24501 33303
rect 23992 33272 24501 33300
rect 23992 33260 23998 33272
rect 24489 33269 24501 33272
rect 24535 33269 24547 33303
rect 29086 33300 29092 33312
rect 29047 33272 29092 33300
rect 24489 33263 24547 33269
rect 29086 33260 29092 33272
rect 29144 33260 29150 33312
rect 29178 33260 29184 33312
rect 29236 33300 29242 33312
rect 29733 33303 29791 33309
rect 29733 33300 29745 33303
rect 29236 33272 29745 33300
rect 29236 33260 29242 33272
rect 29733 33269 29745 33272
rect 29779 33269 29791 33303
rect 29733 33263 29791 33269
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 2041 33099 2099 33105
rect 2041 33065 2053 33099
rect 2087 33096 2099 33099
rect 2498 33096 2504 33108
rect 2087 33068 2504 33096
rect 2087 33065 2099 33068
rect 2041 33059 2099 33065
rect 2498 33056 2504 33068
rect 2556 33056 2562 33108
rect 8481 33099 8539 33105
rect 8481 33065 8493 33099
rect 8527 33096 8539 33099
rect 9674 33096 9680 33108
rect 8527 33068 9680 33096
rect 8527 33065 8539 33068
rect 8481 33059 8539 33065
rect 9674 33056 9680 33068
rect 9732 33056 9738 33108
rect 11054 33056 11060 33108
rect 11112 33056 11118 33108
rect 12250 33056 12256 33108
rect 12308 33096 12314 33108
rect 14734 33096 14740 33108
rect 12308 33068 14740 33096
rect 12308 33056 12314 33068
rect 14734 33056 14740 33068
rect 14792 33056 14798 33108
rect 17678 33056 17684 33108
rect 17736 33096 17742 33108
rect 19150 33096 19156 33108
rect 17736 33068 19156 33096
rect 17736 33056 17742 33068
rect 19150 33056 19156 33068
rect 19208 33056 19214 33108
rect 25317 33099 25375 33105
rect 19720 33068 25268 33096
rect 11072 33028 11100 33056
rect 8128 33000 11100 33028
rect 6733 32963 6791 32969
rect 6733 32929 6745 32963
rect 6779 32960 6791 32963
rect 7466 32960 7472 32972
rect 6779 32932 7472 32960
rect 6779 32929 6791 32932
rect 6733 32923 6791 32929
rect 7466 32920 7472 32932
rect 7524 32920 7530 32972
rect 2041 32895 2099 32901
rect 2041 32861 2053 32895
rect 2087 32892 2099 32895
rect 5810 32892 5816 32904
rect 2087 32864 5816 32892
rect 2087 32861 2099 32864
rect 2041 32855 2099 32861
rect 5810 32852 5816 32864
rect 5868 32852 5874 32904
rect 8128 32878 8156 33000
rect 13446 32988 13452 33040
rect 13504 33028 13510 33040
rect 14918 33028 14924 33040
rect 13504 33000 14924 33028
rect 13504 32988 13510 33000
rect 14918 32988 14924 33000
rect 14976 32988 14982 33040
rect 19518 33028 19524 33040
rect 17144 33000 19524 33028
rect 15194 32960 15200 32972
rect 9646 32932 15056 32960
rect 15155 32932 15200 32960
rect 9646 32892 9674 32932
rect 8404 32864 9674 32892
rect 7009 32827 7067 32833
rect 7009 32793 7021 32827
rect 7055 32793 7067 32827
rect 7009 32787 7067 32793
rect 7024 32756 7052 32787
rect 8404 32756 8432 32864
rect 10778 32852 10784 32904
rect 10836 32892 10842 32904
rect 10965 32895 11023 32901
rect 10965 32892 10977 32895
rect 10836 32864 10977 32892
rect 10836 32852 10842 32864
rect 10965 32861 10977 32864
rect 11011 32861 11023 32895
rect 10965 32855 11023 32861
rect 10870 32784 10876 32836
rect 10928 32824 10934 32836
rect 11241 32827 11299 32833
rect 11241 32824 11253 32827
rect 10928 32796 11253 32824
rect 10928 32784 10934 32796
rect 11241 32793 11253 32796
rect 11287 32793 11299 32827
rect 12618 32824 12624 32836
rect 12466 32796 12624 32824
rect 11241 32787 11299 32793
rect 7024 32728 8432 32756
rect 11256 32756 11284 32787
rect 12618 32784 12624 32796
rect 12676 32784 12682 32836
rect 12986 32824 12992 32836
rect 12947 32796 12992 32824
rect 12986 32784 12992 32796
rect 13044 32784 13050 32836
rect 14461 32827 14519 32833
rect 14461 32793 14473 32827
rect 14507 32793 14519 32827
rect 14461 32787 14519 32793
rect 11882 32756 11888 32768
rect 11256 32728 11888 32756
rect 11882 32716 11888 32728
rect 11940 32716 11946 32768
rect 11974 32716 11980 32768
rect 12032 32756 12038 32768
rect 14476 32756 14504 32787
rect 12032 32728 14504 32756
rect 15028 32756 15056 32932
rect 15194 32920 15200 32932
rect 15252 32960 15258 32972
rect 15841 32963 15899 32969
rect 15841 32960 15853 32963
rect 15252 32932 15853 32960
rect 15252 32920 15258 32932
rect 15841 32929 15853 32932
rect 15887 32929 15899 32963
rect 15841 32923 15899 32929
rect 16206 32920 16212 32972
rect 16264 32960 16270 32972
rect 17144 32960 17172 33000
rect 19518 32988 19524 33000
rect 19576 32988 19582 33040
rect 16264 32932 17172 32960
rect 16264 32920 16270 32932
rect 17310 32920 17316 32972
rect 17368 32960 17374 32972
rect 19610 32960 19616 32972
rect 17368 32932 19616 32960
rect 17368 32920 17374 32932
rect 19610 32920 19616 32932
rect 19668 32920 19674 32972
rect 17402 32852 17408 32904
rect 17460 32892 17466 32904
rect 19720 32892 19748 33068
rect 19886 33028 19892 33040
rect 19847 33000 19892 33028
rect 19886 32988 19892 33000
rect 19944 32988 19950 33040
rect 23566 32988 23572 33040
rect 23624 33028 23630 33040
rect 24673 33031 24731 33037
rect 24673 33028 24685 33031
rect 23624 33000 24685 33028
rect 23624 32988 23630 33000
rect 24673 32997 24685 33000
rect 24719 32997 24731 33031
rect 24673 32991 24731 32997
rect 19978 32920 19984 32972
rect 20036 32960 20042 32972
rect 20254 32960 20260 32972
rect 20036 32932 20260 32960
rect 20036 32920 20042 32932
rect 20254 32920 20260 32932
rect 20312 32920 20318 32972
rect 20530 32960 20536 32972
rect 20491 32932 20536 32960
rect 20530 32920 20536 32932
rect 20588 32920 20594 32972
rect 21269 32963 21327 32969
rect 21269 32929 21281 32963
rect 21315 32960 21327 32963
rect 21450 32960 21456 32972
rect 21315 32932 21456 32960
rect 21315 32929 21327 32932
rect 21269 32923 21327 32929
rect 21450 32920 21456 32932
rect 21508 32920 21514 32972
rect 23124 32932 25176 32960
rect 17460 32864 19748 32892
rect 19797 32895 19855 32901
rect 17460 32852 17466 32864
rect 19797 32861 19809 32895
rect 19843 32892 19855 32895
rect 20070 32892 20076 32904
rect 19843 32864 20076 32892
rect 19843 32861 19855 32864
rect 19797 32855 19855 32861
rect 20070 32852 20076 32864
rect 20128 32892 20134 32904
rect 20441 32895 20499 32901
rect 20441 32892 20453 32895
rect 20128 32864 20453 32892
rect 20128 32852 20134 32864
rect 20441 32861 20453 32864
rect 20487 32861 20499 32895
rect 23124 32892 23152 32932
rect 20441 32855 20499 32861
rect 22296 32864 23152 32892
rect 15286 32784 15292 32836
rect 15344 32824 15350 32836
rect 16117 32827 16175 32833
rect 16117 32824 16129 32827
rect 15344 32796 16129 32824
rect 15344 32784 15350 32796
rect 16117 32793 16129 32796
rect 16163 32824 16175 32827
rect 16390 32824 16396 32836
rect 16163 32796 16396 32824
rect 16163 32793 16175 32796
rect 16117 32787 16175 32793
rect 16390 32784 16396 32796
rect 16448 32784 16454 32836
rect 17954 32824 17960 32836
rect 17342 32796 17960 32824
rect 17954 32784 17960 32796
rect 18012 32784 18018 32836
rect 18598 32784 18604 32836
rect 18656 32824 18662 32836
rect 20530 32824 20536 32836
rect 18656 32796 20536 32824
rect 18656 32784 18662 32796
rect 20530 32784 20536 32796
rect 20588 32784 20594 32836
rect 22296 32833 22324 32864
rect 23198 32852 23204 32904
rect 23256 32892 23262 32904
rect 23293 32895 23351 32901
rect 23293 32892 23305 32895
rect 23256 32864 23305 32892
rect 23256 32852 23262 32864
rect 23293 32861 23305 32864
rect 23339 32861 23351 32895
rect 24578 32892 24584 32904
rect 24539 32864 24584 32892
rect 23293 32855 23351 32861
rect 24578 32852 24584 32864
rect 24636 32892 24642 32904
rect 25038 32892 25044 32904
rect 24636 32864 25044 32892
rect 24636 32852 24642 32864
rect 25038 32852 25044 32864
rect 25096 32852 25102 32904
rect 21361 32827 21419 32833
rect 21361 32793 21373 32827
rect 21407 32793 21419 32827
rect 21361 32787 21419 32793
rect 22281 32827 22339 32833
rect 22281 32793 22293 32827
rect 22327 32793 22339 32827
rect 23842 32824 23848 32836
rect 22281 32787 22339 32793
rect 23032 32796 23848 32824
rect 17126 32756 17132 32768
rect 15028 32728 17132 32756
rect 12032 32716 12038 32728
rect 17126 32716 17132 32728
rect 17184 32716 17190 32768
rect 17586 32756 17592 32768
rect 17547 32728 17592 32756
rect 17586 32716 17592 32728
rect 17644 32716 17650 32768
rect 17770 32716 17776 32768
rect 17828 32756 17834 32768
rect 21082 32756 21088 32768
rect 17828 32728 21088 32756
rect 17828 32716 17834 32728
rect 21082 32716 21088 32728
rect 21140 32716 21146 32768
rect 21376 32756 21404 32787
rect 23032 32756 23060 32796
rect 23842 32784 23848 32796
rect 23900 32784 23906 32836
rect 25148 32824 25176 32932
rect 25240 32901 25268 33068
rect 25317 33065 25329 33099
rect 25363 33096 25375 33099
rect 27338 33096 27344 33108
rect 25363 33068 27344 33096
rect 25363 33065 25375 33068
rect 25317 33059 25375 33065
rect 27338 33056 27344 33068
rect 27396 33056 27402 33108
rect 26142 32920 26148 32972
rect 26200 32960 26206 32972
rect 26421 32963 26479 32969
rect 26421 32960 26433 32963
rect 26200 32932 26433 32960
rect 26200 32920 26206 32932
rect 26421 32929 26433 32932
rect 26467 32929 26479 32963
rect 26421 32923 26479 32929
rect 27709 32963 27767 32969
rect 27709 32929 27721 32963
rect 27755 32960 27767 32963
rect 29086 32960 29092 32972
rect 27755 32932 29092 32960
rect 27755 32929 27767 32932
rect 27709 32923 27767 32929
rect 29086 32920 29092 32932
rect 29144 32920 29150 32972
rect 25225 32895 25283 32901
rect 25225 32861 25237 32895
rect 25271 32861 25283 32895
rect 25225 32855 25283 32861
rect 34146 32852 34152 32904
rect 34204 32892 34210 32904
rect 38013 32895 38071 32901
rect 38013 32892 38025 32895
rect 34204 32864 38025 32892
rect 34204 32852 34210 32864
rect 38013 32861 38025 32864
rect 38059 32861 38071 32895
rect 38013 32855 38071 32861
rect 25498 32824 25504 32836
rect 25148 32796 25504 32824
rect 25498 32784 25504 32796
rect 25556 32784 25562 32836
rect 26142 32824 26148 32836
rect 26103 32796 26148 32824
rect 26142 32784 26148 32796
rect 26200 32784 26206 32836
rect 26237 32827 26295 32833
rect 26237 32793 26249 32827
rect 26283 32793 26295 32827
rect 26237 32787 26295 32793
rect 21376 32728 23060 32756
rect 23385 32759 23443 32765
rect 23385 32725 23397 32759
rect 23431 32756 23443 32759
rect 26050 32756 26056 32768
rect 23431 32728 26056 32756
rect 23431 32725 23443 32728
rect 23385 32719 23443 32725
rect 26050 32716 26056 32728
rect 26108 32716 26114 32768
rect 26252 32756 26280 32787
rect 27338 32784 27344 32836
rect 27396 32824 27402 32836
rect 27801 32827 27859 32833
rect 27801 32824 27813 32827
rect 27396 32796 27813 32824
rect 27396 32784 27402 32796
rect 27801 32793 27813 32796
rect 27847 32793 27859 32827
rect 27801 32787 27859 32793
rect 27982 32784 27988 32836
rect 28040 32824 28046 32836
rect 28721 32827 28779 32833
rect 28721 32824 28733 32827
rect 28040 32796 28733 32824
rect 28040 32784 28046 32796
rect 28721 32793 28733 32796
rect 28767 32793 28779 32827
rect 28721 32787 28779 32793
rect 28442 32756 28448 32768
rect 26252 32728 28448 32756
rect 28442 32716 28448 32728
rect 28500 32716 28506 32768
rect 38194 32756 38200 32768
rect 38155 32728 38200 32756
rect 38194 32716 38200 32728
rect 38252 32716 38258 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 10502 32512 10508 32564
rect 10560 32552 10566 32564
rect 20254 32552 20260 32564
rect 10560 32524 20260 32552
rect 10560 32512 10566 32524
rect 20254 32512 20260 32524
rect 20312 32512 20318 32564
rect 20622 32512 20628 32564
rect 20680 32552 20686 32564
rect 22186 32552 22192 32564
rect 20680 32524 22192 32552
rect 20680 32512 20686 32524
rect 22186 32512 22192 32524
rect 22244 32512 22250 32564
rect 34514 32552 34520 32564
rect 26252 32524 34520 32552
rect 5442 32444 5448 32496
rect 5500 32484 5506 32496
rect 7285 32487 7343 32493
rect 7285 32484 7297 32487
rect 5500 32456 7297 32484
rect 5500 32444 5506 32456
rect 7285 32453 7297 32456
rect 7331 32453 7343 32487
rect 7285 32447 7343 32453
rect 9582 32444 9588 32496
rect 9640 32484 9646 32496
rect 9677 32487 9735 32493
rect 9677 32484 9689 32487
rect 9640 32456 9689 32484
rect 9640 32444 9646 32456
rect 9677 32453 9689 32456
rect 9723 32453 9735 32487
rect 11974 32484 11980 32496
rect 11935 32456 11980 32484
rect 9677 32447 9735 32453
rect 11974 32444 11980 32456
rect 12032 32444 12038 32496
rect 14734 32484 14740 32496
rect 14695 32456 14740 32484
rect 14734 32444 14740 32456
rect 14792 32444 14798 32496
rect 16758 32484 16764 32496
rect 15962 32456 16764 32484
rect 16758 32444 16764 32456
rect 16816 32444 16822 32496
rect 17034 32444 17040 32496
rect 17092 32484 17098 32496
rect 17402 32484 17408 32496
rect 17092 32456 17408 32484
rect 17092 32444 17098 32456
rect 17402 32444 17408 32456
rect 17460 32444 17466 32496
rect 19610 32444 19616 32496
rect 19668 32484 19674 32496
rect 19958 32487 20016 32493
rect 19958 32484 19970 32487
rect 19668 32456 19970 32484
rect 19668 32444 19674 32456
rect 19958 32453 19970 32456
rect 20004 32453 20016 32487
rect 23198 32484 23204 32496
rect 19958 32447 20016 32453
rect 20732 32456 23204 32484
rect 1670 32416 1676 32428
rect 1631 32388 1676 32416
rect 1670 32376 1676 32388
rect 1728 32376 1734 32428
rect 6546 32416 6552 32428
rect 6507 32388 6552 32416
rect 6546 32376 6552 32388
rect 6604 32376 6610 32428
rect 9122 32376 9128 32428
rect 9180 32416 9186 32428
rect 9401 32419 9459 32425
rect 9401 32416 9413 32419
rect 9180 32388 9413 32416
rect 9180 32376 9186 32388
rect 9401 32385 9413 32388
rect 9447 32385 9459 32419
rect 13814 32416 13820 32428
rect 10810 32388 13820 32416
rect 9401 32379 9459 32385
rect 13814 32376 13820 32388
rect 13872 32376 13878 32428
rect 14458 32416 14464 32428
rect 14419 32388 14464 32416
rect 14458 32376 14464 32388
rect 14516 32376 14522 32428
rect 16482 32376 16488 32428
rect 16540 32416 16546 32428
rect 16853 32419 16911 32425
rect 16853 32416 16865 32419
rect 16540 32388 16865 32416
rect 16540 32376 16546 32388
rect 16853 32385 16865 32388
rect 16899 32385 16911 32419
rect 18262 32388 19012 32416
rect 16853 32379 16911 32385
rect 9674 32308 9680 32360
rect 9732 32348 9738 32360
rect 9732 32320 10732 32348
rect 9732 32308 9738 32320
rect 1857 32283 1915 32289
rect 1857 32249 1869 32283
rect 1903 32280 1915 32283
rect 2222 32280 2228 32292
rect 1903 32252 2228 32280
rect 1903 32249 1915 32252
rect 1857 32243 1915 32249
rect 2222 32240 2228 32252
rect 2280 32240 2286 32292
rect 10704 32280 10732 32320
rect 11698 32308 11704 32360
rect 11756 32348 11762 32360
rect 11882 32348 11888 32360
rect 11756 32320 11888 32348
rect 11756 32308 11762 32320
rect 11882 32308 11888 32320
rect 11940 32348 11946 32360
rect 12342 32348 12348 32360
rect 11940 32320 12348 32348
rect 11940 32308 11946 32320
rect 12342 32308 12348 32320
rect 12400 32348 12406 32360
rect 12713 32351 12771 32357
rect 12713 32348 12725 32351
rect 12400 32320 12725 32348
rect 12400 32308 12406 32320
rect 12713 32317 12725 32320
rect 12759 32317 12771 32351
rect 16206 32348 16212 32360
rect 12713 32311 12771 32317
rect 14568 32320 16212 32348
rect 14568 32280 14596 32320
rect 16206 32308 16212 32320
rect 16264 32308 16270 32360
rect 16298 32308 16304 32360
rect 16356 32348 16362 32360
rect 17129 32351 17187 32357
rect 17129 32348 17141 32351
rect 16356 32320 17141 32348
rect 16356 32308 16362 32320
rect 17129 32317 17141 32320
rect 17175 32317 17187 32351
rect 17129 32311 17187 32317
rect 17218 32308 17224 32360
rect 17276 32348 17282 32360
rect 17770 32348 17776 32360
rect 17276 32320 17776 32348
rect 17276 32308 17282 32320
rect 17770 32308 17776 32320
rect 17828 32308 17834 32360
rect 18984 32348 19012 32388
rect 19058 32376 19064 32428
rect 19116 32416 19122 32428
rect 19153 32419 19211 32425
rect 19153 32416 19165 32419
rect 19116 32388 19165 32416
rect 19116 32376 19122 32388
rect 19153 32385 19165 32388
rect 19199 32416 19211 32419
rect 19242 32416 19248 32428
rect 19199 32388 19248 32416
rect 19199 32385 19211 32388
rect 19153 32379 19211 32385
rect 19242 32376 19248 32388
rect 19300 32376 19306 32428
rect 19610 32348 19616 32360
rect 18984 32320 19616 32348
rect 19610 32308 19616 32320
rect 19668 32308 19674 32360
rect 19886 32348 19892 32360
rect 19847 32320 19892 32348
rect 19886 32308 19892 32320
rect 19944 32308 19950 32360
rect 20254 32348 20260 32360
rect 20215 32320 20260 32348
rect 20254 32308 20260 32320
rect 20312 32308 20318 32360
rect 20732 32280 20760 32456
rect 23198 32444 23204 32456
rect 23256 32444 23262 32496
rect 23566 32484 23572 32496
rect 23527 32456 23572 32484
rect 23566 32444 23572 32456
rect 23624 32444 23630 32496
rect 25130 32484 25136 32496
rect 25091 32456 25136 32484
rect 25130 32444 25136 32456
rect 25188 32444 25194 32496
rect 22002 32416 22008 32428
rect 21963 32388 22008 32416
rect 22002 32376 22008 32388
rect 22060 32376 22066 32428
rect 22833 32419 22891 32425
rect 22833 32385 22845 32419
rect 22879 32416 22891 32419
rect 23290 32416 23296 32428
rect 22879 32388 23296 32416
rect 22879 32385 22891 32388
rect 22833 32379 22891 32385
rect 23290 32376 23296 32388
rect 23348 32376 23354 32428
rect 26252 32425 26280 32524
rect 34514 32512 34520 32524
rect 34572 32512 34578 32564
rect 27246 32484 27252 32496
rect 27207 32456 27252 32484
rect 27246 32444 27252 32456
rect 27304 32444 27310 32496
rect 28997 32487 29055 32493
rect 28997 32484 29009 32487
rect 27816 32456 29009 32484
rect 26237 32419 26295 32425
rect 26237 32385 26249 32419
rect 26283 32385 26295 32419
rect 26237 32379 26295 32385
rect 27157 32419 27215 32425
rect 27157 32385 27169 32419
rect 27203 32416 27215 32419
rect 27430 32416 27436 32428
rect 27203 32388 27436 32416
rect 27203 32385 27215 32388
rect 27157 32379 27215 32385
rect 27430 32376 27436 32388
rect 27488 32376 27494 32428
rect 22462 32308 22468 32360
rect 22520 32348 22526 32360
rect 23477 32351 23535 32357
rect 22520 32320 22692 32348
rect 22520 32308 22526 32320
rect 22664 32289 22692 32320
rect 23477 32317 23489 32351
rect 23523 32348 23535 32351
rect 23934 32348 23940 32360
rect 23523 32320 23940 32348
rect 23523 32317 23535 32320
rect 23477 32311 23535 32317
rect 23934 32308 23940 32320
rect 23992 32308 23998 32360
rect 24029 32351 24087 32357
rect 24029 32317 24041 32351
rect 24075 32317 24087 32351
rect 24029 32311 24087 32317
rect 22097 32283 22155 32289
rect 22097 32280 22109 32283
rect 10704 32252 14596 32280
rect 18616 32252 20760 32280
rect 20824 32252 22109 32280
rect 5534 32172 5540 32224
rect 5592 32212 5598 32224
rect 11054 32212 11060 32224
rect 5592 32184 11060 32212
rect 5592 32172 5598 32184
rect 11054 32172 11060 32184
rect 11112 32172 11118 32224
rect 11149 32215 11207 32221
rect 11149 32181 11161 32215
rect 11195 32212 11207 32215
rect 14366 32212 14372 32224
rect 11195 32184 14372 32212
rect 11195 32181 11207 32184
rect 11149 32175 11207 32181
rect 14366 32172 14372 32184
rect 14424 32172 14430 32224
rect 14458 32172 14464 32224
rect 14516 32212 14522 32224
rect 15838 32212 15844 32224
rect 14516 32184 15844 32212
rect 14516 32172 14522 32184
rect 15838 32172 15844 32184
rect 15896 32172 15902 32224
rect 16206 32212 16212 32224
rect 16167 32184 16212 32212
rect 16206 32172 16212 32184
rect 16264 32172 16270 32224
rect 16390 32172 16396 32224
rect 16448 32212 16454 32224
rect 16942 32212 16948 32224
rect 16448 32184 16948 32212
rect 16448 32172 16454 32184
rect 16942 32172 16948 32184
rect 17000 32172 17006 32224
rect 17126 32172 17132 32224
rect 17184 32212 17190 32224
rect 18616 32221 18644 32252
rect 20824 32224 20852 32252
rect 22097 32249 22109 32252
rect 22143 32249 22155 32283
rect 22097 32243 22155 32249
rect 22649 32283 22707 32289
rect 22649 32249 22661 32283
rect 22695 32249 22707 32283
rect 22649 32243 22707 32249
rect 23014 32240 23020 32292
rect 23072 32280 23078 32292
rect 24044 32280 24072 32311
rect 24854 32308 24860 32360
rect 24912 32348 24918 32360
rect 25041 32351 25099 32357
rect 25041 32348 25053 32351
rect 24912 32320 25053 32348
rect 24912 32308 24918 32320
rect 25041 32317 25053 32320
rect 25087 32317 25099 32351
rect 25041 32311 25099 32317
rect 26142 32308 26148 32360
rect 26200 32348 26206 32360
rect 27816 32357 27844 32456
rect 28997 32453 29009 32456
rect 29043 32453 29055 32487
rect 28997 32447 29055 32453
rect 28718 32376 28724 32428
rect 28776 32416 28782 32428
rect 28905 32419 28963 32425
rect 28905 32416 28917 32419
rect 28776 32388 28917 32416
rect 28776 32376 28782 32388
rect 28905 32385 28917 32388
rect 28951 32385 28963 32419
rect 28905 32379 28963 32385
rect 35434 32376 35440 32428
rect 35492 32416 35498 32428
rect 38013 32419 38071 32425
rect 38013 32416 38025 32419
rect 35492 32388 38025 32416
rect 35492 32376 35498 32388
rect 38013 32385 38025 32388
rect 38059 32385 38071 32419
rect 38013 32379 38071 32385
rect 27801 32351 27859 32357
rect 27801 32348 27813 32351
rect 26200 32320 27813 32348
rect 26200 32308 26206 32320
rect 27801 32317 27813 32320
rect 27847 32317 27859 32351
rect 27801 32311 27859 32317
rect 27985 32351 28043 32357
rect 27985 32317 27997 32351
rect 28031 32348 28043 32351
rect 28994 32348 29000 32360
rect 28031 32320 29000 32348
rect 28031 32317 28043 32320
rect 27985 32311 28043 32317
rect 28994 32308 29000 32320
rect 29052 32308 29058 32360
rect 25406 32280 25412 32292
rect 23072 32252 24072 32280
rect 25148 32252 25412 32280
rect 23072 32240 23078 32252
rect 18601 32215 18659 32221
rect 18601 32212 18613 32215
rect 17184 32184 18613 32212
rect 17184 32172 17190 32184
rect 18601 32181 18613 32184
rect 18647 32181 18659 32215
rect 19242 32212 19248 32224
rect 19203 32184 19248 32212
rect 18601 32175 18659 32181
rect 19242 32172 19248 32184
rect 19300 32172 19306 32224
rect 19886 32172 19892 32224
rect 19944 32212 19950 32224
rect 20806 32212 20812 32224
rect 19944 32184 20812 32212
rect 19944 32172 19950 32184
rect 20806 32172 20812 32184
rect 20864 32172 20870 32224
rect 21082 32172 21088 32224
rect 21140 32212 21146 32224
rect 25148 32212 25176 32252
rect 25406 32240 25412 32252
rect 25464 32240 25470 32292
rect 25593 32283 25651 32289
rect 25593 32249 25605 32283
rect 25639 32280 25651 32283
rect 29914 32280 29920 32292
rect 25639 32252 29920 32280
rect 25639 32249 25651 32252
rect 25593 32243 25651 32249
rect 29914 32240 29920 32252
rect 29972 32240 29978 32292
rect 21140 32184 25176 32212
rect 21140 32172 21146 32184
rect 25222 32172 25228 32224
rect 25280 32212 25286 32224
rect 26329 32215 26387 32221
rect 26329 32212 26341 32215
rect 25280 32184 26341 32212
rect 25280 32172 25286 32184
rect 26329 32181 26341 32184
rect 26375 32181 26387 32215
rect 26329 32175 26387 32181
rect 26694 32172 26700 32224
rect 26752 32212 26758 32224
rect 27062 32212 27068 32224
rect 26752 32184 27068 32212
rect 26752 32172 26758 32184
rect 27062 32172 27068 32184
rect 27120 32172 27126 32224
rect 28074 32172 28080 32224
rect 28132 32212 28138 32224
rect 28169 32215 28227 32221
rect 28169 32212 28181 32215
rect 28132 32184 28181 32212
rect 28132 32172 28138 32184
rect 28169 32181 28181 32184
rect 28215 32181 28227 32215
rect 38194 32212 38200 32224
rect 38155 32184 38200 32212
rect 28169 32175 28227 32181
rect 38194 32172 38200 32184
rect 38252 32172 38258 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 6086 32008 6092 32020
rect 5276 31980 6092 32008
rect 5276 31881 5304 31980
rect 6086 31968 6092 31980
rect 6144 31968 6150 32020
rect 6656 31980 11928 32008
rect 5261 31875 5319 31881
rect 5261 31841 5273 31875
rect 5307 31841 5319 31875
rect 5534 31872 5540 31884
rect 5495 31844 5540 31872
rect 5261 31835 5319 31841
rect 5534 31832 5540 31844
rect 5592 31832 5598 31884
rect 1581 31807 1639 31813
rect 1581 31773 1593 31807
rect 1627 31804 1639 31807
rect 1854 31804 1860 31816
rect 1627 31776 1860 31804
rect 1627 31773 1639 31776
rect 1581 31767 1639 31773
rect 1854 31764 1860 31776
rect 1912 31764 1918 31816
rect 2314 31804 2320 31816
rect 2275 31776 2320 31804
rect 2314 31764 2320 31776
rect 2372 31764 2378 31816
rect 2406 31764 2412 31816
rect 2464 31804 2470 31816
rect 2464 31776 2509 31804
rect 6656 31790 6684 31980
rect 7006 31940 7012 31952
rect 6967 31912 7012 31940
rect 7006 31900 7012 31912
rect 7064 31900 7070 31952
rect 9122 31872 9128 31884
rect 9083 31844 9128 31872
rect 9122 31832 9128 31844
rect 9180 31832 9186 31884
rect 9401 31875 9459 31881
rect 9401 31841 9413 31875
rect 9447 31872 9459 31875
rect 11790 31872 11796 31884
rect 9447 31844 11796 31872
rect 9447 31841 9459 31844
rect 9401 31835 9459 31841
rect 11790 31832 11796 31844
rect 11848 31832 11854 31884
rect 11900 31872 11928 31980
rect 13814 31968 13820 32020
rect 13872 32008 13878 32020
rect 15378 32008 15384 32020
rect 13872 31980 15384 32008
rect 13872 31968 13878 31980
rect 15378 31968 15384 31980
rect 15436 31968 15442 32020
rect 15930 31968 15936 32020
rect 15988 32008 15994 32020
rect 19334 32008 19340 32020
rect 15988 31980 19340 32008
rect 15988 31968 15994 31980
rect 19334 31968 19340 31980
rect 19392 31968 19398 32020
rect 19444 31980 25084 32008
rect 18506 31940 18512 31952
rect 17328 31912 18512 31940
rect 13814 31872 13820 31884
rect 11900 31844 13820 31872
rect 13814 31832 13820 31844
rect 13872 31832 13878 31884
rect 14550 31832 14556 31884
rect 14608 31872 14614 31884
rect 14734 31872 14740 31884
rect 14608 31844 14740 31872
rect 14608 31832 14614 31844
rect 14734 31832 14740 31844
rect 14792 31832 14798 31884
rect 16025 31875 16083 31881
rect 16025 31841 16037 31875
rect 16071 31872 16083 31875
rect 16390 31872 16396 31884
rect 16071 31844 16396 31872
rect 16071 31841 16083 31844
rect 16025 31835 16083 31841
rect 16390 31832 16396 31844
rect 16448 31832 16454 31884
rect 16666 31832 16672 31884
rect 16724 31872 16730 31884
rect 17328 31872 17356 31912
rect 18506 31900 18512 31912
rect 18564 31900 18570 31952
rect 17770 31872 17776 31884
rect 16724 31844 17356 31872
rect 17731 31844 17776 31872
rect 16724 31832 16730 31844
rect 17770 31832 17776 31844
rect 17828 31832 17834 31884
rect 17862 31832 17868 31884
rect 17920 31872 17926 31884
rect 19444 31872 19472 31980
rect 20254 31940 20260 31952
rect 19536 31912 20260 31940
rect 19536 31881 19564 31912
rect 20254 31900 20260 31912
rect 20312 31900 20318 31952
rect 24946 31940 24952 31952
rect 20456 31912 24952 31940
rect 17920 31844 19472 31872
rect 19521 31875 19579 31881
rect 17920 31832 17926 31844
rect 19521 31841 19533 31875
rect 19567 31841 19579 31875
rect 19521 31835 19579 31841
rect 20165 31875 20223 31881
rect 20165 31841 20177 31875
rect 20211 31872 20223 31875
rect 20456 31872 20484 31912
rect 23308 31881 23336 31912
rect 24946 31900 24952 31912
rect 25004 31900 25010 31952
rect 20211 31844 20484 31872
rect 23293 31875 23351 31881
rect 20211 31841 20223 31844
rect 20165 31835 20223 31841
rect 23293 31841 23305 31875
rect 23339 31841 23351 31875
rect 25056 31872 25084 31980
rect 25130 31968 25136 32020
rect 25188 32008 25194 32020
rect 27617 32011 27675 32017
rect 27617 32008 27629 32011
rect 25188 31980 27629 32008
rect 25188 31968 25194 31980
rect 27617 31977 27629 31980
rect 27663 31977 27675 32011
rect 28994 32008 29000 32020
rect 28955 31980 29000 32008
rect 27617 31971 27675 31977
rect 28994 31968 29000 31980
rect 29052 31968 29058 32020
rect 25406 31900 25412 31952
rect 25464 31940 25470 31952
rect 25464 31912 26924 31940
rect 25464 31900 25470 31912
rect 25682 31872 25688 31884
rect 25056 31844 25688 31872
rect 23293 31835 23351 31841
rect 25682 31832 25688 31844
rect 25740 31832 25746 31884
rect 25866 31832 25872 31884
rect 25924 31881 26096 31884
rect 25924 31875 26111 31881
rect 25924 31856 26065 31875
rect 25924 31832 25930 31856
rect 26053 31841 26065 31856
rect 26099 31841 26111 31875
rect 26053 31835 26111 31841
rect 2464 31764 2470 31776
rect 10502 31764 10508 31816
rect 10560 31764 10566 31816
rect 10778 31764 10784 31816
rect 10836 31804 10842 31816
rect 11882 31804 11888 31816
rect 10836 31776 11888 31804
rect 10836 31764 10842 31776
rect 11882 31764 11888 31776
rect 11940 31804 11946 31816
rect 11977 31807 12035 31813
rect 11977 31804 11989 31807
rect 11940 31776 11989 31804
rect 11940 31764 11946 31776
rect 11977 31773 11989 31776
rect 12023 31773 12035 31807
rect 17678 31804 17684 31816
rect 17434 31776 17684 31804
rect 11977 31767 12035 31773
rect 17678 31764 17684 31776
rect 17736 31764 17742 31816
rect 18693 31807 18751 31813
rect 18693 31773 18705 31807
rect 18739 31804 18751 31807
rect 19058 31804 19064 31816
rect 18739 31776 19064 31804
rect 18739 31773 18751 31776
rect 18693 31767 18751 31773
rect 19058 31764 19064 31776
rect 19116 31764 19122 31816
rect 20530 31764 20536 31816
rect 20588 31798 20594 31816
rect 20625 31807 20683 31813
rect 20625 31798 20637 31807
rect 20588 31773 20637 31798
rect 20671 31773 20683 31807
rect 20588 31770 20683 31773
rect 20588 31764 20594 31770
rect 20625 31767 20683 31770
rect 25317 31807 25375 31813
rect 25317 31773 25329 31807
rect 25363 31804 25375 31807
rect 25774 31804 25780 31816
rect 25363 31776 25780 31804
rect 25363 31773 25375 31776
rect 25317 31767 25375 31773
rect 25774 31764 25780 31776
rect 25832 31764 25838 31816
rect 26896 31804 26924 31912
rect 27062 31832 27068 31884
rect 27120 31872 27126 31884
rect 27120 31844 27165 31872
rect 27120 31832 27126 31844
rect 27614 31832 27620 31884
rect 27672 31872 27678 31884
rect 27672 31844 28948 31872
rect 27672 31832 27678 31844
rect 27525 31807 27583 31813
rect 27525 31804 27537 31807
rect 26896 31776 27537 31804
rect 27525 31773 27537 31776
rect 27571 31804 27583 31807
rect 28258 31804 28264 31816
rect 27571 31776 28264 31804
rect 27571 31773 27583 31776
rect 27525 31767 27583 31773
rect 28258 31764 28264 31776
rect 28316 31764 28322 31816
rect 28920 31813 28948 31844
rect 28905 31807 28963 31813
rect 28905 31773 28917 31807
rect 28951 31804 28963 31807
rect 30006 31804 30012 31816
rect 28951 31776 30012 31804
rect 28951 31773 28963 31776
rect 28905 31767 28963 31773
rect 30006 31764 30012 31776
rect 30064 31764 30070 31816
rect 11149 31739 11207 31745
rect 11149 31705 11161 31739
rect 11195 31736 11207 31739
rect 11606 31736 11612 31748
rect 11195 31708 11612 31736
rect 11195 31705 11207 31708
rect 11149 31699 11207 31705
rect 11606 31696 11612 31708
rect 11664 31696 11670 31748
rect 12250 31736 12256 31748
rect 12211 31708 12256 31736
rect 12250 31696 12256 31708
rect 12308 31696 12314 31748
rect 15930 31736 15936 31748
rect 13478 31708 15936 31736
rect 15930 31696 15936 31708
rect 15988 31696 15994 31748
rect 16301 31739 16359 31745
rect 16301 31705 16313 31739
rect 16347 31736 16359 31739
rect 16574 31736 16580 31748
rect 16347 31708 16580 31736
rect 16347 31705 16359 31708
rect 16301 31699 16359 31705
rect 16574 31696 16580 31708
rect 16632 31696 16638 31748
rect 19613 31739 19671 31745
rect 19613 31705 19625 31739
rect 19659 31736 19671 31739
rect 20717 31739 20775 31745
rect 20717 31736 20729 31739
rect 19659 31708 20729 31736
rect 19659 31705 19671 31708
rect 19613 31699 19671 31705
rect 20717 31705 20729 31708
rect 20763 31705 20775 31739
rect 23017 31739 23075 31745
rect 23017 31736 23029 31739
rect 20717 31699 20775 31705
rect 22940 31708 23029 31736
rect 22940 31680 22968 31708
rect 23017 31705 23029 31708
rect 23063 31705 23075 31739
rect 23017 31699 23075 31705
rect 23109 31739 23167 31745
rect 23109 31705 23121 31739
rect 23155 31736 23167 31739
rect 23198 31736 23204 31748
rect 23155 31708 23204 31736
rect 23155 31705 23167 31708
rect 23109 31699 23167 31705
rect 23198 31696 23204 31708
rect 23256 31696 23262 31748
rect 26050 31696 26056 31748
rect 26108 31736 26114 31748
rect 26145 31739 26203 31745
rect 26145 31736 26157 31739
rect 26108 31708 26157 31736
rect 26108 31696 26114 31708
rect 26145 31705 26157 31708
rect 26191 31705 26203 31739
rect 26145 31699 26203 31705
rect 1762 31668 1768 31680
rect 1723 31640 1768 31668
rect 1762 31628 1768 31640
rect 1820 31628 1826 31680
rect 3602 31628 3608 31680
rect 3660 31668 3666 31680
rect 13630 31668 13636 31680
rect 3660 31640 13636 31668
rect 3660 31628 3666 31640
rect 13630 31628 13636 31640
rect 13688 31628 13694 31680
rect 13722 31628 13728 31680
rect 13780 31668 13786 31680
rect 13780 31640 13825 31668
rect 13780 31628 13786 31640
rect 14182 31628 14188 31680
rect 14240 31668 14246 31680
rect 14918 31668 14924 31680
rect 14240 31640 14924 31668
rect 14240 31628 14246 31640
rect 14918 31628 14924 31640
rect 14976 31628 14982 31680
rect 17954 31628 17960 31680
rect 18012 31668 18018 31680
rect 18785 31671 18843 31677
rect 18785 31668 18797 31671
rect 18012 31640 18797 31668
rect 18012 31628 18018 31640
rect 18785 31637 18797 31640
rect 18831 31637 18843 31671
rect 18785 31631 18843 31637
rect 19334 31628 19340 31680
rect 19392 31668 19398 31680
rect 20070 31668 20076 31680
rect 19392 31640 20076 31668
rect 19392 31628 19398 31640
rect 20070 31628 20076 31640
rect 20128 31628 20134 31680
rect 22922 31628 22928 31680
rect 22980 31628 22986 31680
rect 25314 31628 25320 31680
rect 25372 31668 25378 31680
rect 25409 31671 25467 31677
rect 25409 31668 25421 31671
rect 25372 31640 25421 31668
rect 25372 31628 25378 31640
rect 25409 31637 25421 31640
rect 25455 31637 25467 31671
rect 28166 31668 28172 31680
rect 28127 31640 28172 31668
rect 25409 31631 25467 31637
rect 28166 31628 28172 31640
rect 28224 31628 28230 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 5442 31464 5448 31476
rect 3160 31436 5448 31464
rect 3160 31396 3188 31436
rect 5442 31424 5448 31436
rect 5500 31424 5506 31476
rect 14844 31436 19932 31464
rect 14844 31408 14872 31436
rect 3068 31368 3188 31396
rect 3329 31399 3387 31405
rect 3068 31337 3096 31368
rect 3329 31365 3341 31399
rect 3375 31396 3387 31399
rect 3602 31396 3608 31408
rect 3375 31368 3608 31396
rect 3375 31365 3387 31368
rect 3329 31359 3387 31365
rect 3602 31356 3608 31368
rect 3660 31356 3666 31408
rect 5350 31396 5356 31408
rect 4554 31368 5356 31396
rect 5350 31356 5356 31368
rect 5408 31356 5414 31408
rect 12066 31396 12072 31408
rect 9154 31368 12072 31396
rect 12066 31356 12072 31368
rect 12124 31356 12130 31408
rect 13725 31399 13783 31405
rect 13725 31365 13737 31399
rect 13771 31396 13783 31399
rect 14826 31396 14832 31408
rect 13771 31368 14832 31396
rect 13771 31365 13783 31368
rect 13725 31359 13783 31365
rect 14826 31356 14832 31368
rect 14884 31356 14890 31408
rect 14918 31356 14924 31408
rect 14976 31396 14982 31408
rect 17770 31396 17776 31408
rect 14976 31368 17776 31396
rect 14976 31356 14982 31368
rect 17770 31356 17776 31368
rect 17828 31356 17834 31408
rect 17865 31399 17923 31405
rect 17865 31365 17877 31399
rect 17911 31396 17923 31399
rect 19610 31396 19616 31408
rect 17911 31368 19616 31396
rect 17911 31365 17923 31368
rect 17865 31359 17923 31365
rect 19610 31356 19616 31368
rect 19668 31356 19674 31408
rect 19904 31396 19932 31436
rect 19978 31424 19984 31476
rect 20036 31464 20042 31476
rect 20533 31467 20591 31473
rect 20533 31464 20545 31467
rect 20036 31436 20545 31464
rect 20036 31424 20042 31436
rect 20533 31433 20545 31436
rect 20579 31433 20591 31467
rect 20533 31427 20591 31433
rect 20714 31424 20720 31476
rect 20772 31464 20778 31476
rect 21361 31467 21419 31473
rect 21361 31464 21373 31467
rect 20772 31436 21373 31464
rect 20772 31424 20778 31436
rect 21361 31433 21373 31436
rect 21407 31433 21419 31467
rect 21361 31427 21419 31433
rect 23474 31424 23480 31476
rect 23532 31464 23538 31476
rect 23750 31464 23756 31476
rect 23532 31436 23756 31464
rect 23532 31424 23538 31436
rect 23750 31424 23756 31436
rect 23808 31424 23814 31476
rect 23842 31424 23848 31476
rect 23900 31464 23906 31476
rect 23937 31467 23995 31473
rect 23937 31464 23949 31467
rect 23900 31436 23949 31464
rect 23900 31424 23906 31436
rect 23937 31433 23949 31436
rect 23983 31433 23995 31467
rect 28074 31464 28080 31476
rect 28035 31436 28080 31464
rect 23937 31427 23995 31433
rect 28074 31424 28080 31436
rect 28132 31424 28138 31476
rect 29825 31467 29883 31473
rect 29825 31433 29837 31467
rect 29871 31433 29883 31467
rect 29825 31427 29883 31433
rect 24118 31396 24124 31408
rect 19904 31368 24124 31396
rect 3053 31331 3111 31337
rect 3053 31297 3065 31331
rect 3099 31297 3111 31331
rect 11698 31328 11704 31340
rect 11659 31300 11704 31328
rect 3053 31291 3111 31297
rect 11698 31288 11704 31300
rect 11756 31288 11762 31340
rect 13110 31300 14688 31328
rect 7653 31263 7711 31269
rect 7653 31229 7665 31263
rect 7699 31260 7711 31263
rect 7929 31263 7987 31269
rect 7699 31232 7788 31260
rect 7699 31229 7711 31232
rect 7653 31223 7711 31229
rect 4706 31084 4712 31136
rect 4764 31124 4770 31136
rect 4801 31127 4859 31133
rect 4801 31124 4813 31127
rect 4764 31096 4813 31124
rect 4764 31084 4770 31096
rect 4801 31093 4813 31096
rect 4847 31093 4859 31127
rect 7760 31124 7788 31232
rect 7929 31229 7941 31263
rect 7975 31260 7987 31263
rect 9306 31260 9312 31272
rect 7975 31232 9312 31260
rect 7975 31229 7987 31232
rect 7929 31223 7987 31229
rect 9306 31220 9312 31232
rect 9364 31220 9370 31272
rect 11146 31220 11152 31272
rect 11204 31260 11210 31272
rect 11606 31260 11612 31272
rect 11204 31232 11612 31260
rect 11204 31220 11210 31232
rect 11606 31220 11612 31232
rect 11664 31260 11670 31272
rect 11977 31263 12035 31269
rect 11977 31260 11989 31263
rect 11664 31232 11989 31260
rect 11664 31220 11670 31232
rect 11977 31229 11989 31232
rect 12023 31229 12035 31263
rect 11977 31223 12035 31229
rect 12066 31220 12072 31272
rect 12124 31260 12130 31272
rect 12124 31232 14596 31260
rect 12124 31220 12130 31232
rect 9122 31124 9128 31136
rect 7760 31096 9128 31124
rect 4801 31087 4859 31093
rect 9122 31084 9128 31096
rect 9180 31084 9186 31136
rect 9401 31127 9459 31133
rect 9401 31093 9413 31127
rect 9447 31124 9459 31127
rect 9766 31124 9772 31136
rect 9447 31096 9772 31124
rect 9447 31093 9459 31096
rect 9401 31087 9459 31093
rect 9766 31084 9772 31096
rect 9824 31084 9830 31136
rect 14568 31124 14596 31232
rect 14660 31192 14688 31300
rect 14734 31288 14740 31340
rect 14792 31328 14798 31340
rect 17494 31328 17500 31340
rect 14792 31300 17500 31328
rect 14792 31288 14798 31300
rect 17494 31288 17500 31300
rect 17552 31288 17558 31340
rect 19797 31331 19855 31337
rect 19797 31297 19809 31331
rect 19843 31328 19855 31331
rect 19978 31328 19984 31340
rect 19843 31300 19984 31328
rect 19843 31297 19855 31300
rect 19797 31291 19855 31297
rect 19978 31288 19984 31300
rect 20036 31328 20042 31340
rect 20162 31328 20168 31340
rect 20036 31300 20168 31328
rect 20036 31288 20042 31300
rect 20162 31288 20168 31300
rect 20220 31288 20226 31340
rect 20456 31337 20484 31368
rect 24118 31356 24124 31368
rect 24176 31356 24182 31408
rect 25314 31396 25320 31408
rect 25275 31368 25320 31396
rect 25314 31356 25320 31368
rect 25372 31356 25378 31408
rect 29840 31396 29868 31427
rect 29840 31368 30696 31396
rect 20441 31331 20499 31337
rect 20441 31297 20453 31331
rect 20487 31297 20499 31331
rect 21269 31331 21327 31337
rect 21269 31328 21281 31331
rect 20441 31291 20499 31297
rect 21100 31300 21281 31328
rect 17037 31263 17095 31269
rect 17037 31229 17049 31263
rect 17083 31260 17095 31263
rect 17773 31263 17831 31269
rect 17773 31260 17785 31263
rect 17083 31232 17785 31260
rect 17083 31229 17095 31232
rect 17037 31223 17095 31229
rect 17773 31229 17785 31232
rect 17819 31229 17831 31263
rect 17773 31223 17831 31229
rect 17862 31220 17868 31272
rect 17920 31260 17926 31272
rect 18782 31260 18788 31272
rect 17920 31232 18788 31260
rect 17920 31220 17926 31232
rect 18782 31220 18788 31232
rect 18840 31220 18846 31272
rect 19058 31220 19064 31272
rect 19116 31260 19122 31272
rect 20714 31260 20720 31272
rect 19116 31232 20720 31260
rect 19116 31220 19122 31232
rect 20714 31220 20720 31232
rect 20772 31220 20778 31272
rect 20990 31192 20996 31204
rect 14660 31164 20996 31192
rect 20990 31152 20996 31164
rect 21048 31152 21054 31204
rect 16390 31124 16396 31136
rect 14568 31096 16396 31124
rect 16390 31084 16396 31096
rect 16448 31084 16454 31136
rect 16482 31084 16488 31136
rect 16540 31124 16546 31136
rect 19889 31127 19947 31133
rect 19889 31124 19901 31127
rect 16540 31096 19901 31124
rect 16540 31084 16546 31096
rect 19889 31093 19901 31096
rect 19935 31093 19947 31127
rect 19889 31087 19947 31093
rect 20530 31084 20536 31136
rect 20588 31124 20594 31136
rect 21100 31124 21128 31300
rect 21269 31297 21281 31300
rect 21315 31297 21327 31331
rect 21269 31291 21327 31297
rect 21450 31288 21456 31340
rect 21508 31328 21514 31340
rect 22002 31328 22008 31340
rect 21508 31300 22008 31328
rect 21508 31288 21514 31300
rect 22002 31288 22008 31300
rect 22060 31288 22066 31340
rect 23385 31331 23443 31337
rect 23385 31297 23397 31331
rect 23431 31328 23443 31331
rect 23750 31328 23756 31340
rect 23431 31300 23756 31328
rect 23431 31297 23443 31300
rect 23385 31291 23443 31297
rect 23750 31288 23756 31300
rect 23808 31288 23814 31340
rect 23842 31288 23848 31340
rect 23900 31328 23906 31340
rect 27433 31331 27491 31337
rect 23900 31300 23945 31328
rect 23900 31288 23906 31300
rect 27433 31297 27445 31331
rect 27479 31328 27491 31331
rect 28166 31328 28172 31340
rect 27479 31300 28172 31328
rect 27479 31297 27491 31300
rect 27433 31291 27491 31297
rect 28166 31288 28172 31300
rect 28224 31288 28230 31340
rect 29822 31288 29828 31340
rect 29880 31328 29886 31340
rect 30006 31328 30012 31340
rect 29880 31300 30012 31328
rect 29880 31288 29886 31300
rect 30006 31288 30012 31300
rect 30064 31288 30070 31340
rect 30668 31337 30696 31368
rect 30653 31331 30711 31337
rect 30653 31297 30665 31331
rect 30699 31297 30711 31331
rect 30653 31291 30711 31297
rect 22189 31263 22247 31269
rect 22189 31229 22201 31263
rect 22235 31260 22247 31263
rect 25222 31260 25228 31272
rect 22235 31232 23244 31260
rect 25183 31232 25228 31260
rect 22235 31229 22247 31232
rect 22189 31223 22247 31229
rect 23216 31201 23244 31232
rect 25222 31220 25228 31232
rect 25280 31220 25286 31272
rect 26145 31263 26203 31269
rect 26145 31229 26157 31263
rect 26191 31260 26203 31263
rect 27246 31260 27252 31272
rect 26191 31232 27252 31260
rect 26191 31229 26203 31232
rect 26145 31223 26203 31229
rect 27246 31220 27252 31232
rect 27304 31220 27310 31272
rect 27617 31263 27675 31269
rect 27617 31229 27629 31263
rect 27663 31260 27675 31263
rect 27663 31232 30512 31260
rect 27663 31229 27675 31232
rect 27617 31223 27675 31229
rect 30484 31201 30512 31232
rect 23201 31195 23259 31201
rect 23201 31161 23213 31195
rect 23247 31161 23259 31195
rect 23201 31155 23259 31161
rect 30469 31195 30527 31201
rect 30469 31161 30481 31195
rect 30515 31161 30527 31195
rect 30469 31155 30527 31161
rect 22554 31124 22560 31136
rect 20588 31096 21128 31124
rect 22515 31096 22560 31124
rect 20588 31084 20594 31096
rect 22554 31084 22560 31096
rect 22612 31084 22618 31136
rect 24762 31084 24768 31136
rect 24820 31124 24826 31136
rect 38010 31124 38016 31136
rect 24820 31096 38016 31124
rect 24820 31084 24826 31096
rect 38010 31084 38016 31096
rect 38068 31084 38074 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 12986 30920 12992 30932
rect 5460 30892 12992 30920
rect 5460 30796 5488 30892
rect 12986 30880 12992 30892
rect 13044 30880 13050 30932
rect 13814 30880 13820 30932
rect 13872 30920 13878 30932
rect 19889 30923 19947 30929
rect 19889 30920 19901 30923
rect 13872 30892 19901 30920
rect 13872 30880 13878 30892
rect 19889 30889 19901 30892
rect 19935 30889 19947 30923
rect 19889 30883 19947 30889
rect 20162 30880 20168 30932
rect 20220 30920 20226 30932
rect 23750 30920 23756 30932
rect 20220 30892 22094 30920
rect 23711 30892 23756 30920
rect 20220 30880 20226 30892
rect 12161 30855 12219 30861
rect 12161 30821 12173 30855
rect 12207 30852 12219 30855
rect 15562 30852 15568 30864
rect 12207 30824 15568 30852
rect 12207 30821 12219 30824
rect 12161 30815 12219 30821
rect 15562 30812 15568 30824
rect 15620 30812 15626 30864
rect 17126 30812 17132 30864
rect 17184 30852 17190 30864
rect 17184 30824 17540 30852
rect 17184 30812 17190 30824
rect 4249 30787 4307 30793
rect 4249 30753 4261 30787
rect 4295 30784 4307 30787
rect 5442 30784 5448 30796
rect 4295 30756 5448 30784
rect 4295 30753 4307 30756
rect 4249 30747 4307 30753
rect 5442 30744 5448 30756
rect 5500 30744 5506 30796
rect 6086 30744 6092 30796
rect 6144 30784 6150 30796
rect 6365 30787 6423 30793
rect 6365 30784 6377 30787
rect 6144 30756 6377 30784
rect 6144 30744 6150 30756
rect 6365 30753 6377 30756
rect 6411 30753 6423 30787
rect 6365 30747 6423 30753
rect 6641 30787 6699 30793
rect 6641 30753 6653 30787
rect 6687 30784 6699 30787
rect 9582 30784 9588 30796
rect 6687 30756 9588 30784
rect 6687 30753 6699 30756
rect 6641 30747 6699 30753
rect 9582 30744 9588 30756
rect 9640 30744 9646 30796
rect 10413 30787 10471 30793
rect 10413 30753 10425 30787
rect 10459 30784 10471 30787
rect 10778 30784 10784 30796
rect 10459 30756 10784 30784
rect 10459 30753 10471 30756
rect 10413 30747 10471 30753
rect 10778 30744 10784 30756
rect 10836 30744 10842 30796
rect 15838 30784 15844 30796
rect 15799 30756 15844 30784
rect 15838 30744 15844 30756
rect 15896 30744 15902 30796
rect 16117 30787 16175 30793
rect 16117 30753 16129 30787
rect 16163 30784 16175 30787
rect 16574 30784 16580 30796
rect 16163 30756 16580 30784
rect 16163 30753 16175 30756
rect 16117 30747 16175 30753
rect 16574 30744 16580 30756
rect 16632 30744 16638 30796
rect 16666 30744 16672 30796
rect 16724 30784 16730 30796
rect 17512 30784 17540 30824
rect 17678 30812 17684 30864
rect 17736 30852 17742 30864
rect 22066 30852 22094 30892
rect 23750 30880 23756 30892
rect 23808 30880 23814 30932
rect 17736 30824 21680 30852
rect 22066 30824 23980 30852
rect 17736 30812 17742 30824
rect 21652 30796 21680 30824
rect 20346 30784 20352 30796
rect 16724 30756 17448 30784
rect 17512 30756 20352 30784
rect 16724 30744 16730 30756
rect 2774 30676 2780 30728
rect 2832 30716 2838 30728
rect 3973 30719 4031 30725
rect 3973 30716 3985 30719
rect 2832 30688 3985 30716
rect 2832 30676 2838 30688
rect 3973 30685 3985 30688
rect 4019 30685 4031 30719
rect 3973 30679 4031 30685
rect 5350 30676 5356 30728
rect 5408 30676 5414 30728
rect 17420 30710 17448 30756
rect 20346 30744 20352 30756
rect 20404 30744 20410 30796
rect 21634 30784 21640 30796
rect 21547 30756 21640 30784
rect 21634 30744 21640 30756
rect 21692 30744 21698 30796
rect 22094 30744 22100 30796
rect 22152 30784 22158 30796
rect 23014 30784 23020 30796
rect 22152 30756 23020 30784
rect 22152 30744 22158 30756
rect 23014 30744 23020 30756
rect 23072 30744 23078 30796
rect 18322 30716 18328 30728
rect 17512 30710 18328 30716
rect 17420 30688 18328 30710
rect 17420 30682 17540 30688
rect 18322 30676 18328 30688
rect 18380 30676 18386 30728
rect 18693 30719 18751 30725
rect 18693 30685 18705 30719
rect 18739 30716 18751 30719
rect 19334 30716 19340 30728
rect 18739 30688 19340 30716
rect 18739 30685 18751 30688
rect 18693 30679 18751 30685
rect 19334 30676 19340 30688
rect 19392 30676 19398 30728
rect 19797 30719 19855 30725
rect 19797 30685 19809 30719
rect 19843 30716 19855 30719
rect 19843 30688 20300 30716
rect 19843 30685 19855 30688
rect 19797 30679 19855 30685
rect 10689 30651 10747 30657
rect 7866 30620 10640 30648
rect 4614 30540 4620 30592
rect 4672 30580 4678 30592
rect 5721 30583 5779 30589
rect 5721 30580 5733 30583
rect 4672 30552 5733 30580
rect 4672 30540 4678 30552
rect 5721 30549 5733 30552
rect 5767 30549 5779 30583
rect 5721 30543 5779 30549
rect 8113 30583 8171 30589
rect 8113 30549 8125 30583
rect 8159 30580 8171 30583
rect 8478 30580 8484 30592
rect 8159 30552 8484 30580
rect 8159 30549 8171 30552
rect 8113 30543 8171 30549
rect 8478 30540 8484 30552
rect 8536 30540 8542 30592
rect 10612 30580 10640 30620
rect 10689 30617 10701 30651
rect 10735 30648 10747 30651
rect 10778 30648 10784 30660
rect 10735 30620 10784 30648
rect 10735 30617 10747 30620
rect 10689 30611 10747 30617
rect 10778 30608 10784 30620
rect 10836 30608 10842 30660
rect 17954 30648 17960 30660
rect 11914 30620 16436 30648
rect 17342 30620 17960 30648
rect 15102 30580 15108 30592
rect 10612 30552 15108 30580
rect 15102 30540 15108 30552
rect 15160 30540 15166 30592
rect 16408 30580 16436 30620
rect 17954 30608 17960 30620
rect 18012 30608 18018 30660
rect 18046 30608 18052 30660
rect 18104 30648 18110 30660
rect 20162 30648 20168 30660
rect 18104 30620 20168 30648
rect 18104 30608 18110 30620
rect 20162 30608 20168 30620
rect 20220 30608 20226 30660
rect 20272 30648 20300 30688
rect 20714 30676 20720 30728
rect 20772 30716 20778 30728
rect 20901 30719 20959 30725
rect 20901 30716 20913 30719
rect 20772 30688 20913 30716
rect 20772 30676 20778 30688
rect 20901 30685 20913 30688
rect 20947 30716 20959 30719
rect 21082 30716 21088 30728
rect 20947 30688 21088 30716
rect 20947 30685 20959 30688
rect 20901 30679 20959 30685
rect 21082 30676 21088 30688
rect 21140 30676 21146 30728
rect 23106 30716 23112 30728
rect 23067 30688 23112 30716
rect 23106 30676 23112 30688
rect 23164 30676 23170 30728
rect 23952 30725 23980 30824
rect 28074 30812 28080 30864
rect 28132 30812 28138 30864
rect 26237 30787 26295 30793
rect 26237 30753 26249 30787
rect 26283 30784 26295 30787
rect 27154 30784 27160 30796
rect 26283 30756 27160 30784
rect 26283 30753 26295 30756
rect 26237 30747 26295 30753
rect 27154 30744 27160 30756
rect 27212 30744 27218 30796
rect 27893 30787 27951 30793
rect 27893 30753 27905 30787
rect 27939 30784 27951 30787
rect 28092 30784 28120 30812
rect 27939 30756 28120 30784
rect 27939 30753 27951 30756
rect 27893 30747 27951 30753
rect 23937 30719 23995 30725
rect 23937 30685 23949 30719
rect 23983 30685 23995 30719
rect 23937 30679 23995 30685
rect 28077 30719 28135 30725
rect 28077 30685 28089 30719
rect 28123 30716 28135 30719
rect 29270 30716 29276 30728
rect 28123 30688 29276 30716
rect 28123 30685 28135 30688
rect 28077 30679 28135 30685
rect 29270 30676 29276 30688
rect 29328 30676 29334 30728
rect 38286 30716 38292 30728
rect 38247 30688 38292 30716
rect 38286 30676 38292 30688
rect 38344 30676 38350 30728
rect 21174 30648 21180 30660
rect 20272 30620 21180 30648
rect 21174 30608 21180 30620
rect 21232 30608 21238 30660
rect 21726 30608 21732 30660
rect 21784 30648 21790 30660
rect 26329 30651 26387 30657
rect 21784 30620 21829 30648
rect 21784 30608 21790 30620
rect 26329 30617 26341 30651
rect 26375 30617 26387 30651
rect 26329 30611 26387 30617
rect 17126 30580 17132 30592
rect 16408 30552 17132 30580
rect 17126 30540 17132 30552
rect 17184 30540 17190 30592
rect 17589 30583 17647 30589
rect 17589 30549 17601 30583
rect 17635 30580 17647 30583
rect 17770 30580 17776 30592
rect 17635 30552 17776 30580
rect 17635 30549 17647 30552
rect 17589 30543 17647 30549
rect 17770 30540 17776 30552
rect 17828 30540 17834 30592
rect 18782 30580 18788 30592
rect 18743 30552 18788 30580
rect 18782 30540 18788 30552
rect 18840 30540 18846 30592
rect 19150 30540 19156 30592
rect 19208 30580 19214 30592
rect 20530 30580 20536 30592
rect 19208 30552 20536 30580
rect 19208 30540 19214 30552
rect 20530 30540 20536 30552
rect 20588 30540 20594 30592
rect 20990 30580 20996 30592
rect 20951 30552 20996 30580
rect 20990 30540 20996 30552
rect 21048 30540 21054 30592
rect 23201 30583 23259 30589
rect 23201 30549 23213 30583
rect 23247 30580 23259 30583
rect 26344 30580 26372 30611
rect 26602 30608 26608 30660
rect 26660 30648 26666 30660
rect 27249 30651 27307 30657
rect 27249 30648 27261 30651
rect 26660 30620 27261 30648
rect 26660 30608 26666 30620
rect 27249 30617 27261 30620
rect 27295 30617 27307 30651
rect 27249 30611 27307 30617
rect 28534 30580 28540 30592
rect 23247 30552 26372 30580
rect 28495 30552 28540 30580
rect 23247 30549 23259 30552
rect 23201 30543 23259 30549
rect 28534 30540 28540 30552
rect 28592 30540 28598 30592
rect 38102 30580 38108 30592
rect 38063 30552 38108 30580
rect 38102 30540 38108 30552
rect 38160 30540 38166 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 8220 30348 9168 30376
rect 6178 30268 6184 30320
rect 6236 30308 6242 30320
rect 6546 30308 6552 30320
rect 6236 30280 6552 30308
rect 6236 30268 6242 30280
rect 6546 30268 6552 30280
rect 6604 30308 6610 30320
rect 8220 30308 8248 30348
rect 6604 30280 8248 30308
rect 9140 30308 9168 30348
rect 15764 30348 16252 30376
rect 9861 30311 9919 30317
rect 9861 30308 9873 30311
rect 9140 30280 9873 30308
rect 6604 30268 6610 30280
rect 9861 30277 9873 30280
rect 9907 30308 9919 30311
rect 11330 30308 11336 30320
rect 9907 30280 11336 30308
rect 9907 30277 9919 30280
rect 9861 30271 9919 30277
rect 11330 30268 11336 30280
rect 11388 30308 11394 30320
rect 11974 30308 11980 30320
rect 11388 30280 11980 30308
rect 11388 30268 11394 30280
rect 11974 30268 11980 30280
rect 12032 30268 12038 30320
rect 15764 30308 15792 30348
rect 14306 30280 15792 30308
rect 15838 30268 15844 30320
rect 15896 30308 15902 30320
rect 16117 30311 16175 30317
rect 16117 30308 16129 30311
rect 15896 30280 16129 30308
rect 15896 30268 15902 30280
rect 16117 30277 16129 30280
rect 16163 30277 16175 30311
rect 16224 30308 16252 30348
rect 16758 30336 16764 30388
rect 16816 30376 16822 30388
rect 17218 30376 17224 30388
rect 16816 30348 17224 30376
rect 16816 30336 16822 30348
rect 17218 30336 17224 30348
rect 17276 30336 17282 30388
rect 18966 30376 18972 30388
rect 17512 30348 18972 30376
rect 17512 30308 17540 30348
rect 18966 30336 18972 30348
rect 19024 30336 19030 30388
rect 19334 30336 19340 30388
rect 19392 30376 19398 30388
rect 20070 30376 20076 30388
rect 19392 30348 20076 30376
rect 19392 30336 19398 30348
rect 20070 30336 20076 30348
rect 20128 30336 20134 30388
rect 21358 30376 21364 30388
rect 20640 30348 21364 30376
rect 19242 30308 19248 30320
rect 16224 30280 17540 30308
rect 18354 30280 19248 30308
rect 16117 30271 16175 30277
rect 1578 30240 1584 30252
rect 1539 30212 1584 30240
rect 1578 30200 1584 30212
rect 1636 30200 1642 30252
rect 6086 30200 6092 30252
rect 6144 30240 6150 30252
rect 7561 30243 7619 30249
rect 7561 30240 7573 30243
rect 6144 30212 7573 30240
rect 6144 30200 6150 30212
rect 7561 30209 7573 30212
rect 7607 30209 7619 30243
rect 12342 30240 12348 30252
rect 8970 30212 12348 30240
rect 7561 30203 7619 30209
rect 7576 30172 7604 30203
rect 12342 30200 12348 30212
rect 12400 30200 12406 30252
rect 15286 30240 15292 30252
rect 14476 30212 15292 30240
rect 9674 30172 9680 30184
rect 7576 30144 9680 30172
rect 9674 30132 9680 30144
rect 9732 30172 9738 30184
rect 10597 30175 10655 30181
rect 10597 30172 10609 30175
rect 9732 30144 10609 30172
rect 9732 30132 9738 30144
rect 10597 30141 10609 30144
rect 10643 30141 10655 30175
rect 10597 30135 10655 30141
rect 11698 30132 11704 30184
rect 11756 30172 11762 30184
rect 12066 30172 12072 30184
rect 11756 30144 12072 30172
rect 11756 30132 11762 30144
rect 12066 30132 12072 30144
rect 12124 30172 12130 30184
rect 12805 30175 12863 30181
rect 12805 30172 12817 30175
rect 12124 30144 12817 30172
rect 12124 30132 12130 30144
rect 12805 30141 12817 30144
rect 12851 30141 12863 30175
rect 12805 30135 12863 30141
rect 13081 30175 13139 30181
rect 13081 30141 13093 30175
rect 13127 30172 13139 30175
rect 14476 30172 14504 30212
rect 15286 30200 15292 30212
rect 15344 30200 15350 30252
rect 15381 30243 15439 30249
rect 15381 30209 15393 30243
rect 15427 30240 15439 30243
rect 16132 30240 16160 30271
rect 19242 30268 19248 30280
rect 19300 30268 19306 30320
rect 16853 30243 16911 30249
rect 16853 30240 16865 30243
rect 15427 30212 15516 30240
rect 16132 30212 16865 30240
rect 15427 30209 15439 30212
rect 15381 30203 15439 30209
rect 13127 30144 14504 30172
rect 13127 30141 13139 30144
rect 13081 30135 13139 30141
rect 15488 30104 15516 30212
rect 16853 30209 16865 30212
rect 16899 30209 16911 30243
rect 19426 30240 19432 30252
rect 19387 30212 19432 30240
rect 16853 30203 16911 30209
rect 19426 30200 19432 30212
rect 19484 30200 19490 30252
rect 19518 30200 19524 30252
rect 19576 30240 19582 30252
rect 19978 30240 19984 30252
rect 19576 30212 19984 30240
rect 19576 30200 19582 30212
rect 19978 30200 19984 30212
rect 20036 30240 20042 30252
rect 20073 30243 20131 30249
rect 20073 30240 20085 30243
rect 20036 30212 20085 30240
rect 20036 30200 20042 30212
rect 20073 30209 20085 30212
rect 20119 30240 20131 30243
rect 20640 30240 20668 30348
rect 21358 30336 21364 30348
rect 21416 30336 21422 30388
rect 29270 30376 29276 30388
rect 24780 30348 25084 30376
rect 29231 30348 29276 30376
rect 20806 30268 20812 30320
rect 20864 30308 20870 30320
rect 20864 30280 23428 30308
rect 20864 30268 20870 30280
rect 20119 30212 20668 30240
rect 20717 30243 20775 30249
rect 20119 30209 20131 30212
rect 20073 30203 20131 30209
rect 20717 30209 20729 30243
rect 20763 30240 20775 30243
rect 21266 30240 21272 30252
rect 20763 30212 21272 30240
rect 20763 30209 20775 30212
rect 20717 30203 20775 30209
rect 21266 30200 21272 30212
rect 21324 30200 21330 30252
rect 22186 30240 22192 30252
rect 22147 30212 22192 30240
rect 22186 30200 22192 30212
rect 22244 30200 22250 30252
rect 22278 30200 22284 30252
rect 22336 30240 22342 30252
rect 23400 30249 23428 30280
rect 23566 30268 23572 30320
rect 23624 30308 23630 30320
rect 24213 30311 24271 30317
rect 24213 30308 24225 30311
rect 23624 30280 24225 30308
rect 23624 30268 23630 30280
rect 24213 30277 24225 30280
rect 24259 30277 24271 30311
rect 24213 30271 24271 30277
rect 24394 30268 24400 30320
rect 24452 30308 24458 30320
rect 24780 30308 24808 30348
rect 24946 30308 24952 30320
rect 24452 30280 24808 30308
rect 24907 30280 24952 30308
rect 24452 30268 24458 30280
rect 24946 30268 24952 30280
rect 25004 30268 25010 30320
rect 25056 30308 25084 30348
rect 29270 30336 29276 30348
rect 29328 30336 29334 30388
rect 27249 30311 27307 30317
rect 25056 30280 27200 30308
rect 27172 30249 27200 30280
rect 27249 30277 27261 30311
rect 27295 30308 27307 30311
rect 27338 30308 27344 30320
rect 27295 30280 27344 30308
rect 27295 30277 27307 30280
rect 27249 30271 27307 30277
rect 27338 30268 27344 30280
rect 27396 30268 27402 30320
rect 36814 30308 36820 30320
rect 31726 30280 36820 30308
rect 23385 30243 23443 30249
rect 22336 30212 22381 30240
rect 22336 30200 22342 30212
rect 23385 30209 23397 30243
rect 23431 30209 23443 30243
rect 23385 30203 23443 30209
rect 24121 30243 24179 30249
rect 24121 30209 24133 30243
rect 24167 30209 24179 30243
rect 24121 30203 24179 30209
rect 26329 30243 26387 30249
rect 26329 30209 26341 30243
rect 26375 30209 26387 30243
rect 26329 30203 26387 30209
rect 27157 30243 27215 30249
rect 27157 30209 27169 30243
rect 27203 30209 27215 30243
rect 27157 30203 27215 30209
rect 16206 30132 16212 30184
rect 16264 30172 16270 30184
rect 17129 30175 17187 30181
rect 17129 30172 17141 30175
rect 16264 30144 17141 30172
rect 16264 30132 16270 30144
rect 17129 30141 17141 30144
rect 17175 30172 17187 30175
rect 17218 30172 17224 30184
rect 17175 30144 17224 30172
rect 17175 30141 17187 30144
rect 17129 30135 17187 30141
rect 17218 30132 17224 30144
rect 17276 30132 17282 30184
rect 17494 30132 17500 30184
rect 17552 30172 17558 30184
rect 20165 30175 20223 30181
rect 20165 30172 20177 30175
rect 17552 30144 20177 30172
rect 17552 30132 17558 30144
rect 20165 30141 20177 30144
rect 20211 30141 20223 30175
rect 22922 30172 22928 30184
rect 20165 30135 20223 30141
rect 20272 30144 22928 30172
rect 14108 30076 15516 30104
rect 1762 30036 1768 30048
rect 1723 30008 1768 30036
rect 1762 29996 1768 30008
rect 1820 29996 1826 30048
rect 7834 30045 7840 30048
rect 7824 30039 7840 30045
rect 7824 30005 7836 30039
rect 7824 29999 7840 30005
rect 7834 29996 7840 29999
rect 7892 29996 7898 30048
rect 9306 30036 9312 30048
rect 9267 30008 9312 30036
rect 9306 29996 9312 30008
rect 9364 29996 9370 30048
rect 11974 29996 11980 30048
rect 12032 30036 12038 30048
rect 14108 30036 14136 30076
rect 18138 30064 18144 30116
rect 18196 30104 18202 30116
rect 20272 30104 20300 30144
rect 22922 30132 22928 30144
rect 22980 30132 22986 30184
rect 23198 30132 23204 30184
rect 23256 30172 23262 30184
rect 23477 30175 23535 30181
rect 23477 30172 23489 30175
rect 23256 30144 23489 30172
rect 23256 30132 23262 30144
rect 23477 30141 23489 30144
rect 23523 30141 23535 30175
rect 24136 30172 24164 30203
rect 24210 30172 24216 30184
rect 24136 30144 24216 30172
rect 23477 30135 23535 30141
rect 24210 30132 24216 30144
rect 24268 30132 24274 30184
rect 24857 30175 24915 30181
rect 24857 30141 24869 30175
rect 24903 30141 24915 30175
rect 25774 30172 25780 30184
rect 25735 30144 25780 30172
rect 24857 30135 24915 30141
rect 18196 30076 20300 30104
rect 18196 30064 18202 30076
rect 21634 30064 21640 30116
rect 21692 30104 21698 30116
rect 24872 30104 24900 30135
rect 25774 30132 25780 30144
rect 25832 30132 25838 30184
rect 26344 30172 26372 30203
rect 27522 30200 27528 30252
rect 27580 30240 27586 30252
rect 28629 30243 28687 30249
rect 28629 30240 28641 30243
rect 27580 30212 28641 30240
rect 27580 30200 27586 30212
rect 28629 30209 28641 30212
rect 28675 30209 28687 30243
rect 28629 30203 28687 30209
rect 29457 30243 29515 30249
rect 29457 30209 29469 30243
rect 29503 30240 29515 30243
rect 29730 30240 29736 30252
rect 29503 30212 29736 30240
rect 29503 30209 29515 30212
rect 29457 30203 29515 30209
rect 29730 30200 29736 30212
rect 29788 30200 29794 30252
rect 31726 30172 31754 30280
rect 36814 30268 36820 30280
rect 36872 30268 36878 30320
rect 26344 30144 31754 30172
rect 21692 30076 24900 30104
rect 25792 30104 25820 30132
rect 27982 30104 27988 30116
rect 25792 30076 27988 30104
rect 21692 30064 21698 30076
rect 27982 30064 27988 30076
rect 28040 30064 28046 30116
rect 14550 30036 14556 30048
rect 12032 30008 14136 30036
rect 14511 30008 14556 30036
rect 12032 29996 12038 30008
rect 14550 29996 14556 30008
rect 14608 29996 14614 30048
rect 15194 29996 15200 30048
rect 15252 30036 15258 30048
rect 16390 30036 16396 30048
rect 15252 30008 16396 30036
rect 15252 29996 15258 30008
rect 16390 29996 16396 30008
rect 16448 29996 16454 30048
rect 16574 29996 16580 30048
rect 16632 30036 16638 30048
rect 18598 30036 18604 30048
rect 16632 30008 18604 30036
rect 16632 29996 16638 30008
rect 18598 29996 18604 30008
rect 18656 29996 18662 30048
rect 18690 29996 18696 30048
rect 18748 30036 18754 30048
rect 19521 30039 19579 30045
rect 19521 30036 19533 30039
rect 18748 30008 19533 30036
rect 18748 29996 18754 30008
rect 19521 30005 19533 30008
rect 19567 30005 19579 30039
rect 20806 30036 20812 30048
rect 20767 30008 20812 30036
rect 19521 29999 19579 30005
rect 20806 29996 20812 30008
rect 20864 29996 20870 30048
rect 20898 29996 20904 30048
rect 20956 30036 20962 30048
rect 23934 30036 23940 30048
rect 20956 30008 23940 30036
rect 20956 29996 20962 30008
rect 23934 29996 23940 30008
rect 23992 29996 23998 30048
rect 24302 29996 24308 30048
rect 24360 30036 24366 30048
rect 26421 30039 26479 30045
rect 26421 30036 26433 30039
rect 24360 30008 26433 30036
rect 24360 29996 24366 30008
rect 26421 30005 26433 30008
rect 26467 30005 26479 30039
rect 26421 29999 26479 30005
rect 28166 29996 28172 30048
rect 28224 30036 28230 30048
rect 28721 30039 28779 30045
rect 28721 30036 28733 30039
rect 28224 30008 28733 30036
rect 28224 29996 28230 30008
rect 28721 30005 28733 30008
rect 28767 30005 28779 30039
rect 28721 29999 28779 30005
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 4709 29835 4767 29841
rect 4709 29801 4721 29835
rect 4755 29832 4767 29835
rect 20898 29832 20904 29844
rect 4755 29804 20904 29832
rect 4755 29801 4767 29804
rect 4709 29795 4767 29801
rect 20898 29792 20904 29804
rect 20956 29792 20962 29844
rect 21726 29792 21732 29844
rect 21784 29832 21790 29844
rect 22373 29835 22431 29841
rect 22373 29832 22385 29835
rect 21784 29804 22385 29832
rect 21784 29792 21790 29804
rect 22373 29801 22385 29804
rect 22419 29801 22431 29835
rect 22373 29795 22431 29801
rect 23934 29792 23940 29844
rect 23992 29832 23998 29844
rect 24854 29832 24860 29844
rect 23992 29804 24860 29832
rect 23992 29792 23998 29804
rect 24854 29792 24860 29804
rect 24912 29792 24918 29844
rect 28534 29832 28540 29844
rect 28495 29804 28540 29832
rect 28534 29792 28540 29804
rect 28592 29792 28598 29844
rect 29730 29832 29736 29844
rect 29691 29804 29736 29832
rect 29730 29792 29736 29804
rect 29788 29792 29794 29844
rect 34885 29835 34943 29841
rect 34885 29801 34897 29835
rect 34931 29832 34943 29835
rect 35434 29832 35440 29844
rect 34931 29804 35440 29832
rect 34931 29801 34943 29804
rect 34885 29795 34943 29801
rect 35434 29792 35440 29804
rect 35492 29792 35498 29844
rect 10873 29767 10931 29773
rect 10873 29733 10885 29767
rect 10919 29764 10931 29767
rect 10919 29736 16160 29764
rect 10919 29733 10931 29736
rect 10873 29727 10931 29733
rect 8202 29656 8208 29708
rect 8260 29696 8266 29708
rect 10888 29696 10916 29727
rect 8260 29668 10916 29696
rect 8260 29656 8266 29668
rect 13538 29656 13544 29708
rect 13596 29696 13602 29708
rect 15194 29696 15200 29708
rect 13596 29668 15200 29696
rect 13596 29656 13602 29668
rect 15194 29656 15200 29668
rect 15252 29656 15258 29708
rect 15838 29656 15844 29708
rect 15896 29696 15902 29708
rect 16025 29699 16083 29705
rect 16025 29696 16037 29699
rect 15896 29668 16037 29696
rect 15896 29656 15902 29668
rect 16025 29665 16037 29668
rect 16071 29665 16083 29699
rect 16132 29696 16160 29736
rect 17310 29724 17316 29776
rect 17368 29764 17374 29776
rect 18138 29764 18144 29776
rect 17368 29736 18144 29764
rect 17368 29724 17374 29736
rect 18138 29724 18144 29736
rect 18196 29724 18202 29776
rect 18598 29724 18604 29776
rect 18656 29764 18662 29776
rect 26326 29764 26332 29776
rect 18656 29736 26332 29764
rect 18656 29724 18662 29736
rect 26326 29724 26332 29736
rect 26384 29724 26390 29776
rect 37458 29764 37464 29776
rect 27080 29736 37464 29764
rect 16132 29668 18184 29696
rect 16025 29659 16083 29665
rect 4617 29631 4675 29637
rect 4617 29597 4629 29631
rect 4663 29628 4675 29631
rect 4798 29628 4804 29640
rect 4663 29600 4804 29628
rect 4663 29597 4675 29600
rect 4617 29591 4675 29597
rect 4798 29588 4804 29600
rect 4856 29588 4862 29640
rect 9122 29628 9128 29640
rect 9083 29600 9128 29628
rect 9122 29588 9128 29600
rect 9180 29588 9186 29640
rect 11330 29628 11336 29640
rect 11291 29600 11336 29628
rect 11330 29588 11336 29600
rect 11388 29588 11394 29640
rect 13906 29628 13912 29640
rect 11900 29600 13912 29628
rect 9398 29560 9404 29572
rect 9359 29532 9404 29560
rect 9398 29520 9404 29532
rect 9456 29520 9462 29572
rect 11900 29560 11928 29600
rect 13906 29588 13912 29600
rect 13964 29588 13970 29640
rect 14458 29588 14464 29640
rect 14516 29628 14522 29640
rect 15930 29628 15936 29640
rect 14516 29600 15936 29628
rect 14516 29588 14522 29600
rect 15930 29588 15936 29600
rect 15988 29588 15994 29640
rect 18046 29628 18052 29640
rect 17434 29600 18052 29628
rect 18046 29588 18052 29600
rect 18104 29588 18110 29640
rect 18156 29628 18184 29668
rect 20622 29656 20628 29708
rect 20680 29696 20686 29708
rect 21085 29699 21143 29705
rect 21085 29696 21097 29699
rect 20680 29668 21097 29696
rect 20680 29656 20686 29668
rect 21085 29665 21097 29668
rect 21131 29665 21143 29699
rect 21085 29659 21143 29665
rect 22002 29656 22008 29708
rect 22060 29696 22066 29708
rect 24302 29696 24308 29708
rect 22060 29668 24308 29696
rect 22060 29656 22066 29668
rect 24302 29656 24308 29668
rect 24360 29656 24366 29708
rect 24762 29656 24768 29708
rect 24820 29696 24826 29708
rect 24949 29699 25007 29705
rect 24949 29696 24961 29699
rect 24820 29668 24961 29696
rect 24820 29656 24826 29668
rect 24949 29665 24961 29668
rect 24995 29665 25007 29699
rect 24949 29659 25007 29665
rect 25314 29656 25320 29708
rect 25372 29696 25378 29708
rect 25961 29699 26019 29705
rect 25961 29696 25973 29699
rect 25372 29668 25973 29696
rect 25372 29656 25378 29668
rect 25961 29665 25973 29668
rect 26007 29696 26019 29699
rect 26234 29696 26240 29708
rect 26007 29668 26240 29696
rect 26007 29665 26019 29668
rect 25961 29659 26019 29665
rect 26234 29656 26240 29668
rect 26292 29656 26298 29708
rect 18693 29631 18751 29637
rect 18693 29628 18705 29631
rect 18156 29600 18705 29628
rect 18693 29597 18705 29600
rect 18739 29597 18751 29631
rect 18693 29591 18751 29597
rect 18785 29631 18843 29637
rect 18785 29597 18797 29631
rect 18831 29628 18843 29631
rect 18966 29628 18972 29640
rect 18831 29600 18972 29628
rect 18831 29597 18843 29600
rect 18785 29591 18843 29597
rect 18966 29588 18972 29600
rect 19024 29588 19030 29640
rect 19429 29631 19487 29637
rect 19429 29597 19441 29631
rect 19475 29628 19487 29631
rect 19518 29628 19524 29640
rect 19475 29600 19524 29628
rect 19475 29597 19487 29600
rect 19429 29591 19487 29597
rect 19518 29588 19524 29600
rect 19576 29588 19582 29640
rect 20254 29628 20260 29640
rect 20215 29600 20260 29628
rect 20254 29588 20260 29600
rect 20312 29588 20318 29640
rect 20990 29628 20996 29640
rect 20951 29600 20996 29628
rect 20990 29588 20996 29600
rect 21048 29588 21054 29640
rect 21174 29588 21180 29640
rect 21232 29628 21238 29640
rect 21634 29628 21640 29640
rect 21232 29600 21640 29628
rect 21232 29588 21238 29600
rect 21634 29588 21640 29600
rect 21692 29588 21698 29640
rect 22281 29631 22339 29637
rect 22281 29597 22293 29631
rect 22327 29628 22339 29631
rect 22738 29628 22744 29640
rect 22327 29600 22744 29628
rect 22327 29597 22339 29600
rect 22281 29591 22339 29597
rect 22738 29588 22744 29600
rect 22796 29588 22802 29640
rect 22922 29628 22928 29640
rect 22883 29600 22928 29628
rect 22922 29588 22928 29600
rect 22980 29588 22986 29640
rect 23569 29631 23627 29637
rect 23569 29597 23581 29631
rect 23615 29597 23627 29631
rect 26418 29628 26424 29640
rect 23569 29591 23627 29597
rect 25884 29600 26280 29628
rect 26379 29600 26424 29628
rect 12066 29560 12072 29572
rect 10626 29532 11928 29560
rect 12027 29532 12072 29560
rect 12066 29520 12072 29532
rect 12124 29520 12130 29572
rect 13446 29520 13452 29572
rect 13504 29560 13510 29572
rect 16301 29563 16359 29569
rect 16301 29560 16313 29563
rect 13504 29532 16313 29560
rect 13504 29520 13510 29532
rect 16301 29529 16313 29532
rect 16347 29529 16359 29563
rect 21729 29563 21787 29569
rect 21729 29560 21741 29563
rect 16301 29523 16359 29529
rect 17604 29532 21741 29560
rect 11514 29452 11520 29504
rect 11572 29492 11578 29504
rect 17604 29492 17632 29532
rect 21729 29529 21741 29532
rect 21775 29529 21787 29563
rect 21729 29523 21787 29529
rect 21910 29520 21916 29572
rect 21968 29560 21974 29572
rect 23584 29560 23612 29591
rect 21968 29532 23612 29560
rect 25041 29563 25099 29569
rect 21968 29520 21974 29532
rect 25041 29529 25053 29563
rect 25087 29560 25099 29563
rect 25884 29560 25912 29600
rect 25087 29532 25912 29560
rect 26252 29560 26280 29600
rect 26418 29588 26424 29600
rect 26476 29588 26482 29640
rect 27080 29637 27108 29736
rect 37458 29724 37464 29736
rect 37516 29724 37522 29776
rect 28166 29696 28172 29708
rect 28127 29668 28172 29696
rect 28166 29656 28172 29668
rect 28224 29656 28230 29708
rect 28534 29656 28540 29708
rect 28592 29696 28598 29708
rect 28592 29668 30788 29696
rect 28592 29656 28598 29668
rect 27065 29631 27123 29637
rect 27065 29597 27077 29631
rect 27111 29597 27123 29631
rect 27065 29591 27123 29597
rect 27985 29631 28043 29637
rect 27985 29597 27997 29631
rect 28031 29628 28043 29631
rect 28442 29628 28448 29640
rect 28031 29600 28448 29628
rect 28031 29597 28043 29600
rect 27985 29591 28043 29597
rect 28442 29588 28448 29600
rect 28500 29588 28506 29640
rect 30760 29637 30788 29668
rect 34606 29656 34612 29708
rect 34664 29696 34670 29708
rect 37737 29699 37795 29705
rect 37737 29696 37749 29699
rect 34664 29668 37749 29696
rect 34664 29656 34670 29668
rect 37737 29665 37749 29668
rect 37783 29665 37795 29699
rect 37737 29659 37795 29665
rect 29917 29631 29975 29637
rect 29917 29597 29929 29631
rect 29963 29597 29975 29631
rect 29917 29591 29975 29597
rect 30745 29631 30803 29637
rect 30745 29597 30757 29631
rect 30791 29597 30803 29631
rect 30745 29591 30803 29597
rect 30837 29631 30895 29637
rect 30837 29597 30849 29631
rect 30883 29628 30895 29631
rect 35069 29631 35127 29637
rect 35069 29628 35081 29631
rect 30883 29600 35081 29628
rect 30883 29597 30895 29600
rect 30837 29591 30895 29597
rect 35069 29597 35081 29600
rect 35115 29597 35127 29631
rect 37458 29628 37464 29640
rect 37419 29600 37464 29628
rect 35069 29591 35127 29597
rect 29178 29560 29184 29572
rect 26252 29532 29184 29560
rect 25087 29529 25099 29532
rect 25041 29523 25099 29529
rect 29178 29520 29184 29532
rect 29236 29520 29242 29572
rect 11572 29464 17632 29492
rect 11572 29452 11578 29464
rect 17678 29452 17684 29504
rect 17736 29492 17742 29504
rect 17773 29495 17831 29501
rect 17773 29492 17785 29495
rect 17736 29464 17785 29492
rect 17736 29452 17742 29464
rect 17773 29461 17785 29464
rect 17819 29461 17831 29495
rect 17773 29455 17831 29461
rect 18046 29452 18052 29504
rect 18104 29492 18110 29504
rect 18782 29492 18788 29504
rect 18104 29464 18788 29492
rect 18104 29452 18110 29464
rect 18782 29452 18788 29464
rect 18840 29452 18846 29504
rect 18874 29452 18880 29504
rect 18932 29492 18938 29504
rect 19521 29495 19579 29501
rect 19521 29492 19533 29495
rect 18932 29464 19533 29492
rect 18932 29452 18938 29464
rect 19521 29461 19533 29464
rect 19567 29461 19579 29495
rect 19521 29455 19579 29461
rect 20073 29495 20131 29501
rect 20073 29461 20085 29495
rect 20119 29492 20131 29495
rect 21542 29492 21548 29504
rect 20119 29464 21548 29492
rect 20119 29461 20131 29464
rect 20073 29455 20131 29461
rect 21542 29452 21548 29464
rect 21600 29452 21606 29504
rect 23014 29492 23020 29504
rect 22975 29464 23020 29492
rect 23014 29452 23020 29464
rect 23072 29452 23078 29504
rect 23661 29495 23719 29501
rect 23661 29461 23673 29495
rect 23707 29492 23719 29495
rect 26142 29492 26148 29504
rect 23707 29464 26148 29492
rect 23707 29461 23719 29464
rect 23661 29455 23719 29461
rect 26142 29452 26148 29464
rect 26200 29452 26206 29504
rect 26510 29492 26516 29504
rect 26471 29464 26516 29492
rect 26510 29452 26516 29464
rect 26568 29452 26574 29504
rect 27154 29492 27160 29504
rect 27115 29464 27160 29492
rect 27154 29452 27160 29464
rect 27212 29452 27218 29504
rect 27522 29452 27528 29504
rect 27580 29492 27586 29504
rect 29932 29492 29960 29591
rect 37458 29588 37464 29600
rect 37516 29588 37522 29640
rect 27580 29464 29960 29492
rect 27580 29452 27586 29464
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 9398 29248 9404 29300
rect 9456 29288 9462 29300
rect 13449 29291 13507 29297
rect 13449 29288 13461 29291
rect 9456 29260 13461 29288
rect 9456 29248 9462 29260
rect 13449 29257 13461 29260
rect 13495 29288 13507 29291
rect 13538 29288 13544 29300
rect 13495 29260 13544 29288
rect 13495 29257 13507 29260
rect 13449 29251 13507 29257
rect 13538 29248 13544 29260
rect 13596 29248 13602 29300
rect 15746 29288 15752 29300
rect 14568 29260 15752 29288
rect 2774 29220 2780 29232
rect 2424 29192 2780 29220
rect 1762 29152 1768 29164
rect 1723 29124 1768 29152
rect 1762 29112 1768 29124
rect 1820 29112 1826 29164
rect 2424 29161 2452 29192
rect 2774 29180 2780 29192
rect 2832 29180 2838 29232
rect 4062 29220 4068 29232
rect 3910 29192 4068 29220
rect 4062 29180 4068 29192
rect 4120 29180 4126 29232
rect 4985 29223 5043 29229
rect 4985 29189 4997 29223
rect 5031 29220 5043 29223
rect 6178 29220 6184 29232
rect 5031 29192 6184 29220
rect 5031 29189 5043 29192
rect 4985 29183 5043 29189
rect 6178 29180 6184 29192
rect 6236 29180 6242 29232
rect 11514 29220 11520 29232
rect 10810 29192 11520 29220
rect 11514 29180 11520 29192
rect 11572 29180 11578 29232
rect 12066 29220 12072 29232
rect 11716 29192 12072 29220
rect 2409 29155 2467 29161
rect 2409 29121 2421 29155
rect 2455 29121 2467 29155
rect 2409 29115 2467 29121
rect 4433 29155 4491 29161
rect 4433 29121 4445 29155
rect 4479 29152 4491 29155
rect 7006 29152 7012 29164
rect 4479 29124 7012 29152
rect 4479 29121 4491 29124
rect 4433 29115 4491 29121
rect 7006 29112 7012 29124
rect 7064 29112 7070 29164
rect 9122 29112 9128 29164
rect 9180 29152 9186 29164
rect 9309 29155 9367 29161
rect 9309 29152 9321 29155
rect 9180 29124 9321 29152
rect 9180 29112 9186 29124
rect 9309 29121 9321 29124
rect 9355 29121 9367 29155
rect 11606 29152 11612 29164
rect 9309 29115 9367 29121
rect 10888 29124 11612 29152
rect 4890 29044 4896 29096
rect 4948 29084 4954 29096
rect 5721 29087 5779 29093
rect 5721 29084 5733 29087
rect 4948 29056 5733 29084
rect 4948 29044 4954 29056
rect 5721 29053 5733 29056
rect 5767 29053 5779 29087
rect 9324 29084 9352 29115
rect 10888 29084 10916 29124
rect 11606 29112 11612 29124
rect 11664 29152 11670 29164
rect 11716 29161 11744 29192
rect 12066 29180 12072 29192
rect 12124 29180 12130 29232
rect 14568 29220 14596 29260
rect 15746 29248 15752 29260
rect 15804 29248 15810 29300
rect 16022 29248 16028 29300
rect 16080 29288 16086 29300
rect 16080 29260 16620 29288
rect 16080 29248 16086 29260
rect 16482 29220 16488 29232
rect 14476 29192 14596 29220
rect 15962 29192 16488 29220
rect 14476 29161 14504 29192
rect 16482 29180 16488 29192
rect 16540 29180 16546 29232
rect 16592 29220 16620 29260
rect 17126 29248 17132 29300
rect 17184 29288 17190 29300
rect 21910 29288 21916 29300
rect 17184 29260 21916 29288
rect 17184 29248 17190 29260
rect 21910 29248 21916 29260
rect 21968 29248 21974 29300
rect 24854 29288 24860 29300
rect 22066 29260 24860 29288
rect 17862 29220 17868 29232
rect 16592 29192 17868 29220
rect 17862 29180 17868 29192
rect 17920 29180 17926 29232
rect 18138 29220 18144 29232
rect 18099 29192 18144 29220
rect 18138 29180 18144 29192
rect 18196 29180 18202 29232
rect 18230 29180 18236 29232
rect 18288 29220 18294 29232
rect 19334 29220 19340 29232
rect 18288 29192 19340 29220
rect 18288 29180 18294 29192
rect 19334 29180 19340 29192
rect 19392 29180 19398 29232
rect 20254 29220 20260 29232
rect 19628 29192 20260 29220
rect 11701 29155 11759 29161
rect 11701 29152 11713 29155
rect 11664 29124 11713 29152
rect 11664 29112 11670 29124
rect 11701 29121 11713 29124
rect 11747 29121 11759 29155
rect 14461 29155 14519 29161
rect 11701 29115 11759 29121
rect 11054 29084 11060 29096
rect 9324 29056 10916 29084
rect 11015 29056 11060 29084
rect 5721 29047 5779 29053
rect 11054 29044 11060 29056
rect 11112 29084 11118 29096
rect 11422 29084 11428 29096
rect 11112 29056 11428 29084
rect 11112 29044 11118 29056
rect 11422 29044 11428 29056
rect 11480 29084 11486 29096
rect 13096 29084 13124 29138
rect 14461 29121 14473 29155
rect 14507 29121 14519 29155
rect 19628 29152 19656 29192
rect 20254 29180 20260 29192
rect 20312 29180 20318 29232
rect 20533 29223 20591 29229
rect 20533 29189 20545 29223
rect 20579 29220 20591 29223
rect 21266 29220 21272 29232
rect 20579 29192 21272 29220
rect 20579 29189 20591 29192
rect 20533 29183 20591 29189
rect 21266 29180 21272 29192
rect 21324 29180 21330 29232
rect 21453 29223 21511 29229
rect 21453 29189 21465 29223
rect 21499 29220 21511 29223
rect 22066 29220 22094 29260
rect 24854 29248 24860 29260
rect 24912 29248 24918 29300
rect 24964 29260 31754 29288
rect 22922 29220 22928 29232
rect 21499 29192 22094 29220
rect 22388 29192 22928 29220
rect 21499 29189 21511 29192
rect 21453 29183 21511 29189
rect 22388 29164 22416 29192
rect 22922 29180 22928 29192
rect 22980 29180 22986 29232
rect 23014 29180 23020 29232
rect 23072 29220 23078 29232
rect 23937 29223 23995 29229
rect 23937 29220 23949 29223
rect 23072 29192 23949 29220
rect 23072 29180 23078 29192
rect 23937 29189 23949 29192
rect 23983 29189 23995 29223
rect 23937 29183 23995 29189
rect 24486 29180 24492 29232
rect 24544 29220 24550 29232
rect 24964 29220 24992 29260
rect 25516 29220 25544 29260
rect 24544 29192 24992 29220
rect 25424 29192 25544 29220
rect 24544 29180 24550 29192
rect 14461 29115 14519 29121
rect 16132 29124 17356 29152
rect 16132 29084 16160 29124
rect 11480 29056 13032 29084
rect 13096 29056 16160 29084
rect 11480 29044 11486 29056
rect 13004 29016 13032 29056
rect 14458 29016 14464 29028
rect 13004 28988 14464 29016
rect 14458 28976 14464 28988
rect 14516 28976 14522 29028
rect 16298 29016 16304 29028
rect 16224 28988 16304 29016
rect 1581 28951 1639 28957
rect 1581 28917 1593 28951
rect 1627 28948 1639 28951
rect 1854 28948 1860 28960
rect 1627 28920 1860 28948
rect 1627 28917 1639 28920
rect 1581 28911 1639 28917
rect 1854 28908 1860 28920
rect 1912 28908 1918 28960
rect 2672 28951 2730 28957
rect 2672 28917 2684 28951
rect 2718 28948 2730 28951
rect 4706 28948 4712 28960
rect 2718 28920 4712 28948
rect 2718 28917 2730 28920
rect 2672 28911 2730 28917
rect 4706 28908 4712 28920
rect 4764 28948 4770 28960
rect 5258 28948 5264 28960
rect 4764 28920 5264 28948
rect 4764 28908 4770 28920
rect 5258 28908 5264 28920
rect 5316 28908 5322 28960
rect 9572 28951 9630 28957
rect 9572 28917 9584 28951
rect 9618 28948 9630 28951
rect 10962 28948 10968 28960
rect 9618 28920 10968 28948
rect 9618 28917 9630 28920
rect 9572 28911 9630 28917
rect 10962 28908 10968 28920
rect 11020 28908 11026 28960
rect 11964 28951 12022 28957
rect 11964 28917 11976 28951
rect 12010 28948 12022 28951
rect 12066 28948 12072 28960
rect 12010 28920 12072 28948
rect 12010 28917 12022 28920
rect 11964 28911 12022 28917
rect 12066 28908 12072 28920
rect 12124 28908 12130 28960
rect 14734 28957 14740 28960
rect 14724 28951 14740 28957
rect 14724 28917 14736 28951
rect 14724 28911 14740 28917
rect 14734 28908 14740 28911
rect 14792 28908 14798 28960
rect 16224 28957 16252 28988
rect 16298 28976 16304 28988
rect 16356 29016 16362 29028
rect 16482 29016 16488 29028
rect 16356 28988 16488 29016
rect 16356 28976 16362 28988
rect 16482 28976 16488 28988
rect 16540 28976 16546 29028
rect 17328 29016 17356 29124
rect 18892 29124 19656 29152
rect 18049 29087 18107 29093
rect 18049 29053 18061 29087
rect 18095 29084 18107 29087
rect 18230 29084 18236 29096
rect 18095 29056 18236 29084
rect 18095 29053 18107 29056
rect 18049 29047 18107 29053
rect 18230 29044 18236 29056
rect 18288 29044 18294 29096
rect 18414 29084 18420 29096
rect 18375 29056 18420 29084
rect 18414 29044 18420 29056
rect 18472 29044 18478 29096
rect 18506 29044 18512 29096
rect 18564 29084 18570 29096
rect 18892 29084 18920 29124
rect 19702 29112 19708 29164
rect 19760 29152 19766 29164
rect 22370 29152 22376 29164
rect 19760 29124 20116 29152
rect 19760 29112 19766 29124
rect 18564 29056 18920 29084
rect 18564 29044 18570 29056
rect 19334 29044 19340 29096
rect 19392 29084 19398 29096
rect 19797 29087 19855 29093
rect 19797 29084 19809 29087
rect 19392 29056 19809 29084
rect 19392 29044 19398 29056
rect 19797 29053 19809 29056
rect 19843 29053 19855 29087
rect 19797 29047 19855 29053
rect 19702 29016 19708 29028
rect 17328 28988 19708 29016
rect 19702 28976 19708 28988
rect 19760 28976 19766 29028
rect 20088 29016 20116 29124
rect 21376 29124 22376 29152
rect 20254 29044 20260 29096
rect 20312 29072 20318 29096
rect 20441 29087 20499 29093
rect 20312 29044 20392 29072
rect 20441 29053 20453 29087
rect 20487 29084 20499 29087
rect 21376 29084 21404 29124
rect 22370 29112 22376 29124
rect 22428 29112 22434 29164
rect 22649 29155 22707 29161
rect 22649 29121 22661 29155
rect 22695 29121 22707 29155
rect 25038 29152 25044 29164
rect 22649 29115 22707 29121
rect 24780 29124 25044 29152
rect 20487 29056 21404 29084
rect 20487 29053 20499 29056
rect 20441 29047 20499 29053
rect 20162 29016 20168 29028
rect 20088 28988 20168 29016
rect 20162 28976 20168 28988
rect 20220 28976 20226 29028
rect 20364 29016 20392 29044
rect 22664 29016 22692 29115
rect 23845 29087 23903 29093
rect 23845 29053 23857 29087
rect 23891 29084 23903 29087
rect 23934 29084 23940 29096
rect 23891 29056 23940 29084
rect 23891 29053 23903 29056
rect 23845 29047 23903 29053
rect 23934 29044 23940 29056
rect 23992 29084 23998 29096
rect 24780 29084 24808 29124
rect 25038 29112 25044 29124
rect 25096 29112 25102 29164
rect 25424 29152 25452 29192
rect 25590 29180 25596 29232
rect 25648 29220 25654 29232
rect 25685 29223 25743 29229
rect 25685 29220 25697 29223
rect 25648 29192 25697 29220
rect 25648 29180 25654 29192
rect 25685 29189 25697 29192
rect 25731 29189 25743 29223
rect 31726 29220 31754 29260
rect 32950 29220 32956 29232
rect 31726 29192 32956 29220
rect 25685 29183 25743 29189
rect 32950 29180 32956 29192
rect 33008 29180 33014 29232
rect 25148 29124 25452 29152
rect 23992 29056 24808 29084
rect 24857 29087 24915 29093
rect 23992 29044 23998 29056
rect 24857 29053 24869 29087
rect 24903 29084 24915 29087
rect 25148 29084 25176 29124
rect 26970 29112 26976 29164
rect 27028 29152 27034 29164
rect 27157 29155 27215 29161
rect 27157 29152 27169 29155
rect 27028 29124 27169 29152
rect 27028 29112 27034 29124
rect 27157 29121 27169 29124
rect 27203 29121 27215 29155
rect 27157 29115 27215 29121
rect 24903 29056 25176 29084
rect 24903 29053 24915 29056
rect 24857 29047 24915 29053
rect 25222 29044 25228 29096
rect 25280 29084 25286 29096
rect 25593 29087 25651 29093
rect 25593 29084 25605 29087
rect 25280 29056 25605 29084
rect 25280 29044 25286 29056
rect 25593 29053 25605 29056
rect 25639 29053 25651 29087
rect 26602 29084 26608 29096
rect 26563 29056 26608 29084
rect 25593 29047 25651 29053
rect 26602 29044 26608 29056
rect 26660 29044 26666 29096
rect 27246 29084 27252 29096
rect 27207 29056 27252 29084
rect 27246 29044 27252 29056
rect 27304 29084 27310 29096
rect 27801 29087 27859 29093
rect 27801 29084 27813 29087
rect 27304 29056 27813 29084
rect 27304 29044 27310 29056
rect 27801 29053 27813 29056
rect 27847 29053 27859 29087
rect 27982 29084 27988 29096
rect 27943 29056 27988 29084
rect 27801 29047 27859 29053
rect 27982 29044 27988 29056
rect 28040 29044 28046 29096
rect 20272 28988 20392 29016
rect 20456 28988 22692 29016
rect 22741 29019 22799 29025
rect 16209 28951 16267 28957
rect 16209 28917 16221 28951
rect 16255 28948 16267 28951
rect 16255 28920 16289 28948
rect 16255 28917 16267 28920
rect 16209 28911 16267 28917
rect 18230 28908 18236 28960
rect 18288 28948 18294 28960
rect 20070 28948 20076 28960
rect 18288 28920 20076 28948
rect 18288 28908 18294 28920
rect 20070 28908 20076 28920
rect 20128 28908 20134 28960
rect 20272 28948 20300 28988
rect 20456 28948 20484 28988
rect 22741 28985 22753 29019
rect 22787 29016 22799 29019
rect 27614 29016 27620 29028
rect 22787 28988 27620 29016
rect 22787 28985 22799 28988
rect 22741 28979 22799 28985
rect 27614 28976 27620 28988
rect 27672 28976 27678 29028
rect 28442 29016 28448 29028
rect 28403 28988 28448 29016
rect 28442 28976 28448 28988
rect 28500 28976 28506 29028
rect 20272 28920 20484 28948
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 13078 28744 13084 28756
rect 9232 28716 13084 28744
rect 6917 28611 6975 28617
rect 6917 28577 6929 28611
rect 6963 28608 6975 28611
rect 9232 28608 9260 28716
rect 13078 28704 13084 28716
rect 13136 28744 13142 28756
rect 13357 28747 13415 28753
rect 13136 28716 13308 28744
rect 13136 28704 13142 28716
rect 9306 28636 9312 28688
rect 9364 28676 9370 28688
rect 13280 28676 13308 28716
rect 13357 28713 13369 28747
rect 13403 28744 13415 28747
rect 16206 28744 16212 28756
rect 13403 28716 16212 28744
rect 13403 28713 13415 28716
rect 13357 28707 13415 28713
rect 16206 28704 16212 28716
rect 16264 28704 16270 28756
rect 17310 28704 17316 28756
rect 17368 28744 17374 28756
rect 17589 28747 17647 28753
rect 17589 28744 17601 28747
rect 17368 28716 17601 28744
rect 17368 28704 17374 28716
rect 17589 28713 17601 28716
rect 17635 28713 17647 28747
rect 17589 28707 17647 28713
rect 17678 28704 17684 28756
rect 17736 28744 17742 28756
rect 17736 28716 19656 28744
rect 17736 28704 17742 28716
rect 13630 28676 13636 28688
rect 9364 28648 11744 28676
rect 13280 28648 13636 28676
rect 9364 28636 9370 28648
rect 11606 28608 11612 28620
rect 6963 28580 9260 28608
rect 11567 28580 11612 28608
rect 6963 28577 6975 28580
rect 6917 28571 6975 28577
rect 11606 28568 11612 28580
rect 11664 28568 11670 28620
rect 11716 28608 11744 28648
rect 13630 28636 13636 28648
rect 13688 28636 13694 28688
rect 13740 28648 15976 28676
rect 13740 28608 13768 28648
rect 11716 28580 13768 28608
rect 15746 28568 15752 28620
rect 15804 28608 15810 28620
rect 15841 28611 15899 28617
rect 15841 28608 15853 28611
rect 15804 28580 15853 28608
rect 15804 28568 15810 28580
rect 15841 28577 15853 28580
rect 15887 28577 15899 28611
rect 15948 28608 15976 28648
rect 18138 28636 18144 28688
rect 18196 28676 18202 28688
rect 19521 28679 19579 28685
rect 19521 28676 19533 28679
rect 18196 28648 19533 28676
rect 18196 28636 18202 28648
rect 19521 28645 19533 28648
rect 19567 28645 19579 28679
rect 19628 28676 19656 28716
rect 20346 28704 20352 28756
rect 20404 28744 20410 28756
rect 21177 28747 21235 28753
rect 21177 28744 21189 28747
rect 20404 28716 21189 28744
rect 20404 28704 20410 28716
rect 21177 28713 21189 28716
rect 21223 28713 21235 28747
rect 21177 28707 21235 28713
rect 22373 28747 22431 28753
rect 22373 28713 22385 28747
rect 22419 28744 22431 28747
rect 22646 28744 22652 28756
rect 22419 28716 22652 28744
rect 22419 28713 22431 28716
rect 22373 28707 22431 28713
rect 22646 28704 22652 28716
rect 22704 28704 22710 28756
rect 22756 28716 25360 28744
rect 22756 28676 22784 28716
rect 23842 28676 23848 28688
rect 19628 28648 22784 28676
rect 22848 28648 23848 28676
rect 19521 28639 19579 28645
rect 15948 28580 17356 28608
rect 15841 28571 15899 28577
rect 1854 28540 1860 28552
rect 1815 28512 1860 28540
rect 1854 28500 1860 28512
rect 1912 28500 1918 28552
rect 4890 28540 4896 28552
rect 4851 28512 4896 28540
rect 4890 28500 4896 28512
rect 4948 28500 4954 28552
rect 17328 28540 17356 28580
rect 17512 28580 22094 28608
rect 17512 28540 17540 28580
rect 17328 28512 17540 28540
rect 18506 28500 18512 28552
rect 18564 28540 18570 28552
rect 19429 28543 19487 28549
rect 19429 28540 19441 28543
rect 18564 28512 19441 28540
rect 18564 28500 18570 28512
rect 19429 28509 19441 28512
rect 19475 28540 19487 28543
rect 19518 28540 19524 28552
rect 19475 28512 19524 28540
rect 19475 28509 19487 28512
rect 19429 28503 19487 28509
rect 19518 28500 19524 28512
rect 19576 28500 19582 28552
rect 20073 28543 20131 28549
rect 20073 28509 20085 28543
rect 20119 28540 20131 28543
rect 20162 28540 20168 28552
rect 20119 28512 20168 28540
rect 20119 28509 20131 28512
rect 20073 28503 20131 28509
rect 20162 28500 20168 28512
rect 20220 28500 20226 28552
rect 21085 28543 21143 28549
rect 21085 28509 21097 28543
rect 21131 28542 21143 28543
rect 21174 28542 21180 28552
rect 21131 28514 21180 28542
rect 21131 28509 21143 28514
rect 21085 28503 21143 28509
rect 21174 28500 21180 28514
rect 21232 28500 21238 28552
rect 21726 28540 21732 28552
rect 21687 28512 21732 28540
rect 21726 28500 21732 28512
rect 21784 28500 21790 28552
rect 21910 28540 21916 28552
rect 21871 28512 21916 28540
rect 21910 28500 21916 28512
rect 21968 28500 21974 28552
rect 3418 28432 3424 28484
rect 3476 28472 3482 28484
rect 5169 28475 5227 28481
rect 5169 28472 5181 28475
rect 3476 28444 5181 28472
rect 3476 28432 3482 28444
rect 5169 28441 5181 28444
rect 5215 28441 5227 28475
rect 6454 28472 6460 28484
rect 6394 28444 6460 28472
rect 5169 28435 5227 28441
rect 6454 28432 6460 28444
rect 6512 28432 6518 28484
rect 11882 28472 11888 28484
rect 11843 28444 11888 28472
rect 11882 28432 11888 28444
rect 11940 28432 11946 28484
rect 16117 28475 16175 28481
rect 13110 28444 16068 28472
rect 1949 28407 2007 28413
rect 1949 28373 1961 28407
rect 1995 28404 2007 28407
rect 2130 28404 2136 28416
rect 1995 28376 2136 28404
rect 1995 28373 2007 28376
rect 1949 28367 2007 28373
rect 2130 28364 2136 28376
rect 2188 28364 2194 28416
rect 16040 28404 16068 28444
rect 16117 28441 16129 28475
rect 16163 28472 16175 28475
rect 16206 28472 16212 28484
rect 16163 28444 16212 28472
rect 16163 28441 16175 28444
rect 16117 28435 16175 28441
rect 16206 28432 16212 28444
rect 16264 28432 16270 28484
rect 18874 28472 18880 28484
rect 17342 28444 18880 28472
rect 18874 28432 18880 28444
rect 18932 28432 18938 28484
rect 19242 28432 19248 28484
rect 19300 28472 19306 28484
rect 20530 28472 20536 28484
rect 19300 28444 20536 28472
rect 19300 28432 19306 28444
rect 20530 28432 20536 28444
rect 20588 28432 20594 28484
rect 22066 28472 22094 28580
rect 22848 28472 22876 28648
rect 23842 28636 23848 28648
rect 23900 28676 23906 28688
rect 24578 28676 24584 28688
rect 23900 28648 24584 28676
rect 23900 28636 23906 28648
rect 24578 28636 24584 28648
rect 24636 28636 24642 28688
rect 25332 28676 25360 28716
rect 25406 28704 25412 28756
rect 25464 28744 25470 28756
rect 25958 28744 25964 28756
rect 25464 28716 25964 28744
rect 25464 28704 25470 28716
rect 25958 28704 25964 28716
rect 26016 28704 26022 28756
rect 27522 28744 27528 28756
rect 26252 28716 27528 28744
rect 26252 28676 26280 28716
rect 27522 28704 27528 28716
rect 27580 28704 27586 28756
rect 25332 28648 26280 28676
rect 26326 28636 26332 28688
rect 26384 28676 26390 28688
rect 26384 28648 28672 28676
rect 26384 28636 26390 28648
rect 23014 28608 23020 28620
rect 22975 28580 23020 28608
rect 23014 28568 23020 28580
rect 23072 28568 23078 28620
rect 25317 28611 25375 28617
rect 25317 28608 25329 28611
rect 23952 28580 25329 28608
rect 22066 28444 22876 28472
rect 23109 28475 23167 28481
rect 23109 28441 23121 28475
rect 23155 28472 23167 28475
rect 23952 28472 23980 28580
rect 25317 28577 25329 28580
rect 25363 28577 25375 28611
rect 25317 28571 25375 28577
rect 25961 28611 26019 28617
rect 25961 28577 25973 28611
rect 26007 28608 26019 28611
rect 26234 28608 26240 28620
rect 26007 28580 26240 28608
rect 26007 28577 26019 28580
rect 25961 28571 26019 28577
rect 26234 28568 26240 28580
rect 26292 28608 26298 28620
rect 27154 28608 27160 28620
rect 26292 28580 27160 28608
rect 26292 28568 26298 28580
rect 27154 28568 27160 28580
rect 27212 28568 27218 28620
rect 27798 28608 27804 28620
rect 27759 28580 27804 28608
rect 27798 28568 27804 28580
rect 27856 28568 27862 28620
rect 24578 28540 24584 28552
rect 24539 28512 24584 28540
rect 24578 28500 24584 28512
rect 24636 28500 24642 28552
rect 24673 28543 24731 28549
rect 24673 28509 24685 28543
rect 24719 28540 24731 28543
rect 24946 28540 24952 28552
rect 24719 28512 24952 28540
rect 24719 28509 24731 28512
rect 24673 28503 24731 28509
rect 24946 28500 24952 28512
rect 25004 28500 25010 28552
rect 25130 28500 25136 28552
rect 25188 28540 25194 28552
rect 28644 28549 28672 28648
rect 31220 28648 31754 28676
rect 31220 28549 31248 28648
rect 31297 28611 31355 28617
rect 31297 28577 31309 28611
rect 31343 28608 31355 28611
rect 31726 28608 31754 28648
rect 38102 28608 38108 28620
rect 31343 28580 31524 28608
rect 31726 28580 38108 28608
rect 31343 28577 31355 28580
rect 31297 28571 31355 28577
rect 25225 28543 25283 28549
rect 25225 28540 25237 28543
rect 25188 28512 25237 28540
rect 25188 28500 25194 28512
rect 25225 28509 25237 28512
rect 25271 28509 25283 28543
rect 25225 28503 25283 28509
rect 28629 28543 28687 28549
rect 28629 28509 28641 28543
rect 28675 28509 28687 28543
rect 28629 28503 28687 28509
rect 31205 28543 31263 28549
rect 31205 28509 31217 28543
rect 31251 28509 31263 28543
rect 31205 28503 31263 28509
rect 23155 28444 23980 28472
rect 24029 28475 24087 28481
rect 23155 28441 23167 28444
rect 23109 28435 23167 28441
rect 24029 28441 24041 28475
rect 24075 28472 24087 28475
rect 26053 28475 26111 28481
rect 24075 28444 26004 28472
rect 24075 28441 24087 28444
rect 24029 28435 24087 28441
rect 25976 28416 26004 28444
rect 26053 28441 26065 28475
rect 26099 28472 26111 28475
rect 26510 28472 26516 28484
rect 26099 28444 26516 28472
rect 26099 28441 26111 28444
rect 26053 28435 26111 28441
rect 26510 28432 26516 28444
rect 26568 28432 26574 28484
rect 26973 28475 27031 28481
rect 26973 28441 26985 28475
rect 27019 28441 27031 28475
rect 26973 28435 27031 28441
rect 17494 28404 17500 28416
rect 16040 28376 17500 28404
rect 17494 28364 17500 28376
rect 17552 28364 17558 28416
rect 19150 28364 19156 28416
rect 19208 28404 19214 28416
rect 20165 28407 20223 28413
rect 20165 28404 20177 28407
rect 19208 28376 20177 28404
rect 19208 28364 19214 28376
rect 20165 28373 20177 28376
rect 20211 28373 20223 28407
rect 20165 28367 20223 28373
rect 21082 28364 21088 28416
rect 21140 28404 21146 28416
rect 22278 28404 22284 28416
rect 21140 28376 22284 28404
rect 21140 28364 21146 28376
rect 22278 28364 22284 28376
rect 22336 28364 22342 28416
rect 22370 28364 22376 28416
rect 22428 28404 22434 28416
rect 24762 28404 24768 28416
rect 22428 28376 24768 28404
rect 22428 28364 22434 28376
rect 24762 28364 24768 28376
rect 24820 28364 24826 28416
rect 25958 28364 25964 28416
rect 26016 28404 26022 28416
rect 26988 28404 27016 28435
rect 27338 28432 27344 28484
rect 27396 28472 27402 28484
rect 27525 28475 27583 28481
rect 27525 28472 27537 28475
rect 27396 28444 27537 28472
rect 27396 28432 27402 28444
rect 27525 28441 27537 28444
rect 27571 28441 27583 28475
rect 27525 28435 27583 28441
rect 27614 28432 27620 28484
rect 27672 28472 27678 28484
rect 28721 28475 28779 28481
rect 27672 28444 27717 28472
rect 27672 28432 27678 28444
rect 28721 28441 28733 28475
rect 28767 28472 28779 28475
rect 31496 28472 31524 28580
rect 38102 28568 38108 28580
rect 38160 28568 38166 28620
rect 31941 28475 31999 28481
rect 31941 28472 31953 28475
rect 28767 28444 31432 28472
rect 31496 28444 31953 28472
rect 28767 28441 28779 28444
rect 28721 28435 28779 28441
rect 26016 28376 27016 28404
rect 31404 28404 31432 28444
rect 31941 28441 31953 28444
rect 31987 28441 31999 28475
rect 31941 28435 31999 28441
rect 32033 28475 32091 28481
rect 32033 28441 32045 28475
rect 32079 28441 32091 28475
rect 32950 28472 32956 28484
rect 32911 28444 32956 28472
rect 32033 28435 32091 28441
rect 32048 28404 32076 28435
rect 32950 28432 32956 28444
rect 33008 28432 33014 28484
rect 31404 28376 32076 28404
rect 26016 28364 26022 28376
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 9582 28160 9588 28212
rect 9640 28200 9646 28212
rect 11057 28203 11115 28209
rect 11057 28200 11069 28203
rect 9640 28172 11069 28200
rect 9640 28160 9646 28172
rect 11057 28169 11069 28172
rect 11103 28169 11115 28203
rect 20990 28200 20996 28212
rect 11057 28163 11115 28169
rect 12406 28172 20996 28200
rect 4982 28132 4988 28144
rect 4738 28104 4988 28132
rect 4982 28092 4988 28104
rect 5040 28092 5046 28144
rect 9674 28132 9680 28144
rect 9324 28104 9680 28132
rect 9324 28073 9352 28104
rect 9674 28092 9680 28104
rect 9732 28092 9738 28144
rect 11072 28132 11100 28163
rect 12406 28132 12434 28172
rect 20990 28160 20996 28172
rect 21048 28160 21054 28212
rect 21266 28200 21272 28212
rect 21227 28172 21272 28200
rect 21266 28160 21272 28172
rect 21324 28160 21330 28212
rect 22278 28160 22284 28212
rect 22336 28200 22342 28212
rect 22336 28172 24900 28200
rect 22336 28160 22342 28172
rect 18690 28132 18696 28144
rect 11072 28104 12434 28132
rect 15134 28104 18696 28132
rect 18690 28092 18696 28104
rect 18748 28092 18754 28144
rect 23198 28092 23204 28144
rect 23256 28132 23262 28144
rect 23382 28132 23388 28144
rect 23256 28104 23388 28132
rect 23256 28092 23262 28104
rect 23382 28092 23388 28104
rect 23440 28092 23446 28144
rect 24872 28132 24900 28172
rect 24946 28160 24952 28212
rect 25004 28200 25010 28212
rect 25590 28200 25596 28212
rect 25004 28172 25049 28200
rect 25551 28172 25596 28200
rect 25004 28160 25010 28172
rect 25590 28160 25596 28172
rect 25648 28160 25654 28212
rect 26142 28160 26148 28212
rect 26200 28200 26206 28212
rect 26200 28172 27384 28200
rect 26200 28160 26206 28172
rect 27356 28141 27384 28172
rect 27341 28135 27399 28141
rect 24872 28104 26372 28132
rect 9309 28067 9367 28073
rect 9309 28033 9321 28067
rect 9355 28033 9367 28067
rect 9309 28027 9367 28033
rect 10686 28024 10692 28076
rect 10744 28024 10750 28076
rect 15838 28024 15844 28076
rect 15896 28064 15902 28076
rect 15896 28036 15941 28064
rect 15896 28024 15902 28036
rect 18414 28024 18420 28076
rect 18472 28064 18478 28076
rect 19242 28064 19248 28076
rect 18472 28036 19248 28064
rect 18472 28024 18478 28036
rect 19242 28024 19248 28036
rect 19300 28024 19306 28076
rect 19889 28067 19947 28073
rect 19889 28033 19901 28067
rect 19935 28064 19947 28067
rect 20162 28064 20168 28076
rect 19935 28036 20168 28064
rect 19935 28033 19947 28036
rect 19889 28027 19947 28033
rect 20162 28024 20168 28036
rect 20220 28024 20226 28076
rect 20533 28067 20591 28073
rect 20533 28033 20545 28067
rect 20579 28033 20591 28067
rect 21174 28064 21180 28076
rect 21135 28036 21180 28064
rect 20533 28027 20591 28033
rect 2774 27956 2780 28008
rect 2832 27996 2838 28008
rect 3237 27999 3295 28005
rect 3237 27996 3249 27999
rect 2832 27968 3249 27996
rect 2832 27956 2838 27968
rect 3237 27965 3249 27968
rect 3283 27965 3295 27999
rect 3510 27996 3516 28008
rect 3471 27968 3516 27996
rect 3237 27959 3295 27965
rect 3252 27860 3280 27959
rect 3510 27956 3516 27968
rect 3568 27956 3574 28008
rect 3878 27956 3884 28008
rect 3936 27996 3942 28008
rect 4985 27999 5043 28005
rect 4985 27996 4997 27999
rect 3936 27968 4997 27996
rect 3936 27956 3942 27968
rect 4985 27965 4997 27968
rect 5031 27965 5043 27999
rect 9582 27996 9588 28008
rect 9543 27968 9588 27996
rect 4985 27959 5043 27965
rect 9582 27956 9588 27968
rect 9640 27956 9646 28008
rect 13817 27999 13875 28005
rect 13817 27965 13829 27999
rect 13863 27996 13875 27999
rect 15470 27996 15476 28008
rect 13863 27968 15476 27996
rect 13863 27965 13875 27968
rect 13817 27959 13875 27965
rect 15470 27956 15476 27968
rect 15528 27956 15534 28008
rect 15565 27999 15623 28005
rect 15565 27965 15577 27999
rect 15611 27996 15623 27999
rect 17678 27996 17684 28008
rect 15611 27968 17684 27996
rect 15611 27965 15623 27968
rect 15565 27959 15623 27965
rect 4890 27860 4896 27872
rect 3252 27832 4896 27860
rect 4890 27820 4896 27832
rect 4948 27820 4954 27872
rect 8018 27820 8024 27872
rect 8076 27860 8082 27872
rect 9398 27860 9404 27872
rect 8076 27832 9404 27860
rect 8076 27820 8082 27832
rect 9398 27820 9404 27832
rect 9456 27820 9462 27872
rect 13541 27863 13599 27869
rect 13541 27829 13553 27863
rect 13587 27860 13599 27863
rect 13722 27860 13728 27872
rect 13587 27832 13728 27860
rect 13587 27829 13599 27832
rect 13541 27823 13599 27829
rect 13722 27820 13728 27832
rect 13780 27860 13786 27872
rect 15764 27860 15792 27968
rect 17678 27956 17684 27968
rect 17736 27956 17742 28008
rect 18322 27956 18328 28008
rect 18380 27996 18386 28008
rect 19981 27999 20039 28005
rect 19981 27996 19993 27999
rect 18380 27968 19993 27996
rect 18380 27956 18386 27968
rect 19981 27965 19993 27968
rect 20027 27965 20039 27999
rect 20548 27996 20576 28027
rect 21174 28024 21180 28036
rect 21232 28024 21238 28076
rect 22646 28024 22652 28076
rect 22704 28064 22710 28076
rect 22833 28067 22891 28073
rect 22833 28064 22845 28067
rect 22704 28036 22845 28064
rect 22704 28024 22710 28036
rect 22833 28033 22845 28036
rect 22879 28033 22891 28067
rect 22833 28027 22891 28033
rect 23014 28024 23020 28076
rect 23072 28064 23078 28076
rect 23293 28067 23351 28073
rect 23293 28064 23305 28067
rect 23072 28036 23305 28064
rect 23072 28024 23078 28036
rect 23293 28033 23305 28036
rect 23339 28033 23351 28067
rect 23293 28027 23351 28033
rect 23566 28024 23572 28076
rect 23624 28064 23630 28076
rect 24872 28073 24900 28104
rect 24213 28067 24271 28073
rect 24213 28064 24225 28067
rect 23624 28036 24225 28064
rect 23624 28024 23630 28036
rect 24213 28033 24225 28036
rect 24259 28033 24271 28067
rect 24213 28027 24271 28033
rect 24857 28067 24915 28073
rect 24857 28033 24869 28067
rect 24903 28033 24915 28067
rect 24857 28027 24915 28033
rect 24946 28024 24952 28076
rect 25004 28064 25010 28076
rect 26344 28073 26372 28104
rect 27341 28101 27353 28135
rect 27387 28101 27399 28135
rect 27341 28095 27399 28101
rect 25501 28067 25559 28073
rect 25501 28064 25513 28067
rect 25004 28036 25513 28064
rect 25004 28024 25010 28036
rect 25501 28033 25513 28036
rect 25547 28033 25559 28067
rect 25501 28027 25559 28033
rect 26329 28067 26387 28073
rect 26329 28033 26341 28067
rect 26375 28033 26387 28067
rect 38286 28064 38292 28076
rect 38247 28036 38292 28064
rect 26329 28027 26387 28033
rect 38286 28024 38292 28036
rect 38344 28024 38350 28076
rect 21082 27996 21088 28008
rect 20548 27968 21088 27996
rect 19981 27959 20039 27965
rect 21082 27956 21088 27968
rect 21140 27996 21146 28008
rect 21818 27996 21824 28008
rect 21140 27968 21824 27996
rect 21140 27956 21146 27968
rect 21818 27956 21824 27968
rect 21876 27956 21882 28008
rect 22189 27999 22247 28005
rect 22189 27965 22201 27999
rect 22235 27965 22247 27999
rect 22370 27996 22376 28008
rect 22331 27968 22376 27996
rect 22189 27959 22247 27965
rect 22204 27928 22232 27959
rect 22370 27956 22376 27968
rect 22428 27956 22434 28008
rect 24302 27996 24308 28008
rect 24263 27968 24308 27996
rect 24302 27956 24308 27968
rect 24360 27956 24366 28008
rect 27249 27999 27307 28005
rect 27249 27965 27261 27999
rect 27295 27996 27307 27999
rect 27706 27996 27712 28008
rect 27295 27968 27712 27996
rect 27295 27965 27307 27968
rect 27249 27959 27307 27965
rect 27706 27956 27712 27968
rect 27764 27956 27770 28008
rect 23382 27928 23388 27940
rect 22204 27900 23388 27928
rect 23382 27888 23388 27900
rect 23440 27888 23446 27940
rect 27798 27928 27804 27940
rect 27759 27900 27804 27928
rect 27798 27888 27804 27900
rect 27856 27888 27862 27940
rect 13780 27832 15792 27860
rect 13780 27820 13786 27832
rect 17954 27820 17960 27872
rect 18012 27860 18018 27872
rect 19337 27863 19395 27869
rect 19337 27860 19349 27863
rect 18012 27832 19349 27860
rect 18012 27820 18018 27832
rect 19337 27829 19349 27832
rect 19383 27829 19395 27863
rect 20622 27860 20628 27872
rect 20583 27832 20628 27860
rect 19337 27823 19395 27829
rect 20622 27820 20628 27832
rect 20680 27820 20686 27872
rect 25774 27820 25780 27872
rect 25832 27860 25838 27872
rect 26145 27863 26203 27869
rect 26145 27860 26157 27863
rect 25832 27832 26157 27860
rect 25832 27820 25838 27832
rect 26145 27829 26157 27832
rect 26191 27829 26203 27863
rect 26145 27823 26203 27829
rect 35894 27820 35900 27872
rect 35952 27860 35958 27872
rect 38105 27863 38163 27869
rect 38105 27860 38117 27863
rect 35952 27832 38117 27860
rect 35952 27820 35958 27832
rect 38105 27829 38117 27832
rect 38151 27829 38163 27863
rect 38105 27823 38163 27829
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 2866 27616 2872 27668
rect 2924 27656 2930 27668
rect 8018 27656 8024 27668
rect 2924 27628 8024 27656
rect 2924 27616 2930 27628
rect 8018 27616 8024 27628
rect 8076 27616 8082 27668
rect 8110 27616 8116 27668
rect 8168 27656 8174 27668
rect 10578 27659 10636 27665
rect 10578 27656 10590 27659
rect 8168 27628 10590 27656
rect 8168 27616 8174 27628
rect 10578 27625 10590 27628
rect 10624 27625 10636 27659
rect 10578 27619 10636 27625
rect 10686 27616 10692 27668
rect 10744 27656 10750 27668
rect 20622 27656 20628 27668
rect 10744 27628 20628 27656
rect 10744 27616 10750 27628
rect 20622 27616 20628 27628
rect 20680 27616 20686 27668
rect 20898 27616 20904 27668
rect 20956 27656 20962 27668
rect 24946 27656 24952 27668
rect 20956 27628 24952 27656
rect 20956 27616 20962 27628
rect 24946 27616 24952 27628
rect 25004 27616 25010 27668
rect 7009 27591 7067 27597
rect 7009 27557 7021 27591
rect 7055 27588 7067 27591
rect 7098 27588 7104 27600
rect 7055 27560 7104 27588
rect 7055 27557 7067 27560
rect 7009 27551 7067 27557
rect 7098 27548 7104 27560
rect 7156 27588 7162 27600
rect 9582 27588 9588 27600
rect 7156 27560 9588 27588
rect 7156 27548 7162 27560
rect 9582 27548 9588 27560
rect 9640 27548 9646 27600
rect 18138 27588 18144 27600
rect 11716 27560 18144 27588
rect 4890 27480 4896 27532
rect 4948 27520 4954 27532
rect 5261 27523 5319 27529
rect 5261 27520 5273 27523
rect 4948 27492 5273 27520
rect 4948 27480 4954 27492
rect 5261 27489 5273 27492
rect 5307 27489 5319 27523
rect 5261 27483 5319 27489
rect 9674 27480 9680 27532
rect 9732 27520 9738 27532
rect 10321 27523 10379 27529
rect 10321 27520 10333 27523
rect 9732 27492 10333 27520
rect 9732 27480 9738 27492
rect 10321 27489 10333 27492
rect 10367 27489 10379 27523
rect 10321 27483 10379 27489
rect 1578 27452 1584 27464
rect 1539 27424 1584 27452
rect 1578 27412 1584 27424
rect 1636 27412 1642 27464
rect 11716 27438 11744 27560
rect 18138 27548 18144 27560
rect 18196 27548 18202 27600
rect 22186 27548 22192 27600
rect 22244 27588 22250 27600
rect 24026 27588 24032 27600
rect 22244 27560 24032 27588
rect 22244 27548 22250 27560
rect 24026 27548 24032 27560
rect 24084 27548 24090 27600
rect 26694 27588 26700 27600
rect 25792 27560 26700 27588
rect 11790 27480 11796 27532
rect 11848 27520 11854 27532
rect 12342 27520 12348 27532
rect 11848 27492 12348 27520
rect 11848 27480 11854 27492
rect 12342 27480 12348 27492
rect 12400 27480 12406 27532
rect 17589 27523 17647 27529
rect 17589 27489 17601 27523
rect 17635 27520 17647 27523
rect 21910 27520 21916 27532
rect 17635 27492 21916 27520
rect 17635 27489 17647 27492
rect 17589 27483 17647 27489
rect 21910 27480 21916 27492
rect 21968 27480 21974 27532
rect 22097 27523 22155 27529
rect 22097 27489 22109 27523
rect 22143 27520 22155 27523
rect 23109 27523 23167 27529
rect 22143 27492 23060 27520
rect 22143 27489 22155 27492
rect 22097 27483 22155 27489
rect 20622 27412 20628 27464
rect 20680 27452 20686 27464
rect 21177 27455 21235 27461
rect 21177 27452 21189 27455
rect 20680 27424 21189 27452
rect 20680 27412 20686 27424
rect 21177 27421 21189 27424
rect 21223 27452 21235 27455
rect 21634 27452 21640 27464
rect 21223 27424 21640 27452
rect 21223 27421 21235 27424
rect 21177 27415 21235 27421
rect 21634 27412 21640 27424
rect 21692 27412 21698 27464
rect 5537 27387 5595 27393
rect 5537 27353 5549 27387
rect 5583 27384 5595 27387
rect 5626 27384 5632 27396
rect 5583 27356 5632 27384
rect 5583 27353 5595 27356
rect 5537 27347 5595 27353
rect 5626 27344 5632 27356
rect 5684 27344 5690 27396
rect 6762 27356 6914 27384
rect 1762 27316 1768 27328
rect 1723 27288 1768 27316
rect 1762 27276 1768 27288
rect 1820 27276 1826 27328
rect 6886 27316 6914 27356
rect 12342 27344 12348 27396
rect 12400 27384 12406 27396
rect 12400 27356 17632 27384
rect 12400 27344 12406 27356
rect 13170 27316 13176 27328
rect 6886 27288 13176 27316
rect 13170 27276 13176 27288
rect 13228 27276 13234 27328
rect 17604 27316 17632 27356
rect 17678 27344 17684 27396
rect 17736 27384 17742 27396
rect 18601 27387 18659 27393
rect 17736 27356 17781 27384
rect 17736 27344 17742 27356
rect 18601 27353 18613 27387
rect 18647 27384 18659 27387
rect 18690 27384 18696 27396
rect 18647 27356 18696 27384
rect 18647 27353 18659 27356
rect 18601 27347 18659 27353
rect 18690 27344 18696 27356
rect 18748 27344 18754 27396
rect 19705 27387 19763 27393
rect 19705 27353 19717 27387
rect 19751 27353 19763 27387
rect 19705 27347 19763 27353
rect 18966 27316 18972 27328
rect 17604 27288 18972 27316
rect 18966 27276 18972 27288
rect 19024 27276 19030 27328
rect 19720 27316 19748 27347
rect 19794 27344 19800 27396
rect 19852 27384 19858 27396
rect 19852 27356 19897 27384
rect 19852 27344 19858 27356
rect 20530 27344 20536 27396
rect 20588 27384 20594 27396
rect 20717 27387 20775 27393
rect 20717 27384 20729 27387
rect 20588 27356 20729 27384
rect 20588 27344 20594 27356
rect 20717 27353 20729 27356
rect 20763 27353 20775 27387
rect 20717 27347 20775 27353
rect 22182 27387 22240 27393
rect 22182 27353 22194 27387
rect 22228 27353 22240 27387
rect 23032 27384 23060 27492
rect 23109 27489 23121 27523
rect 23155 27520 23167 27523
rect 25792 27520 25820 27560
rect 26694 27548 26700 27560
rect 26752 27548 26758 27600
rect 27982 27548 27988 27600
rect 28040 27588 28046 27600
rect 29825 27591 29883 27597
rect 29825 27588 29837 27591
rect 28040 27560 29837 27588
rect 28040 27548 28046 27560
rect 29825 27557 29837 27560
rect 29871 27557 29883 27591
rect 29825 27551 29883 27557
rect 23155 27492 25820 27520
rect 25869 27523 25927 27529
rect 23155 27489 23167 27492
rect 23109 27483 23167 27489
rect 25869 27489 25881 27523
rect 25915 27520 25927 27523
rect 26234 27520 26240 27532
rect 25915 27492 26240 27520
rect 25915 27489 25927 27492
rect 25869 27483 25927 27489
rect 26234 27480 26240 27492
rect 26292 27480 26298 27532
rect 23566 27452 23572 27464
rect 23527 27424 23572 27452
rect 23566 27412 23572 27424
rect 23624 27412 23630 27464
rect 24578 27452 24584 27464
rect 24539 27424 24584 27452
rect 24578 27412 24584 27424
rect 24636 27412 24642 27464
rect 29730 27452 29736 27464
rect 29691 27424 29736 27452
rect 29730 27412 29736 27424
rect 29788 27412 29794 27464
rect 38010 27452 38016 27464
rect 37971 27424 38016 27452
rect 38010 27412 38016 27424
rect 38068 27412 38074 27464
rect 23032 27356 25912 27384
rect 22182 27347 22240 27353
rect 20898 27316 20904 27328
rect 19720 27288 20904 27316
rect 20898 27276 20904 27288
rect 20956 27276 20962 27328
rect 21266 27316 21272 27328
rect 21227 27288 21272 27316
rect 21266 27276 21272 27288
rect 21324 27276 21330 27328
rect 22204 27316 22232 27347
rect 23661 27319 23719 27325
rect 23661 27316 23673 27319
rect 22204 27288 23673 27316
rect 23661 27285 23673 27288
rect 23707 27285 23719 27319
rect 24670 27316 24676 27328
rect 24631 27288 24676 27316
rect 23661 27279 23719 27285
rect 24670 27276 24676 27288
rect 24728 27276 24734 27328
rect 25884 27316 25912 27356
rect 25958 27344 25964 27396
rect 26016 27384 26022 27396
rect 26878 27384 26884 27396
rect 26016 27356 26061 27384
rect 26839 27356 26884 27384
rect 26016 27344 26022 27356
rect 26878 27344 26884 27356
rect 26936 27344 26942 27396
rect 28074 27316 28080 27328
rect 25884 27288 28080 27316
rect 28074 27276 28080 27288
rect 28132 27276 28138 27328
rect 38194 27316 38200 27328
rect 38155 27288 38200 27316
rect 38194 27276 38200 27288
rect 38252 27276 38258 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 1581 27115 1639 27121
rect 1581 27081 1593 27115
rect 1627 27112 1639 27115
rect 2314 27112 2320 27124
rect 1627 27084 2320 27112
rect 1627 27081 1639 27084
rect 1581 27075 1639 27081
rect 2314 27072 2320 27084
rect 2372 27072 2378 27124
rect 3326 27072 3332 27124
rect 3384 27112 3390 27124
rect 3384 27084 9444 27112
rect 3384 27072 3390 27084
rect 4525 27047 4583 27053
rect 4525 27013 4537 27047
rect 4571 27044 4583 27047
rect 4614 27044 4620 27056
rect 4571 27016 4620 27044
rect 4571 27013 4583 27016
rect 4525 27007 4583 27013
rect 4614 27004 4620 27016
rect 4672 27004 4678 27056
rect 9416 27053 9444 27084
rect 16482 27072 16488 27124
rect 16540 27112 16546 27124
rect 17405 27115 17463 27121
rect 16540 27084 16712 27112
rect 16540 27072 16546 27084
rect 9401 27047 9459 27053
rect 9401 27013 9413 27047
rect 9447 27013 9459 27047
rect 9401 27007 9459 27013
rect 10965 27047 11023 27053
rect 10965 27013 10977 27047
rect 11011 27044 11023 27047
rect 11330 27044 11336 27056
rect 11011 27016 11336 27044
rect 11011 27013 11023 27016
rect 10965 27007 11023 27013
rect 11330 27004 11336 27016
rect 11388 27004 11394 27056
rect 13722 27004 13728 27056
rect 13780 27044 13786 27056
rect 16684 27044 16712 27084
rect 17405 27081 17417 27115
rect 17451 27112 17463 27115
rect 17678 27112 17684 27124
rect 17451 27084 17684 27112
rect 17451 27081 17463 27084
rect 17405 27075 17463 27081
rect 17678 27072 17684 27084
rect 17736 27072 17742 27124
rect 20898 27112 20904 27124
rect 17788 27084 19334 27112
rect 20811 27084 20904 27112
rect 17788 27044 17816 27084
rect 18138 27044 18144 27056
rect 13780 27016 16620 27044
rect 16684 27016 17816 27044
rect 18099 27016 18144 27044
rect 13780 27004 13786 27016
rect 1762 26976 1768 26988
rect 1723 26948 1768 26976
rect 1762 26936 1768 26948
rect 1820 26936 1826 26988
rect 16482 26976 16488 26988
rect 5658 26948 5764 26976
rect 8602 26948 16488 26976
rect 5736 26920 5764 26948
rect 16482 26936 16488 26948
rect 16540 26936 16546 26988
rect 16592 26976 16620 27016
rect 18138 27004 18144 27016
rect 18196 27004 18202 27056
rect 19306 27044 19334 27084
rect 20898 27072 20904 27084
rect 20956 27112 20962 27124
rect 21726 27112 21732 27124
rect 20956 27084 21732 27112
rect 20956 27072 20962 27084
rect 21726 27072 21732 27084
rect 21784 27072 21790 27124
rect 23566 27112 23572 27124
rect 21836 27084 23572 27112
rect 21836 27044 21864 27084
rect 23566 27072 23572 27084
rect 23624 27072 23630 27124
rect 24026 27072 24032 27124
rect 24084 27112 24090 27124
rect 24394 27112 24400 27124
rect 24084 27084 24400 27112
rect 24084 27072 24090 27084
rect 24394 27072 24400 27084
rect 24452 27072 24458 27124
rect 24578 27072 24584 27124
rect 24636 27112 24642 27124
rect 34146 27112 34152 27124
rect 24636 27084 31754 27112
rect 34107 27084 34152 27112
rect 24636 27072 24642 27084
rect 19306 27016 21864 27044
rect 22097 27047 22155 27053
rect 22097 27013 22109 27047
rect 22143 27044 22155 27047
rect 22462 27044 22468 27056
rect 22143 27016 22468 27044
rect 22143 27013 22155 27016
rect 22097 27007 22155 27013
rect 22462 27004 22468 27016
rect 22520 27004 22526 27056
rect 23842 27044 23848 27056
rect 23803 27016 23848 27044
rect 23842 27004 23848 27016
rect 23900 27004 23906 27056
rect 24964 27053 24992 27084
rect 24949 27047 25007 27053
rect 24949 27013 24961 27047
rect 24995 27013 25007 27047
rect 27341 27047 27399 27053
rect 27341 27044 27353 27047
rect 24949 27007 25007 27013
rect 25056 27016 27353 27044
rect 17313 26979 17371 26985
rect 17313 26976 17325 26979
rect 16592 26948 17325 26976
rect 17313 26945 17325 26948
rect 17359 26945 17371 26979
rect 17313 26939 17371 26945
rect 17586 26936 17592 26988
rect 17644 26976 17650 26988
rect 19426 26976 19432 26988
rect 17644 26948 17908 26976
rect 17644 26936 17650 26948
rect 4249 26911 4307 26917
rect 4249 26877 4261 26911
rect 4295 26877 4307 26911
rect 4249 26871 4307 26877
rect 4264 26772 4292 26871
rect 4614 26868 4620 26920
rect 4672 26908 4678 26920
rect 4890 26908 4896 26920
rect 4672 26880 4896 26908
rect 4672 26868 4678 26880
rect 4890 26868 4896 26880
rect 4948 26868 4954 26920
rect 5074 26868 5080 26920
rect 5132 26908 5138 26920
rect 5132 26880 5580 26908
rect 5132 26868 5138 26880
rect 5552 26840 5580 26880
rect 5718 26868 5724 26920
rect 5776 26868 5782 26920
rect 6730 26868 6736 26920
rect 6788 26908 6794 26920
rect 7193 26911 7251 26917
rect 7193 26908 7205 26911
rect 6788 26880 7205 26908
rect 6788 26868 6794 26880
rect 7193 26877 7205 26880
rect 7239 26877 7251 26911
rect 7193 26871 7251 26877
rect 7469 26911 7527 26917
rect 7469 26877 7481 26911
rect 7515 26908 7527 26911
rect 7558 26908 7564 26920
rect 7515 26880 7564 26908
rect 7515 26877 7527 26880
rect 7469 26871 7527 26877
rect 7558 26868 7564 26880
rect 7616 26868 7622 26920
rect 11606 26868 11612 26920
rect 11664 26908 11670 26920
rect 17678 26908 17684 26920
rect 11664 26880 17684 26908
rect 11664 26868 11670 26880
rect 17678 26868 17684 26880
rect 17736 26868 17742 26920
rect 17880 26908 17908 26948
rect 18892 26948 19432 26976
rect 18049 26911 18107 26917
rect 18049 26908 18061 26911
rect 17880 26880 18061 26908
rect 18049 26877 18061 26880
rect 18095 26877 18107 26911
rect 18049 26871 18107 26877
rect 18892 26840 18920 26948
rect 19426 26936 19432 26948
rect 19484 26936 19490 26988
rect 19521 26979 19579 26985
rect 19521 26945 19533 26979
rect 19567 26976 19579 26979
rect 19978 26976 19984 26988
rect 19567 26948 19984 26976
rect 19567 26945 19579 26948
rect 19521 26939 19579 26945
rect 19978 26936 19984 26948
rect 20036 26936 20042 26988
rect 20162 26976 20168 26988
rect 20123 26948 20168 26976
rect 20162 26936 20168 26948
rect 20220 26936 20226 26988
rect 20809 26979 20867 26985
rect 20809 26945 20821 26979
rect 20855 26945 20867 26979
rect 20809 26939 20867 26945
rect 19061 26911 19119 26917
rect 19061 26877 19073 26911
rect 19107 26877 19119 26911
rect 20824 26908 20852 26939
rect 21634 26936 21640 26988
rect 21692 26976 21698 26988
rect 22005 26979 22063 26985
rect 22005 26976 22017 26979
rect 21692 26948 22017 26976
rect 21692 26936 21698 26948
rect 22005 26945 22017 26948
rect 22051 26976 22063 26979
rect 22649 26979 22707 26985
rect 22649 26976 22661 26979
rect 22051 26948 22661 26976
rect 22051 26945 22063 26948
rect 22005 26939 22063 26945
rect 22649 26945 22661 26948
rect 22695 26945 22707 26979
rect 22649 26939 22707 26945
rect 23382 26936 23388 26988
rect 23440 26936 23446 26988
rect 24394 26936 24400 26988
rect 24452 26976 24458 26988
rect 25056 26976 25084 27016
rect 27341 27013 27353 27016
rect 27387 27013 27399 27047
rect 31726 27044 31754 27084
rect 34146 27072 34152 27084
rect 34204 27072 34210 27124
rect 34606 27044 34612 27056
rect 31726 27016 34612 27044
rect 27341 27007 27399 27013
rect 34606 27004 34612 27016
rect 34664 27004 34670 27056
rect 25774 26976 25780 26988
rect 24452 26948 25084 26976
rect 25735 26948 25780 26976
rect 24452 26936 24458 26948
rect 25774 26936 25780 26948
rect 25832 26936 25838 26988
rect 28350 26976 28356 26988
rect 28311 26948 28356 26976
rect 28350 26936 28356 26948
rect 28408 26936 28414 26988
rect 29181 26979 29239 26985
rect 29181 26945 29193 26979
rect 29227 26976 29239 26979
rect 29227 26948 31754 26976
rect 29227 26945 29239 26948
rect 29181 26939 29239 26945
rect 22094 26908 22100 26920
rect 20824 26880 22100 26908
rect 19061 26871 19119 26877
rect 5552 26812 6914 26840
rect 4614 26772 4620 26784
rect 4264 26744 4620 26772
rect 4614 26732 4620 26744
rect 4672 26732 4678 26784
rect 5166 26732 5172 26784
rect 5224 26772 5230 26784
rect 5997 26775 6055 26781
rect 5997 26772 6009 26775
rect 5224 26744 6009 26772
rect 5224 26732 5230 26744
rect 5997 26741 6009 26744
rect 6043 26741 6055 26775
rect 6886 26772 6914 26812
rect 8588 26812 18920 26840
rect 19076 26840 19104 26871
rect 22094 26868 22100 26880
rect 22152 26868 22158 26920
rect 22462 26868 22468 26920
rect 22520 26908 22526 26920
rect 23400 26908 23428 26936
rect 23753 26911 23811 26917
rect 23753 26908 23765 26911
rect 22520 26880 23152 26908
rect 23400 26880 23765 26908
rect 22520 26868 22526 26880
rect 23124 26852 23152 26880
rect 23753 26877 23765 26880
rect 23799 26877 23811 26911
rect 23753 26871 23811 26877
rect 24029 26911 24087 26917
rect 24029 26877 24041 26911
rect 24075 26877 24087 26911
rect 24029 26871 24087 26877
rect 27249 26911 27307 26917
rect 27249 26877 27261 26911
rect 27295 26908 27307 26911
rect 29273 26911 29331 26917
rect 29273 26908 29285 26911
rect 27295 26880 29285 26908
rect 27295 26877 27307 26880
rect 27249 26871 27307 26877
rect 29273 26877 29285 26880
rect 29319 26877 29331 26911
rect 31726 26908 31754 26948
rect 31938 26936 31944 26988
rect 31996 26976 32002 26988
rect 34333 26979 34391 26985
rect 34333 26976 34345 26979
rect 31996 26948 34345 26976
rect 31996 26936 32002 26948
rect 34333 26945 34345 26948
rect 34379 26945 34391 26979
rect 34333 26939 34391 26945
rect 38102 26908 38108 26920
rect 31726 26880 38108 26908
rect 29273 26871 29331 26877
rect 19076 26812 21036 26840
rect 8588 26772 8616 26812
rect 6886 26744 8616 26772
rect 8941 26775 8999 26781
rect 5997 26735 6055 26741
rect 8941 26741 8953 26775
rect 8987 26772 8999 26775
rect 12066 26772 12072 26784
rect 8987 26744 12072 26772
rect 8987 26741 8999 26744
rect 8941 26735 8999 26741
rect 12066 26732 12072 26744
rect 12124 26732 12130 26784
rect 17126 26732 17132 26784
rect 17184 26772 17190 26784
rect 19613 26775 19671 26781
rect 19613 26772 19625 26775
rect 17184 26744 19625 26772
rect 17184 26732 17190 26744
rect 19613 26741 19625 26744
rect 19659 26741 19671 26775
rect 19613 26735 19671 26741
rect 19978 26732 19984 26784
rect 20036 26772 20042 26784
rect 20257 26775 20315 26781
rect 20257 26772 20269 26775
rect 20036 26744 20269 26772
rect 20036 26732 20042 26744
rect 20257 26741 20269 26744
rect 20303 26741 20315 26775
rect 21008 26772 21036 26812
rect 21082 26800 21088 26852
rect 21140 26840 21146 26852
rect 22741 26843 22799 26849
rect 22741 26840 22753 26843
rect 21140 26812 22753 26840
rect 21140 26800 21146 26812
rect 22741 26809 22753 26812
rect 22787 26809 22799 26843
rect 22741 26803 22799 26809
rect 23106 26800 23112 26852
rect 23164 26840 23170 26852
rect 24044 26840 24072 26871
rect 38102 26868 38108 26880
rect 38160 26868 38166 26920
rect 23164 26812 24072 26840
rect 23164 26800 23170 26812
rect 24762 26800 24768 26852
rect 24820 26840 24826 26852
rect 25593 26843 25651 26849
rect 25593 26840 25605 26843
rect 24820 26812 25605 26840
rect 24820 26800 24826 26812
rect 25593 26809 25605 26812
rect 25639 26809 25651 26843
rect 25593 26803 25651 26809
rect 27706 26800 27712 26852
rect 27764 26840 27770 26852
rect 27801 26843 27859 26849
rect 27801 26840 27813 26843
rect 27764 26812 27813 26840
rect 27764 26800 27770 26812
rect 27801 26809 27813 26812
rect 27847 26809 27859 26843
rect 27801 26803 27859 26809
rect 24486 26772 24492 26784
rect 21008 26744 24492 26772
rect 20257 26735 20315 26741
rect 24486 26732 24492 26744
rect 24544 26732 24550 26784
rect 25038 26772 25044 26784
rect 24999 26744 25044 26772
rect 25038 26732 25044 26744
rect 25096 26732 25102 26784
rect 27890 26732 27896 26784
rect 27948 26772 27954 26784
rect 28445 26775 28503 26781
rect 28445 26772 28457 26775
rect 27948 26744 28457 26772
rect 27948 26732 27954 26744
rect 28445 26741 28457 26744
rect 28491 26741 28503 26775
rect 28445 26735 28503 26741
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 2958 26528 2964 26580
rect 3016 26568 3022 26580
rect 3510 26568 3516 26580
rect 3016 26540 3516 26568
rect 3016 26528 3022 26540
rect 3510 26528 3516 26540
rect 3568 26568 3574 26580
rect 8481 26571 8539 26577
rect 8481 26568 8493 26571
rect 3568 26540 8493 26568
rect 3568 26528 3574 26540
rect 8481 26537 8493 26540
rect 8527 26568 8539 26571
rect 8938 26568 8944 26580
rect 8527 26540 8944 26568
rect 8527 26537 8539 26540
rect 8481 26531 8539 26537
rect 8938 26528 8944 26540
rect 8996 26528 9002 26580
rect 16012 26571 16070 26577
rect 16012 26537 16024 26571
rect 16058 26568 16070 26571
rect 17770 26568 17776 26580
rect 16058 26540 17776 26568
rect 16058 26537 16070 26540
rect 16012 26531 16070 26537
rect 17770 26528 17776 26540
rect 17828 26528 17834 26580
rect 17862 26528 17868 26580
rect 17920 26568 17926 26580
rect 18785 26571 18843 26577
rect 18785 26568 18797 26571
rect 17920 26540 18797 26568
rect 17920 26528 17926 26540
rect 18785 26537 18797 26540
rect 18831 26537 18843 26571
rect 18785 26531 18843 26537
rect 20346 26528 20352 26580
rect 20404 26568 20410 26580
rect 21082 26568 21088 26580
rect 20404 26540 21088 26568
rect 20404 26528 20410 26540
rect 21082 26528 21088 26540
rect 21140 26528 21146 26580
rect 23842 26528 23848 26580
rect 23900 26568 23906 26580
rect 25041 26571 25099 26577
rect 25041 26568 25053 26571
rect 23900 26540 25053 26568
rect 23900 26528 23906 26540
rect 25041 26537 25053 26540
rect 25087 26537 25099 26571
rect 25041 26531 25099 26537
rect 25685 26571 25743 26577
rect 25685 26537 25697 26571
rect 25731 26568 25743 26571
rect 25958 26568 25964 26580
rect 25731 26540 25964 26568
rect 25731 26537 25743 26540
rect 25685 26531 25743 26537
rect 25958 26528 25964 26540
rect 26016 26528 26022 26580
rect 29454 26568 29460 26580
rect 26344 26540 29460 26568
rect 13262 26460 13268 26512
rect 13320 26500 13326 26512
rect 13725 26503 13783 26509
rect 13725 26500 13737 26503
rect 13320 26472 13737 26500
rect 13320 26460 13326 26472
rect 13725 26469 13737 26472
rect 13771 26469 13783 26503
rect 17788 26500 17816 26528
rect 19426 26500 19432 26512
rect 17788 26472 19432 26500
rect 13725 26463 13783 26469
rect 19426 26460 19432 26472
rect 19484 26460 19490 26512
rect 19518 26460 19524 26512
rect 19576 26500 19582 26512
rect 24670 26500 24676 26512
rect 19576 26472 24676 26500
rect 19576 26460 19582 26472
rect 24670 26460 24676 26472
rect 24728 26460 24734 26512
rect 2130 26432 2136 26444
rect 2091 26404 2136 26432
rect 2130 26392 2136 26404
rect 2188 26392 2194 26444
rect 7006 26432 7012 26444
rect 6967 26404 7012 26432
rect 7006 26392 7012 26404
rect 7064 26392 7070 26444
rect 21266 26432 21272 26444
rect 13372 26404 21272 26432
rect 6730 26364 6736 26376
rect 6691 26336 6736 26364
rect 6730 26324 6736 26336
rect 6788 26324 6794 26376
rect 11606 26364 11612 26376
rect 8142 26336 11612 26364
rect 11606 26324 11612 26336
rect 11664 26324 11670 26376
rect 11698 26324 11704 26376
rect 11756 26364 11762 26376
rect 11977 26367 12035 26373
rect 11977 26364 11989 26367
rect 11756 26336 11989 26364
rect 11756 26324 11762 26336
rect 11977 26333 11989 26336
rect 12023 26333 12035 26367
rect 13372 26350 13400 26404
rect 21266 26392 21272 26404
rect 21324 26392 21330 26444
rect 26344 26441 26372 26540
rect 29454 26528 29460 26540
rect 29512 26528 29518 26580
rect 31938 26568 31944 26580
rect 31899 26540 31944 26568
rect 31938 26528 31944 26540
rect 31996 26528 32002 26580
rect 38102 26568 38108 26580
rect 38063 26540 38108 26568
rect 38102 26528 38108 26540
rect 38160 26528 38166 26580
rect 26881 26503 26939 26509
rect 26881 26469 26893 26503
rect 26927 26500 26939 26503
rect 27798 26500 27804 26512
rect 26927 26472 27804 26500
rect 26927 26469 26939 26472
rect 26881 26463 26939 26469
rect 27798 26460 27804 26472
rect 27856 26500 27862 26512
rect 33226 26500 33232 26512
rect 27856 26472 33232 26500
rect 27856 26460 27862 26472
rect 33226 26460 33232 26472
rect 33284 26460 33290 26512
rect 23201 26435 23259 26441
rect 23201 26401 23213 26435
rect 23247 26432 23259 26435
rect 26329 26435 26387 26441
rect 23247 26404 26188 26432
rect 23247 26401 23259 26404
rect 23201 26395 23259 26401
rect 15746 26364 15752 26376
rect 15707 26336 15752 26364
rect 11977 26327 12035 26333
rect 15746 26324 15752 26336
rect 15804 26324 15810 26376
rect 17126 26324 17132 26376
rect 17184 26324 17190 26376
rect 17586 26324 17592 26376
rect 17644 26364 17650 26376
rect 18693 26367 18751 26373
rect 17644 26336 18460 26364
rect 17644 26324 17650 26336
rect 2225 26299 2283 26305
rect 2225 26265 2237 26299
rect 2271 26296 2283 26299
rect 3050 26296 3056 26308
rect 2271 26268 3056 26296
rect 2271 26265 2283 26268
rect 2225 26259 2283 26265
rect 3050 26256 3056 26268
rect 3108 26256 3114 26308
rect 3145 26299 3203 26305
rect 3145 26265 3157 26299
rect 3191 26296 3203 26299
rect 5074 26296 5080 26308
rect 3191 26268 5080 26296
rect 3191 26265 3203 26268
rect 3145 26259 3203 26265
rect 5074 26256 5080 26268
rect 5132 26256 5138 26308
rect 8386 26256 8392 26308
rect 8444 26296 8450 26308
rect 12250 26296 12256 26308
rect 8444 26268 8616 26296
rect 12211 26268 12256 26296
rect 8444 26256 8450 26268
rect 8588 26228 8616 26268
rect 12250 26256 12256 26268
rect 12308 26256 12314 26308
rect 17770 26296 17776 26308
rect 17731 26268 17776 26296
rect 17770 26256 17776 26268
rect 17828 26256 17834 26308
rect 18432 26296 18460 26336
rect 18693 26333 18705 26367
rect 18739 26364 18751 26367
rect 19058 26364 19064 26376
rect 18739 26336 19064 26364
rect 18739 26333 18751 26336
rect 18693 26327 18751 26333
rect 19058 26324 19064 26336
rect 19116 26364 19122 26376
rect 19242 26364 19248 26376
rect 19116 26336 19248 26364
rect 19116 26324 19122 26336
rect 19242 26324 19248 26336
rect 19300 26324 19306 26376
rect 20806 26364 20812 26376
rect 20456 26336 20812 26364
rect 19518 26296 19524 26308
rect 18432 26268 19380 26296
rect 19479 26268 19524 26296
rect 12986 26228 12992 26240
rect 8588 26200 12992 26228
rect 12986 26188 12992 26200
rect 13044 26188 13050 26240
rect 15102 26188 15108 26240
rect 15160 26228 15166 26240
rect 18874 26228 18880 26240
rect 15160 26200 18880 26228
rect 15160 26188 15166 26200
rect 18874 26188 18880 26200
rect 18932 26188 18938 26240
rect 19352 26228 19380 26268
rect 19518 26256 19524 26268
rect 19576 26256 19582 26308
rect 19613 26299 19671 26305
rect 19613 26265 19625 26299
rect 19659 26296 19671 26299
rect 20456 26296 20484 26336
rect 20806 26324 20812 26336
rect 20864 26324 20870 26376
rect 23106 26364 23112 26376
rect 23067 26336 23112 26364
rect 23106 26324 23112 26336
rect 23164 26324 23170 26376
rect 23750 26364 23756 26376
rect 23711 26336 23756 26364
rect 23750 26324 23756 26336
rect 23808 26324 23814 26376
rect 23845 26367 23903 26373
rect 23845 26333 23857 26367
rect 23891 26364 23903 26367
rect 24394 26364 24400 26376
rect 23891 26336 24400 26364
rect 23891 26333 23903 26336
rect 23845 26327 23903 26333
rect 24394 26324 24400 26336
rect 24452 26324 24458 26376
rect 24949 26367 25007 26373
rect 24949 26364 24961 26367
rect 24504 26336 24961 26364
rect 19659 26268 20484 26296
rect 19659 26265 19671 26268
rect 19613 26259 19671 26265
rect 20530 26256 20536 26308
rect 20588 26296 20594 26308
rect 20588 26268 20681 26296
rect 20588 26256 20594 26268
rect 21082 26256 21088 26308
rect 21140 26296 21146 26308
rect 21140 26268 23428 26296
rect 21140 26256 21146 26268
rect 20548 26228 20576 26256
rect 19352 26200 20576 26228
rect 21450 26188 21456 26240
rect 21508 26228 21514 26240
rect 23290 26228 23296 26240
rect 21508 26200 23296 26228
rect 21508 26188 21514 26200
rect 23290 26188 23296 26200
rect 23348 26188 23354 26240
rect 23400 26228 23428 26268
rect 24504 26228 24532 26336
rect 24949 26333 24961 26336
rect 24995 26364 25007 26367
rect 25406 26364 25412 26376
rect 24995 26336 25412 26364
rect 24995 26333 25007 26336
rect 24949 26327 25007 26333
rect 25406 26324 25412 26336
rect 25464 26324 25470 26376
rect 25593 26367 25651 26373
rect 25593 26333 25605 26367
rect 25639 26364 25651 26367
rect 25866 26364 25872 26376
rect 25639 26336 25872 26364
rect 25639 26333 25651 26336
rect 25593 26327 25651 26333
rect 25866 26324 25872 26336
rect 25924 26324 25930 26376
rect 23400 26200 24532 26228
rect 26160 26228 26188 26404
rect 26329 26401 26341 26435
rect 26375 26401 26387 26435
rect 26329 26395 26387 26401
rect 31846 26364 31852 26376
rect 31807 26336 31852 26364
rect 31846 26324 31852 26336
rect 31904 26324 31910 26376
rect 38286 26364 38292 26376
rect 38247 26336 38292 26364
rect 38286 26324 38292 26336
rect 38344 26324 38350 26376
rect 26418 26296 26424 26308
rect 26379 26268 26424 26296
rect 26418 26256 26424 26268
rect 26476 26256 26482 26308
rect 32582 26296 32588 26308
rect 28966 26268 32444 26296
rect 32543 26268 32588 26296
rect 28966 26228 28994 26268
rect 26160 26200 28994 26228
rect 32416 26228 32444 26268
rect 32582 26256 32588 26268
rect 32640 26256 32646 26308
rect 32677 26299 32735 26305
rect 32677 26265 32689 26299
rect 32723 26265 32735 26299
rect 33226 26296 33232 26308
rect 33187 26268 33232 26296
rect 32677 26259 32735 26265
rect 32692 26228 32720 26259
rect 33226 26256 33232 26268
rect 33284 26256 33290 26308
rect 32416 26200 32720 26228
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 3050 26024 3056 26036
rect 3011 25996 3056 26024
rect 3050 25984 3056 25996
rect 3108 25984 3114 26036
rect 5353 26027 5411 26033
rect 5353 26024 5365 26027
rect 3160 25996 5365 26024
rect 1946 25916 1952 25968
rect 2004 25956 2010 25968
rect 3160 25956 3188 25996
rect 5353 25993 5365 25996
rect 5399 25993 5411 26027
rect 17954 26024 17960 26036
rect 5353 25987 5411 25993
rect 12360 25996 17960 26024
rect 12360 25956 12388 25996
rect 17954 25984 17960 25996
rect 18012 25984 18018 26036
rect 18138 25984 18144 26036
rect 18196 26024 18202 26036
rect 19705 26027 19763 26033
rect 19705 26024 19717 26027
rect 18196 25996 19717 26024
rect 18196 25984 18202 25996
rect 19705 25993 19717 25996
rect 19751 25993 19763 26027
rect 19705 25987 19763 25993
rect 21174 25984 21180 26036
rect 21232 25984 21238 26036
rect 22189 26027 22247 26033
rect 22189 25993 22201 26027
rect 22235 26024 22247 26027
rect 26418 26024 26424 26036
rect 22235 25996 26424 26024
rect 22235 25993 22247 25996
rect 22189 25987 22247 25993
rect 26418 25984 26424 25996
rect 26476 25984 26482 26036
rect 32582 25984 32588 26036
rect 32640 26024 32646 26036
rect 32677 26027 32735 26033
rect 32677 26024 32689 26027
rect 32640 25996 32689 26024
rect 32640 25984 32646 25996
rect 32677 25993 32689 25996
rect 32723 25993 32735 26027
rect 32677 25987 32735 25993
rect 2004 25928 3188 25956
rect 10810 25928 12388 25956
rect 2004 25916 2010 25928
rect 14642 25916 14648 25968
rect 14700 25956 14706 25968
rect 17218 25956 17224 25968
rect 14700 25928 17224 25956
rect 14700 25916 14706 25928
rect 17218 25916 17224 25928
rect 17276 25916 17282 25968
rect 19150 25956 19156 25968
rect 18354 25928 19156 25956
rect 19150 25916 19156 25928
rect 19208 25916 19214 25968
rect 21192 25956 21220 25984
rect 22370 25956 22376 25968
rect 19536 25928 22376 25956
rect 2958 25888 2964 25900
rect 2919 25860 2964 25888
rect 2958 25848 2964 25860
rect 3016 25848 3022 25900
rect 4982 25848 4988 25900
rect 5040 25848 5046 25900
rect 7926 25888 7932 25900
rect 7887 25860 7932 25888
rect 7926 25848 7932 25860
rect 7984 25848 7990 25900
rect 3605 25823 3663 25829
rect 3605 25789 3617 25823
rect 3651 25820 3663 25823
rect 3878 25820 3884 25832
rect 3651 25792 3740 25820
rect 3839 25792 3884 25820
rect 3651 25789 3663 25792
rect 3605 25783 3663 25789
rect 3712 25684 3740 25792
rect 3878 25780 3884 25792
rect 3936 25780 3942 25832
rect 6730 25780 6736 25832
rect 6788 25820 6794 25832
rect 8386 25820 8392 25832
rect 6788 25792 8392 25820
rect 6788 25780 6794 25792
rect 8386 25780 8392 25792
rect 8444 25820 8450 25832
rect 8665 25823 8723 25829
rect 8665 25820 8677 25823
rect 8444 25792 8677 25820
rect 8444 25780 8450 25792
rect 8665 25789 8677 25792
rect 8711 25820 8723 25823
rect 9122 25820 9128 25832
rect 8711 25792 9128 25820
rect 8711 25789 8723 25792
rect 8665 25783 8723 25789
rect 9122 25780 9128 25792
rect 9180 25820 9186 25832
rect 9309 25823 9367 25829
rect 9309 25820 9321 25823
rect 9180 25792 9321 25820
rect 9180 25780 9186 25792
rect 9309 25789 9321 25792
rect 9355 25789 9367 25823
rect 9309 25783 9367 25789
rect 9585 25823 9643 25829
rect 9585 25789 9597 25823
rect 9631 25820 9643 25823
rect 10962 25820 10968 25832
rect 9631 25792 10968 25820
rect 9631 25789 9643 25792
rect 9585 25783 9643 25789
rect 10962 25780 10968 25792
rect 11020 25780 11026 25832
rect 11698 25820 11704 25832
rect 11659 25792 11704 25820
rect 11698 25780 11704 25792
rect 11756 25780 11762 25832
rect 11977 25823 12035 25829
rect 11977 25820 11989 25823
rect 11808 25792 11989 25820
rect 10870 25712 10876 25764
rect 10928 25752 10934 25764
rect 11808 25752 11836 25792
rect 11977 25789 11989 25792
rect 12023 25820 12035 25823
rect 12023 25792 13032 25820
rect 12023 25789 12035 25792
rect 11977 25783 12035 25789
rect 10928 25724 11836 25752
rect 10928 25712 10934 25724
rect 4614 25684 4620 25696
rect 3712 25656 4620 25684
rect 4614 25644 4620 25656
rect 4672 25644 4678 25696
rect 11054 25684 11060 25696
rect 11015 25656 11060 25684
rect 11054 25644 11060 25656
rect 11112 25644 11118 25696
rect 13004 25684 13032 25792
rect 13096 25752 13124 25874
rect 14826 25848 14832 25900
rect 14884 25888 14890 25900
rect 16758 25888 16764 25900
rect 14884 25860 16764 25888
rect 14884 25848 14890 25860
rect 16758 25848 16764 25860
rect 16816 25848 16822 25900
rect 18598 25848 18604 25900
rect 18656 25888 18662 25900
rect 19536 25888 19564 25928
rect 22370 25916 22376 25928
rect 22428 25916 22434 25968
rect 18656 25860 19564 25888
rect 19613 25891 19671 25897
rect 18656 25848 18662 25860
rect 19613 25857 19625 25891
rect 19659 25857 19671 25891
rect 19613 25851 19671 25857
rect 13446 25820 13452 25832
rect 13407 25792 13452 25820
rect 13446 25780 13452 25792
rect 13504 25780 13510 25832
rect 15746 25780 15752 25832
rect 15804 25820 15810 25832
rect 16853 25823 16911 25829
rect 16853 25820 16865 25823
rect 15804 25792 16865 25820
rect 15804 25780 15810 25792
rect 16853 25789 16865 25792
rect 16899 25789 16911 25823
rect 17126 25820 17132 25832
rect 17087 25792 17132 25820
rect 16853 25783 16911 25789
rect 17126 25780 17132 25792
rect 17184 25780 17190 25832
rect 17218 25780 17224 25832
rect 17276 25820 17282 25832
rect 19628 25820 19656 25851
rect 20162 25848 20168 25900
rect 20220 25888 20226 25900
rect 20257 25891 20315 25897
rect 20257 25888 20269 25891
rect 20220 25860 20269 25888
rect 20220 25848 20226 25860
rect 20257 25857 20269 25860
rect 20303 25888 20315 25891
rect 21174 25888 21180 25900
rect 20303 25860 21180 25888
rect 20303 25857 20315 25860
rect 20257 25851 20315 25857
rect 21174 25848 21180 25860
rect 21232 25848 21238 25900
rect 21269 25891 21327 25897
rect 21269 25857 21281 25891
rect 21315 25888 21327 25891
rect 21358 25888 21364 25900
rect 21315 25860 21364 25888
rect 21315 25857 21327 25860
rect 21269 25851 21327 25857
rect 21358 25848 21364 25860
rect 21416 25848 21422 25900
rect 21634 25848 21640 25900
rect 21692 25888 21698 25900
rect 22097 25891 22155 25897
rect 22097 25888 22109 25891
rect 21692 25860 22109 25888
rect 21692 25848 21698 25860
rect 22097 25857 22109 25860
rect 22143 25857 22155 25891
rect 22097 25851 22155 25857
rect 22186 25848 22192 25900
rect 22244 25888 22250 25900
rect 22925 25891 22983 25897
rect 22925 25888 22937 25891
rect 22244 25860 22937 25888
rect 22244 25848 22250 25860
rect 22925 25857 22937 25860
rect 22971 25857 22983 25891
rect 22925 25851 22983 25857
rect 23290 25848 23296 25900
rect 23348 25888 23354 25900
rect 23385 25891 23443 25897
rect 23385 25888 23397 25891
rect 23348 25860 23397 25888
rect 23348 25848 23354 25860
rect 23385 25857 23397 25860
rect 23431 25888 23443 25891
rect 23934 25888 23940 25900
rect 23431 25860 23940 25888
rect 23431 25857 23443 25860
rect 23385 25851 23443 25857
rect 23934 25848 23940 25860
rect 23992 25848 23998 25900
rect 28258 25888 28264 25900
rect 28219 25860 28264 25888
rect 28258 25848 28264 25860
rect 28316 25848 28322 25900
rect 29089 25891 29147 25897
rect 29089 25857 29101 25891
rect 29135 25857 29147 25891
rect 29089 25851 29147 25857
rect 29181 25891 29239 25897
rect 29181 25857 29193 25891
rect 29227 25888 29239 25891
rect 31205 25891 31263 25897
rect 31205 25888 31217 25891
rect 29227 25860 31217 25888
rect 29227 25857 29239 25860
rect 29181 25851 29239 25857
rect 31205 25857 31217 25860
rect 31251 25857 31263 25891
rect 31205 25851 31263 25857
rect 17276 25792 19656 25820
rect 17276 25780 17282 25792
rect 20806 25780 20812 25832
rect 20864 25820 20870 25832
rect 23477 25823 23535 25829
rect 23477 25820 23489 25823
rect 20864 25792 23489 25820
rect 20864 25780 20870 25792
rect 23477 25789 23489 25792
rect 23523 25789 23535 25823
rect 29104 25820 29132 25851
rect 29914 25820 29920 25832
rect 29104 25792 29224 25820
rect 29875 25792 29920 25820
rect 23477 25783 23535 25789
rect 29196 25764 29224 25792
rect 29914 25780 29920 25792
rect 29972 25780 29978 25832
rect 30098 25820 30104 25832
rect 30059 25792 30104 25820
rect 30098 25780 30104 25792
rect 30156 25780 30162 25832
rect 30466 25780 30472 25832
rect 30524 25820 30530 25832
rect 31021 25823 31079 25829
rect 31021 25820 31033 25823
rect 30524 25792 31033 25820
rect 30524 25780 30530 25792
rect 31021 25789 31033 25792
rect 31067 25789 31079 25823
rect 31021 25783 31079 25789
rect 20990 25752 20996 25764
rect 13096 25724 16988 25752
rect 16666 25684 16672 25696
rect 13004 25656 16672 25684
rect 16666 25644 16672 25656
rect 16724 25644 16730 25696
rect 16960 25684 16988 25724
rect 18524 25724 20996 25752
rect 18524 25684 18552 25724
rect 20990 25712 20996 25724
rect 21048 25712 21054 25764
rect 22741 25755 22799 25761
rect 22741 25721 22753 25755
rect 22787 25752 22799 25755
rect 29086 25752 29092 25764
rect 22787 25724 29092 25752
rect 22787 25721 22799 25724
rect 22741 25715 22799 25721
rect 29086 25712 29092 25724
rect 29144 25712 29150 25764
rect 29178 25712 29184 25764
rect 29236 25712 29242 25764
rect 31846 25752 31852 25764
rect 31726 25724 31852 25752
rect 16960 25656 18552 25684
rect 18598 25644 18604 25696
rect 18656 25684 18662 25696
rect 18656 25656 18701 25684
rect 18656 25644 18662 25656
rect 19426 25644 19432 25696
rect 19484 25684 19490 25696
rect 20349 25687 20407 25693
rect 20349 25684 20361 25687
rect 19484 25656 20361 25684
rect 19484 25644 19490 25656
rect 20349 25653 20361 25656
rect 20395 25653 20407 25687
rect 21358 25684 21364 25696
rect 21319 25656 21364 25684
rect 20349 25647 20407 25653
rect 21358 25644 21364 25656
rect 21416 25644 21422 25696
rect 28077 25687 28135 25693
rect 28077 25653 28089 25687
rect 28123 25684 28135 25687
rect 28534 25684 28540 25696
rect 28123 25656 28540 25684
rect 28123 25653 28135 25656
rect 28077 25647 28135 25653
rect 28534 25644 28540 25656
rect 28592 25644 28598 25696
rect 30561 25687 30619 25693
rect 30561 25653 30573 25687
rect 30607 25684 30619 25687
rect 31389 25687 31447 25693
rect 31389 25684 31401 25687
rect 30607 25656 31401 25684
rect 30607 25653 30619 25656
rect 30561 25647 30619 25653
rect 31389 25653 31401 25656
rect 31435 25684 31447 25687
rect 31726 25684 31754 25724
rect 31846 25712 31852 25724
rect 31904 25712 31910 25764
rect 31435 25656 31754 25684
rect 31435 25653 31447 25656
rect 31389 25647 31447 25653
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 10870 25480 10876 25492
rect 10831 25452 10876 25480
rect 10870 25440 10876 25452
rect 10928 25440 10934 25492
rect 13722 25480 13728 25492
rect 11900 25452 13728 25480
rect 6730 25344 6736 25356
rect 6691 25316 6736 25344
rect 6730 25304 6736 25316
rect 6788 25304 6794 25356
rect 7009 25347 7067 25353
rect 7009 25313 7021 25347
rect 7055 25344 7067 25347
rect 9122 25344 9128 25356
rect 7055 25316 8984 25344
rect 9083 25316 9128 25344
rect 7055 25313 7067 25316
rect 7009 25307 7067 25313
rect 1670 25276 1676 25288
rect 1631 25248 1676 25276
rect 1670 25236 1676 25248
rect 1728 25236 1734 25288
rect 1857 25211 1915 25217
rect 1857 25177 1869 25211
rect 1903 25208 1915 25211
rect 2682 25208 2688 25220
rect 1903 25180 2688 25208
rect 1903 25177 1915 25180
rect 1857 25171 1915 25177
rect 2682 25168 2688 25180
rect 2740 25168 2746 25220
rect 8018 25168 8024 25220
rect 8076 25168 8082 25220
rect 3970 25100 3976 25152
rect 4028 25140 4034 25152
rect 8481 25143 8539 25149
rect 8481 25140 8493 25143
rect 4028 25112 8493 25140
rect 4028 25100 4034 25112
rect 8481 25109 8493 25112
rect 8527 25140 8539 25143
rect 8662 25140 8668 25152
rect 8527 25112 8668 25140
rect 8527 25109 8539 25112
rect 8481 25103 8539 25109
rect 8662 25100 8668 25112
rect 8720 25100 8726 25152
rect 8956 25140 8984 25316
rect 9122 25304 9128 25316
rect 9180 25304 9186 25356
rect 9401 25347 9459 25353
rect 9401 25313 9413 25347
rect 9447 25344 9459 25347
rect 11900 25344 11928 25452
rect 13722 25440 13728 25452
rect 13780 25440 13786 25492
rect 19334 25480 19340 25492
rect 15304 25452 19340 25480
rect 9447 25316 11928 25344
rect 12069 25347 12127 25353
rect 9447 25313 9459 25316
rect 9401 25307 9459 25313
rect 12069 25313 12081 25347
rect 12115 25344 12127 25347
rect 14826 25344 14832 25356
rect 12115 25316 14832 25344
rect 12115 25313 12127 25316
rect 12069 25307 12127 25313
rect 14826 25304 14832 25316
rect 14884 25304 14890 25356
rect 10502 25236 10508 25288
rect 10560 25236 10566 25288
rect 11790 25276 11796 25288
rect 11751 25248 11796 25276
rect 11790 25236 11796 25248
rect 11848 25236 11854 25288
rect 15304 25276 15332 25452
rect 19334 25440 19340 25452
rect 19392 25440 19398 25492
rect 19518 25440 19524 25492
rect 19576 25480 19582 25492
rect 20530 25480 20536 25492
rect 19576 25452 20536 25480
rect 19576 25440 19582 25452
rect 20530 25440 20536 25452
rect 20588 25440 20594 25492
rect 21913 25483 21971 25489
rect 21913 25449 21925 25483
rect 21959 25480 21971 25483
rect 22554 25480 22560 25492
rect 21959 25452 22560 25480
rect 21959 25449 21971 25452
rect 21913 25443 21971 25449
rect 22554 25440 22560 25452
rect 22612 25440 22618 25492
rect 29733 25483 29791 25489
rect 29733 25449 29745 25483
rect 29779 25480 29791 25483
rect 30098 25480 30104 25492
rect 29779 25452 30104 25480
rect 29779 25449 29791 25452
rect 29733 25443 29791 25449
rect 30098 25440 30104 25452
rect 30156 25440 30162 25492
rect 17681 25415 17739 25421
rect 17681 25381 17693 25415
rect 17727 25412 17739 25415
rect 25866 25412 25872 25424
rect 17727 25384 25872 25412
rect 17727 25381 17739 25384
rect 17681 25375 17739 25381
rect 16574 25304 16580 25356
rect 16632 25344 16638 25356
rect 17696 25344 17724 25375
rect 25866 25372 25872 25384
rect 25924 25372 25930 25424
rect 27157 25415 27215 25421
rect 27157 25381 27169 25415
rect 27203 25412 27215 25415
rect 27203 25384 31754 25412
rect 27203 25381 27215 25384
rect 27157 25375 27215 25381
rect 16632 25316 17724 25344
rect 16632 25304 16638 25316
rect 20070 25304 20076 25356
rect 20128 25344 20134 25356
rect 21269 25347 21327 25353
rect 21269 25344 21281 25347
rect 20128 25316 21281 25344
rect 20128 25304 20134 25316
rect 21269 25313 21281 25316
rect 21315 25313 21327 25347
rect 21269 25307 21327 25313
rect 13202 25248 15332 25276
rect 15378 25236 15384 25288
rect 15436 25276 15442 25288
rect 15746 25276 15752 25288
rect 15436 25248 15752 25276
rect 15436 25236 15442 25248
rect 15746 25236 15752 25248
rect 15804 25276 15810 25288
rect 15933 25279 15991 25285
rect 15933 25276 15945 25279
rect 15804 25248 15945 25276
rect 15804 25236 15810 25248
rect 15933 25245 15945 25248
rect 15979 25245 15991 25279
rect 15933 25239 15991 25245
rect 18693 25279 18751 25285
rect 18693 25245 18705 25279
rect 18739 25276 18751 25279
rect 18782 25276 18788 25288
rect 18739 25248 18788 25276
rect 18739 25245 18751 25248
rect 18693 25239 18751 25245
rect 18782 25236 18788 25248
rect 18840 25236 18846 25288
rect 19334 25236 19340 25288
rect 19392 25276 19398 25288
rect 19429 25279 19487 25285
rect 19429 25276 19441 25279
rect 19392 25248 19441 25276
rect 19392 25236 19398 25248
rect 19429 25245 19441 25248
rect 19475 25245 19487 25279
rect 19978 25276 19984 25288
rect 19429 25239 19487 25245
rect 19536 25248 19984 25276
rect 16209 25211 16267 25217
rect 16209 25177 16221 25211
rect 16255 25177 16267 25211
rect 19536 25208 19564 25248
rect 19978 25236 19984 25248
rect 20036 25236 20042 25288
rect 20438 25236 20444 25288
rect 20496 25276 20502 25288
rect 20622 25276 20628 25288
rect 20496 25248 20628 25276
rect 20496 25236 20502 25248
rect 20622 25236 20628 25248
rect 20680 25236 20686 25288
rect 20714 25236 20720 25288
rect 20772 25236 20778 25288
rect 21450 25276 21456 25288
rect 21411 25248 21456 25276
rect 21450 25236 21456 25248
rect 21508 25236 21514 25288
rect 22922 25236 22928 25288
rect 22980 25276 22986 25288
rect 23750 25276 23756 25288
rect 22980 25248 23756 25276
rect 22980 25236 22986 25248
rect 23750 25236 23756 25248
rect 23808 25236 23814 25288
rect 27154 25236 27160 25288
rect 27212 25276 27218 25288
rect 27341 25279 27399 25285
rect 27341 25276 27353 25279
rect 27212 25248 27353 25276
rect 27212 25236 27218 25248
rect 27341 25245 27353 25248
rect 27387 25245 27399 25279
rect 28534 25276 28540 25288
rect 28495 25248 28540 25276
rect 27341 25239 27399 25245
rect 28534 25236 28540 25248
rect 28592 25236 28598 25288
rect 29178 25276 29184 25288
rect 29139 25248 29184 25276
rect 29178 25236 29184 25248
rect 29236 25236 29242 25288
rect 29917 25279 29975 25285
rect 29917 25245 29929 25279
rect 29963 25245 29975 25279
rect 29917 25239 29975 25245
rect 17434 25180 19564 25208
rect 19705 25211 19763 25217
rect 16209 25171 16267 25177
rect 19705 25177 19717 25211
rect 19751 25208 19763 25211
rect 20732 25208 20760 25236
rect 29932 25208 29960 25239
rect 19751 25180 20760 25208
rect 29012 25180 29960 25208
rect 31726 25208 31754 25384
rect 36170 25208 36176 25220
rect 31726 25180 36176 25208
rect 19751 25177 19763 25180
rect 19705 25171 19763 25177
rect 9674 25140 9680 25152
rect 8956 25112 9680 25140
rect 9674 25100 9680 25112
rect 9732 25100 9738 25152
rect 13541 25143 13599 25149
rect 13541 25109 13553 25143
rect 13587 25140 13599 25143
rect 15746 25140 15752 25152
rect 13587 25112 15752 25140
rect 13587 25109 13599 25112
rect 13541 25103 13599 25109
rect 15746 25100 15752 25112
rect 15804 25100 15810 25152
rect 16224 25140 16252 25171
rect 18598 25140 18604 25152
rect 16224 25112 18604 25140
rect 18598 25100 18604 25112
rect 18656 25100 18662 25152
rect 18785 25143 18843 25149
rect 18785 25109 18797 25143
rect 18831 25140 18843 25143
rect 18874 25140 18880 25152
rect 18831 25112 18880 25140
rect 18831 25109 18843 25112
rect 18785 25103 18843 25109
rect 18874 25100 18880 25112
rect 18932 25100 18938 25152
rect 20714 25140 20720 25152
rect 20675 25112 20720 25140
rect 20714 25100 20720 25112
rect 20772 25100 20778 25152
rect 28353 25143 28411 25149
rect 28353 25109 28365 25143
rect 28399 25140 28411 25143
rect 28626 25140 28632 25152
rect 28399 25112 28632 25140
rect 28399 25109 28411 25112
rect 28353 25103 28411 25109
rect 28626 25100 28632 25112
rect 28684 25100 28690 25152
rect 29012 25149 29040 25180
rect 36170 25168 36176 25180
rect 36228 25168 36234 25220
rect 28997 25143 29055 25149
rect 28997 25109 29009 25143
rect 29043 25109 29055 25143
rect 28997 25103 29055 25109
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 14108 24908 15700 24936
rect 1762 24800 1768 24812
rect 1723 24772 1768 24800
rect 1762 24760 1768 24772
rect 1820 24760 1826 24812
rect 4709 24803 4767 24809
rect 4709 24769 4721 24803
rect 4755 24800 4767 24803
rect 6914 24800 6920 24812
rect 4755 24772 6920 24800
rect 4755 24769 4767 24772
rect 4709 24763 4767 24769
rect 6914 24760 6920 24772
rect 6972 24760 6978 24812
rect 8386 24800 8392 24812
rect 8347 24772 8392 24800
rect 8386 24760 8392 24772
rect 8444 24760 8450 24812
rect 9766 24760 9772 24812
rect 9824 24760 9830 24812
rect 11701 24803 11759 24809
rect 11701 24798 11713 24803
rect 11624 24770 11713 24798
rect 4614 24692 4620 24744
rect 4672 24732 4678 24744
rect 5445 24735 5503 24741
rect 5445 24732 5457 24735
rect 4672 24704 5457 24732
rect 4672 24692 4678 24704
rect 5445 24701 5457 24704
rect 5491 24701 5503 24735
rect 5445 24695 5503 24701
rect 5994 24692 6000 24744
rect 6052 24732 6058 24744
rect 8665 24735 8723 24741
rect 8665 24732 8677 24735
rect 6052 24704 8677 24732
rect 6052 24692 6058 24704
rect 8665 24701 8677 24704
rect 8711 24701 8723 24735
rect 11330 24732 11336 24744
rect 8665 24695 8723 24701
rect 10060 24704 11336 24732
rect 1210 24556 1216 24608
rect 1268 24596 1274 24608
rect 1581 24599 1639 24605
rect 1581 24596 1593 24599
rect 1268 24568 1593 24596
rect 1268 24556 1274 24568
rect 1581 24565 1593 24568
rect 1627 24565 1639 24599
rect 1581 24559 1639 24565
rect 4062 24556 4068 24608
rect 4120 24596 4126 24608
rect 4706 24596 4712 24608
rect 4120 24568 4712 24596
rect 4120 24556 4126 24568
rect 4706 24556 4712 24568
rect 4764 24556 4770 24608
rect 6914 24556 6920 24608
rect 6972 24596 6978 24608
rect 7926 24596 7932 24608
rect 6972 24568 7932 24596
rect 6972 24556 6978 24568
rect 7926 24556 7932 24568
rect 7984 24596 7990 24608
rect 10060 24596 10088 24704
rect 11330 24692 11336 24704
rect 11388 24732 11394 24744
rect 11624 24732 11652 24770
rect 11701 24769 11713 24770
rect 11747 24769 11759 24803
rect 11701 24763 11759 24769
rect 13081 24803 13139 24809
rect 13081 24769 13093 24803
rect 13127 24769 13139 24803
rect 13081 24763 13139 24769
rect 11388 24704 11652 24732
rect 11388 24692 11394 24704
rect 11790 24692 11796 24744
rect 11848 24732 11854 24744
rect 12437 24735 12495 24741
rect 12437 24732 12449 24735
rect 11848 24704 12449 24732
rect 11848 24692 11854 24704
rect 12437 24701 12449 24704
rect 12483 24701 12495 24735
rect 12437 24695 12495 24701
rect 13096 24732 13124 24763
rect 13170 24760 13176 24812
rect 13228 24800 13234 24812
rect 14108 24800 14136 24908
rect 13228 24772 13273 24800
rect 13372 24772 14136 24800
rect 13228 24760 13234 24772
rect 13372 24732 13400 24772
rect 15470 24760 15476 24812
rect 15528 24760 15534 24812
rect 15672 24800 15700 24908
rect 15746 24896 15752 24948
rect 15804 24936 15810 24948
rect 29178 24936 29184 24948
rect 15804 24908 29184 24936
rect 15804 24896 15810 24908
rect 29178 24896 29184 24908
rect 29236 24896 29242 24948
rect 16758 24828 16764 24880
rect 16816 24828 16822 24880
rect 17037 24871 17095 24877
rect 17037 24837 17049 24871
rect 17083 24868 17095 24871
rect 17083 24840 17816 24868
rect 17083 24837 17095 24840
rect 17037 24831 17095 24837
rect 16776 24800 16804 24828
rect 15672 24772 16804 24800
rect 17788 24800 17816 24840
rect 18966 24828 18972 24880
rect 19024 24868 19030 24880
rect 22925 24871 22983 24877
rect 19024 24840 20208 24868
rect 19024 24828 19030 24840
rect 20180 24812 20208 24840
rect 22925 24837 22937 24871
rect 22971 24868 22983 24871
rect 27522 24868 27528 24880
rect 22971 24840 23520 24868
rect 27483 24840 27528 24868
rect 22971 24837 22983 24840
rect 22925 24831 22983 24837
rect 18785 24803 18843 24809
rect 17788 24772 18092 24800
rect 13096 24704 13400 24732
rect 14093 24735 14151 24741
rect 10134 24624 10140 24676
rect 10192 24664 10198 24676
rect 12986 24664 12992 24676
rect 10192 24636 12992 24664
rect 10192 24624 10198 24636
rect 12986 24624 12992 24636
rect 13044 24624 13050 24676
rect 7984 24568 10088 24596
rect 7984 24556 7990 24568
rect 10594 24556 10600 24608
rect 10652 24596 10658 24608
rect 13096 24596 13124 24704
rect 14093 24701 14105 24735
rect 14139 24701 14151 24735
rect 14093 24695 14151 24701
rect 14369 24735 14427 24741
rect 14369 24701 14381 24735
rect 14415 24732 14427 24735
rect 16945 24735 17003 24741
rect 14415 24704 15516 24732
rect 14415 24701 14427 24704
rect 14369 24695 14427 24701
rect 10652 24568 13124 24596
rect 14108 24596 14136 24695
rect 15488 24664 15516 24704
rect 16945 24701 16957 24735
rect 16991 24732 17003 24735
rect 17218 24732 17224 24744
rect 16991 24704 17080 24732
rect 17179 24704 17224 24732
rect 16991 24701 17003 24704
rect 16945 24695 17003 24701
rect 16758 24664 16764 24676
rect 15488 24636 16764 24664
rect 16758 24624 16764 24636
rect 16816 24624 16822 24676
rect 17052 24664 17080 24704
rect 17218 24692 17224 24704
rect 17276 24732 17282 24744
rect 17586 24732 17592 24744
rect 17276 24704 17592 24732
rect 17276 24692 17282 24704
rect 17586 24692 17592 24704
rect 17644 24692 17650 24744
rect 18064 24732 18092 24772
rect 18785 24769 18797 24803
rect 18831 24800 18843 24803
rect 18874 24800 18880 24812
rect 18831 24772 18880 24800
rect 18831 24769 18843 24772
rect 18785 24763 18843 24769
rect 18874 24760 18880 24772
rect 18932 24760 18938 24812
rect 19061 24803 19119 24809
rect 19061 24769 19073 24803
rect 19107 24800 19119 24803
rect 19978 24800 19984 24812
rect 19107 24772 19984 24800
rect 19107 24769 19119 24772
rect 19061 24763 19119 24769
rect 19978 24760 19984 24772
rect 20036 24760 20042 24812
rect 20162 24760 20168 24812
rect 20220 24800 20226 24812
rect 20257 24803 20315 24809
rect 20257 24800 20269 24803
rect 20220 24772 20269 24800
rect 20220 24760 20226 24772
rect 20257 24769 20269 24772
rect 20303 24769 20315 24803
rect 20257 24763 20315 24769
rect 20622 24760 20628 24812
rect 20680 24800 20686 24812
rect 20893 24803 20951 24809
rect 20893 24800 20905 24803
rect 20680 24772 20905 24800
rect 20680 24760 20686 24772
rect 20893 24769 20905 24772
rect 20939 24769 20951 24803
rect 20893 24763 20951 24769
rect 20990 24760 20996 24812
rect 21048 24800 21054 24812
rect 21048 24772 21093 24800
rect 21048 24760 21054 24772
rect 20806 24732 20812 24744
rect 18064 24704 20812 24732
rect 20806 24692 20812 24704
rect 20864 24692 20870 24744
rect 21910 24692 21916 24744
rect 21968 24732 21974 24744
rect 22833 24735 22891 24741
rect 22833 24732 22845 24735
rect 21968 24704 22845 24732
rect 21968 24692 21974 24704
rect 22833 24701 22845 24704
rect 22879 24732 22891 24735
rect 23492 24732 23520 24840
rect 27522 24828 27528 24840
rect 27580 24828 27586 24880
rect 23934 24800 23940 24812
rect 23895 24772 23940 24800
rect 23934 24760 23940 24772
rect 23992 24760 23998 24812
rect 25406 24760 25412 24812
rect 25464 24800 25470 24812
rect 25593 24803 25651 24809
rect 25593 24800 25605 24803
rect 25464 24772 25605 24800
rect 25464 24760 25470 24772
rect 25593 24769 25605 24772
rect 25639 24800 25651 24803
rect 27154 24800 27160 24812
rect 25639 24772 27160 24800
rect 25639 24769 25651 24772
rect 25593 24763 25651 24769
rect 27154 24760 27160 24772
rect 27212 24760 27218 24812
rect 29086 24760 29092 24812
rect 29144 24800 29150 24812
rect 38013 24803 38071 24809
rect 38013 24800 38025 24803
rect 29144 24772 38025 24800
rect 29144 24760 29150 24772
rect 38013 24769 38025 24772
rect 38059 24769 38071 24803
rect 38013 24763 38071 24769
rect 24029 24735 24087 24741
rect 24029 24732 24041 24735
rect 22879 24704 23060 24732
rect 23492 24704 24041 24732
rect 22879 24701 22891 24704
rect 22833 24695 22891 24701
rect 17126 24664 17132 24676
rect 17052 24636 17132 24664
rect 17126 24624 17132 24636
rect 17184 24624 17190 24676
rect 17402 24624 17408 24676
rect 17460 24664 17466 24676
rect 21358 24664 21364 24676
rect 17460 24636 21364 24664
rect 17460 24624 17466 24636
rect 21358 24624 21364 24636
rect 21416 24624 21422 24676
rect 21634 24624 21640 24676
rect 21692 24664 21698 24676
rect 22922 24664 22928 24676
rect 21692 24636 22928 24664
rect 21692 24624 21698 24636
rect 22922 24624 22928 24636
rect 22980 24624 22986 24676
rect 15378 24596 15384 24608
rect 14108 24568 15384 24596
rect 10652 24556 10658 24568
rect 15378 24556 15384 24568
rect 15436 24556 15442 24608
rect 15841 24599 15899 24605
rect 15841 24565 15853 24599
rect 15887 24596 15899 24599
rect 15930 24596 15936 24608
rect 15887 24568 15936 24596
rect 15887 24565 15899 24568
rect 15841 24559 15899 24565
rect 15930 24556 15936 24568
rect 15988 24556 15994 24608
rect 18230 24556 18236 24608
rect 18288 24596 18294 24608
rect 20349 24599 20407 24605
rect 20349 24596 20361 24599
rect 18288 24568 20361 24596
rect 18288 24556 18294 24568
rect 20349 24565 20361 24568
rect 20395 24565 20407 24599
rect 20349 24559 20407 24565
rect 20530 24556 20536 24608
rect 20588 24596 20594 24608
rect 22002 24596 22008 24608
rect 20588 24568 22008 24596
rect 20588 24556 20594 24568
rect 22002 24556 22008 24568
rect 22060 24556 22066 24608
rect 23032 24596 23060 24704
rect 24029 24701 24041 24704
rect 24075 24701 24087 24735
rect 24029 24695 24087 24701
rect 27246 24692 27252 24744
rect 27304 24732 27310 24744
rect 27433 24735 27491 24741
rect 27433 24732 27445 24735
rect 27304 24704 27445 24732
rect 27304 24692 27310 24704
rect 27433 24701 27445 24704
rect 27479 24701 27491 24735
rect 28350 24732 28356 24744
rect 28311 24704 28356 24732
rect 27433 24695 27491 24701
rect 28350 24692 28356 24704
rect 28408 24692 28414 24744
rect 28534 24692 28540 24744
rect 28592 24732 28598 24744
rect 28997 24735 29055 24741
rect 28997 24732 29009 24735
rect 28592 24704 29009 24732
rect 28592 24692 28598 24704
rect 28997 24701 29009 24704
rect 29043 24701 29055 24735
rect 28997 24695 29055 24701
rect 23385 24667 23443 24673
rect 23385 24633 23397 24667
rect 23431 24664 23443 24667
rect 23842 24664 23848 24676
rect 23431 24636 23848 24664
rect 23431 24633 23443 24636
rect 23385 24627 23443 24633
rect 23842 24624 23848 24636
rect 23900 24624 23906 24676
rect 24210 24596 24216 24608
rect 23032 24568 24216 24596
rect 24210 24556 24216 24568
rect 24268 24556 24274 24608
rect 25590 24556 25596 24608
rect 25648 24596 25654 24608
rect 25685 24599 25743 24605
rect 25685 24596 25697 24599
rect 25648 24568 25697 24596
rect 25648 24556 25654 24568
rect 25685 24565 25697 24568
rect 25731 24565 25743 24599
rect 38194 24596 38200 24608
rect 38155 24568 38200 24596
rect 25685 24559 25743 24565
rect 38194 24556 38200 24568
rect 38252 24556 38258 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 2682 24352 2688 24404
rect 2740 24392 2746 24404
rect 2740 24364 6408 24392
rect 2740 24352 2746 24364
rect 6380 24324 6408 24364
rect 6454 24352 6460 24404
rect 6512 24392 6518 24404
rect 9582 24392 9588 24404
rect 6512 24364 9588 24392
rect 6512 24352 6518 24364
rect 9582 24352 9588 24364
rect 9640 24352 9646 24404
rect 9766 24352 9772 24404
rect 9824 24392 9830 24404
rect 13906 24392 13912 24404
rect 9824 24364 13912 24392
rect 9824 24352 9830 24364
rect 13906 24352 13912 24364
rect 13964 24352 13970 24404
rect 21726 24392 21732 24404
rect 14016 24364 21732 24392
rect 6380 24296 6592 24324
rect 1673 24259 1731 24265
rect 1673 24225 1685 24259
rect 1719 24256 1731 24259
rect 3973 24259 4031 24265
rect 3973 24256 3985 24259
rect 1719 24228 3985 24256
rect 1719 24225 1731 24228
rect 1673 24219 1731 24225
rect 3973 24225 3985 24228
rect 4019 24256 4031 24259
rect 4246 24256 4252 24268
rect 4019 24228 4252 24256
rect 4019 24225 4031 24228
rect 3973 24219 4031 24225
rect 4246 24216 4252 24228
rect 4304 24256 4310 24268
rect 4614 24256 4620 24268
rect 4304 24228 4620 24256
rect 4304 24216 4310 24228
rect 4614 24216 4620 24228
rect 4672 24256 4678 24268
rect 6564 24256 6592 24296
rect 7742 24284 7748 24336
rect 7800 24324 7806 24336
rect 11698 24324 11704 24336
rect 7800 24296 11704 24324
rect 7800 24284 7806 24296
rect 11698 24284 11704 24296
rect 11756 24284 11762 24336
rect 12986 24284 12992 24336
rect 13044 24324 13050 24336
rect 14016 24324 14044 24364
rect 21726 24352 21732 24364
rect 21784 24352 21790 24404
rect 25406 24392 25412 24404
rect 21928 24364 25412 24392
rect 21928 24324 21956 24364
rect 25406 24352 25412 24364
rect 25464 24352 25470 24404
rect 29638 24392 29644 24404
rect 27908 24364 29644 24392
rect 13044 24296 14044 24324
rect 17236 24296 21956 24324
rect 13044 24284 13050 24296
rect 17236 24256 17264 24296
rect 22002 24284 22008 24336
rect 22060 24324 22066 24336
rect 22646 24324 22652 24336
rect 22060 24296 22652 24324
rect 22060 24284 22066 24296
rect 22646 24284 22652 24296
rect 22704 24284 22710 24336
rect 27908 24324 27936 24364
rect 29638 24352 29644 24364
rect 29696 24352 29702 24404
rect 29730 24324 29736 24336
rect 24596 24296 27936 24324
rect 28000 24296 29736 24324
rect 4672 24228 6408 24256
rect 6564 24228 17264 24256
rect 4672 24216 4678 24228
rect 5997 24191 6055 24197
rect 5997 24157 6009 24191
rect 6043 24188 6055 24191
rect 6270 24188 6276 24200
rect 6043 24160 6276 24188
rect 6043 24157 6055 24160
rect 5997 24151 6055 24157
rect 6270 24148 6276 24160
rect 6328 24148 6334 24200
rect 6380 24188 6408 24228
rect 18874 24216 18880 24268
rect 18932 24256 18938 24268
rect 19334 24256 19340 24268
rect 18932 24228 19340 24256
rect 18932 24216 18938 24228
rect 19334 24216 19340 24228
rect 19392 24216 19398 24268
rect 19426 24216 19432 24268
rect 19484 24216 19490 24268
rect 20257 24259 20315 24265
rect 20257 24225 20269 24259
rect 20303 24256 20315 24259
rect 20303 24228 22692 24256
rect 20303 24225 20315 24228
rect 20257 24219 20315 24225
rect 6457 24191 6515 24197
rect 6457 24188 6469 24191
rect 6380 24160 6469 24188
rect 6457 24157 6469 24160
rect 6503 24157 6515 24191
rect 15378 24188 15384 24200
rect 15339 24160 15384 24188
rect 6457 24151 6515 24157
rect 15378 24148 15384 24160
rect 15436 24148 15442 24200
rect 19444 24188 19472 24216
rect 16790 24160 19472 24188
rect 21085 24191 21143 24197
rect 21085 24157 21097 24191
rect 21131 24188 21143 24191
rect 21542 24188 21548 24200
rect 21131 24160 21548 24188
rect 21131 24157 21143 24160
rect 21085 24151 21143 24157
rect 21542 24148 21548 24160
rect 21600 24148 21606 24200
rect 22664 24188 22692 24228
rect 22830 24216 22836 24268
rect 22888 24256 22894 24268
rect 23198 24256 23204 24268
rect 22888 24228 23204 24256
rect 22888 24216 22894 24228
rect 23198 24216 23204 24228
rect 23256 24216 23262 24268
rect 24596 24197 24624 24296
rect 28000 24197 28028 24296
rect 29730 24284 29736 24296
rect 29788 24284 29794 24336
rect 28534 24256 28540 24268
rect 28495 24228 28540 24256
rect 28534 24216 28540 24228
rect 28592 24216 28598 24268
rect 29181 24259 29239 24265
rect 29181 24225 29193 24259
rect 29227 24256 29239 24259
rect 29914 24256 29920 24268
rect 29227 24228 29920 24256
rect 29227 24225 29239 24228
rect 29181 24219 29239 24225
rect 29914 24216 29920 24228
rect 29972 24216 29978 24268
rect 24581 24191 24639 24197
rect 22664 24160 24532 24188
rect 1118 24080 1124 24132
rect 1176 24120 1182 24132
rect 1946 24120 1952 24132
rect 1176 24092 1952 24120
rect 1176 24080 1182 24092
rect 1946 24080 1952 24092
rect 2004 24080 2010 24132
rect 2498 24080 2504 24132
rect 2556 24080 2562 24132
rect 4249 24123 4307 24129
rect 4249 24089 4261 24123
rect 4295 24120 4307 24123
rect 4522 24120 4528 24132
rect 4295 24092 4528 24120
rect 4295 24089 4307 24092
rect 4249 24083 4307 24089
rect 4522 24080 4528 24092
rect 4580 24080 4586 24132
rect 4798 24080 4804 24132
rect 4856 24080 4862 24132
rect 6362 24080 6368 24132
rect 6420 24120 6426 24132
rect 6733 24123 6791 24129
rect 6733 24120 6745 24123
rect 6420 24092 6745 24120
rect 6420 24080 6426 24092
rect 6733 24089 6745 24092
rect 6779 24089 6791 24123
rect 9214 24120 9220 24132
rect 7958 24092 9220 24120
rect 6733 24083 6791 24089
rect 9214 24080 9220 24092
rect 9272 24080 9278 24132
rect 15657 24123 15715 24129
rect 15657 24089 15669 24123
rect 15703 24089 15715 24123
rect 15657 24083 15715 24089
rect 2038 24012 2044 24064
rect 2096 24052 2102 24064
rect 3421 24055 3479 24061
rect 3421 24052 3433 24055
rect 2096 24024 3433 24052
rect 2096 24012 2102 24024
rect 3421 24021 3433 24024
rect 3467 24021 3479 24055
rect 8202 24052 8208 24064
rect 8163 24024 8208 24052
rect 3421 24015 3479 24021
rect 8202 24012 8208 24024
rect 8260 24012 8266 24064
rect 9582 24012 9588 24064
rect 9640 24052 9646 24064
rect 10778 24052 10784 24064
rect 9640 24024 10784 24052
rect 9640 24012 9646 24024
rect 10778 24012 10784 24024
rect 10836 24052 10842 24064
rect 13722 24052 13728 24064
rect 10836 24024 13728 24052
rect 10836 24012 10842 24024
rect 13722 24012 13728 24024
rect 13780 24012 13786 24064
rect 15672 24052 15700 24083
rect 19426 24080 19432 24132
rect 19484 24120 19490 24132
rect 19613 24123 19671 24129
rect 19613 24120 19625 24123
rect 19484 24092 19625 24120
rect 19484 24080 19490 24092
rect 19613 24089 19625 24092
rect 19659 24089 19671 24123
rect 19613 24083 19671 24089
rect 19705 24123 19763 24129
rect 19705 24089 19717 24123
rect 19751 24120 19763 24123
rect 20622 24120 20628 24132
rect 19751 24092 20628 24120
rect 19751 24089 19763 24092
rect 19705 24083 19763 24089
rect 20622 24080 20628 24092
rect 20680 24080 20686 24132
rect 21821 24123 21879 24129
rect 21821 24120 21833 24123
rect 21744 24092 21833 24120
rect 21744 24064 21772 24092
rect 21821 24089 21833 24092
rect 21867 24089 21879 24123
rect 21821 24083 21879 24089
rect 21913 24123 21971 24129
rect 21913 24089 21925 24123
rect 21959 24089 21971 24123
rect 24504 24120 24532 24160
rect 24581 24157 24593 24191
rect 24627 24157 24639 24191
rect 24581 24151 24639 24157
rect 27985 24191 28043 24197
rect 27985 24157 27997 24191
rect 28031 24157 28043 24191
rect 27985 24151 28043 24157
rect 34698 24148 34704 24200
rect 34756 24188 34762 24200
rect 38013 24191 38071 24197
rect 38013 24188 38025 24191
rect 34756 24160 38025 24188
rect 34756 24148 34762 24160
rect 38013 24157 38025 24160
rect 38059 24157 38071 24191
rect 38013 24151 38071 24157
rect 27706 24120 27712 24132
rect 24504 24092 27712 24120
rect 21913 24083 21971 24089
rect 16574 24052 16580 24064
rect 15672 24024 16580 24052
rect 16574 24012 16580 24024
rect 16632 24012 16638 24064
rect 17126 24052 17132 24064
rect 17087 24024 17132 24052
rect 17126 24012 17132 24024
rect 17184 24012 17190 24064
rect 18138 24012 18144 24064
rect 18196 24052 18202 24064
rect 18233 24055 18291 24061
rect 18233 24052 18245 24055
rect 18196 24024 18245 24052
rect 18196 24012 18202 24024
rect 18233 24021 18245 24024
rect 18279 24021 18291 24055
rect 18233 24015 18291 24021
rect 19978 24012 19984 24064
rect 20036 24052 20042 24064
rect 21177 24055 21235 24061
rect 21177 24052 21189 24055
rect 20036 24024 21189 24052
rect 20036 24012 20042 24024
rect 21177 24021 21189 24024
rect 21223 24021 21235 24055
rect 21177 24015 21235 24021
rect 21726 24012 21732 24064
rect 21784 24012 21790 24064
rect 21928 24052 21956 24083
rect 27706 24080 27712 24092
rect 27764 24080 27770 24132
rect 28626 24120 28632 24132
rect 28587 24092 28632 24120
rect 28626 24080 28632 24092
rect 28684 24080 28690 24132
rect 24673 24055 24731 24061
rect 24673 24052 24685 24055
rect 21928 24024 24685 24052
rect 24673 24021 24685 24024
rect 24719 24021 24731 24055
rect 24673 24015 24731 24021
rect 27801 24055 27859 24061
rect 27801 24021 27813 24055
rect 27847 24052 27859 24055
rect 28902 24052 28908 24064
rect 27847 24024 28908 24052
rect 27847 24021 27859 24024
rect 27801 24015 27859 24021
rect 28902 24012 28908 24024
rect 28960 24012 28966 24064
rect 38194 24052 38200 24064
rect 38155 24024 38200 24052
rect 38194 24012 38200 24024
rect 38252 24012 38258 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 4706 23808 4712 23860
rect 4764 23848 4770 23860
rect 5166 23848 5172 23860
rect 4764 23820 5172 23848
rect 4764 23808 4770 23820
rect 5166 23808 5172 23820
rect 5224 23808 5230 23860
rect 11790 23848 11796 23860
rect 7944 23820 11796 23848
rect 4154 23780 4160 23792
rect 1964 23752 4160 23780
rect 1964 23721 1992 23752
rect 4154 23740 4160 23752
rect 4212 23740 4218 23792
rect 4525 23783 4583 23789
rect 4525 23749 4537 23783
rect 4571 23780 4583 23783
rect 4724 23780 4752 23808
rect 7742 23780 7748 23792
rect 4571 23752 4752 23780
rect 5750 23752 7748 23780
rect 4571 23749 4583 23752
rect 4525 23743 4583 23749
rect 7742 23740 7748 23752
rect 7800 23740 7806 23792
rect 1949 23715 2007 23721
rect 1949 23681 1961 23715
rect 1995 23681 2007 23715
rect 1949 23675 2007 23681
rect 2593 23715 2651 23721
rect 2593 23681 2605 23715
rect 2639 23712 2651 23715
rect 2774 23712 2780 23724
rect 2639 23684 2780 23712
rect 2639 23681 2651 23684
rect 2593 23675 2651 23681
rect 2774 23672 2780 23684
rect 2832 23672 2838 23724
rect 4246 23712 4252 23724
rect 4207 23684 4252 23712
rect 4246 23672 4252 23684
rect 4304 23672 4310 23724
rect 7944 23721 7972 23820
rect 11790 23808 11796 23820
rect 11848 23808 11854 23860
rect 16482 23808 16488 23860
rect 16540 23848 16546 23860
rect 16945 23851 17003 23857
rect 16945 23848 16957 23851
rect 16540 23820 16957 23848
rect 16540 23808 16546 23820
rect 16945 23817 16957 23820
rect 16991 23817 17003 23851
rect 23661 23851 23719 23857
rect 23661 23848 23673 23851
rect 16945 23811 17003 23817
rect 18340 23820 23673 23848
rect 8662 23740 8668 23792
rect 8720 23740 8726 23792
rect 11330 23740 11336 23792
rect 11388 23780 11394 23792
rect 15381 23783 15439 23789
rect 15381 23780 15393 23783
rect 11388 23752 15393 23780
rect 11388 23740 11394 23752
rect 15381 23749 15393 23752
rect 15427 23749 15439 23783
rect 18138 23780 18144 23792
rect 15381 23743 15439 23749
rect 16684 23752 17448 23780
rect 18099 23752 18144 23780
rect 7929 23715 7987 23721
rect 7929 23681 7941 23715
rect 7975 23681 7987 23715
rect 7929 23675 7987 23681
rect 13722 23672 13728 23724
rect 13780 23712 13786 23724
rect 16684 23712 16712 23752
rect 16850 23712 16856 23724
rect 13780 23684 16712 23712
rect 16811 23684 16856 23712
rect 13780 23672 13786 23684
rect 16850 23672 16856 23684
rect 16908 23672 16914 23724
rect 2866 23604 2872 23656
rect 2924 23644 2930 23656
rect 8205 23647 8263 23653
rect 2924 23616 6914 23644
rect 2924 23604 2930 23616
rect 1486 23468 1492 23520
rect 1544 23508 1550 23520
rect 1765 23511 1823 23517
rect 1765 23508 1777 23511
rect 1544 23480 1777 23508
rect 1544 23468 1550 23480
rect 1765 23477 1777 23480
rect 1811 23477 1823 23511
rect 1765 23471 1823 23477
rect 2409 23511 2467 23517
rect 2409 23477 2421 23511
rect 2455 23508 2467 23511
rect 2682 23508 2688 23520
rect 2455 23480 2688 23508
rect 2455 23477 2467 23480
rect 2409 23471 2467 23477
rect 2682 23468 2688 23480
rect 2740 23468 2746 23520
rect 5997 23511 6055 23517
rect 5997 23477 6009 23511
rect 6043 23508 6055 23511
rect 6362 23508 6368 23520
rect 6043 23480 6368 23508
rect 6043 23477 6055 23480
rect 5997 23471 6055 23477
rect 6362 23468 6368 23480
rect 6420 23468 6426 23520
rect 6886 23508 6914 23616
rect 8205 23613 8217 23647
rect 8251 23644 8263 23647
rect 10134 23644 10140 23656
rect 8251 23616 10140 23644
rect 8251 23613 8263 23616
rect 8205 23607 8263 23613
rect 10134 23604 10140 23616
rect 10192 23604 10198 23656
rect 15378 23604 15384 23656
rect 15436 23644 15442 23656
rect 16117 23647 16175 23653
rect 16117 23644 16129 23647
rect 15436 23616 16129 23644
rect 15436 23604 15442 23616
rect 16117 23613 16129 23616
rect 16163 23613 16175 23647
rect 17420 23644 17448 23752
rect 18138 23740 18144 23752
rect 18196 23740 18202 23792
rect 18242 23783 18300 23789
rect 18242 23749 18254 23783
rect 18288 23780 18300 23783
rect 18340 23780 18368 23820
rect 23661 23817 23673 23820
rect 23707 23817 23719 23851
rect 23661 23811 23719 23817
rect 24026 23808 24032 23860
rect 24084 23848 24090 23860
rect 29086 23848 29092 23860
rect 24084 23820 25728 23848
rect 24084 23808 24090 23820
rect 18288 23752 18368 23780
rect 18785 23783 18843 23789
rect 18288 23749 18300 23752
rect 18242 23743 18300 23749
rect 18785 23749 18797 23783
rect 18831 23780 18843 23783
rect 20162 23780 20168 23792
rect 18831 23752 20168 23780
rect 18831 23749 18843 23752
rect 18785 23743 18843 23749
rect 20162 23740 20168 23752
rect 20220 23740 20226 23792
rect 20625 23783 20683 23789
rect 20625 23749 20637 23783
rect 20671 23780 20683 23783
rect 21450 23780 21456 23792
rect 20671 23752 21456 23780
rect 20671 23749 20683 23752
rect 20625 23743 20683 23749
rect 21450 23740 21456 23752
rect 21508 23740 21514 23792
rect 23014 23740 23020 23792
rect 23072 23780 23078 23792
rect 24305 23783 24363 23789
rect 24305 23780 24317 23783
rect 23072 23752 24317 23780
rect 23072 23740 23078 23752
rect 24305 23749 24317 23752
rect 24351 23749 24363 23783
rect 25590 23780 25596 23792
rect 25551 23752 25596 23780
rect 24305 23743 24363 23749
rect 25590 23740 25596 23752
rect 25648 23740 25654 23792
rect 25700 23789 25728 23820
rect 27724 23820 29092 23848
rect 27724 23789 27752 23820
rect 29086 23808 29092 23820
rect 29144 23808 29150 23860
rect 25685 23783 25743 23789
rect 25685 23749 25697 23783
rect 25731 23749 25743 23783
rect 25685 23743 25743 23749
rect 27709 23783 27767 23789
rect 27709 23749 27721 23783
rect 27755 23749 27767 23783
rect 27709 23743 27767 23749
rect 27801 23783 27859 23789
rect 27801 23749 27813 23783
rect 27847 23780 27859 23783
rect 27890 23780 27896 23792
rect 27847 23752 27896 23780
rect 27847 23749 27859 23752
rect 27801 23743 27859 23749
rect 27890 23740 27896 23752
rect 27948 23740 27954 23792
rect 19150 23672 19156 23724
rect 19208 23712 19214 23724
rect 20533 23715 20591 23721
rect 20533 23712 20545 23715
rect 19208 23684 20545 23712
rect 19208 23672 19214 23684
rect 20533 23681 20545 23684
rect 20579 23681 20591 23715
rect 20533 23675 20591 23681
rect 20806 23672 20812 23724
rect 20864 23712 20870 23724
rect 22005 23715 22063 23721
rect 22005 23712 22017 23715
rect 20864 23684 22017 23712
rect 20864 23672 20870 23684
rect 22005 23681 22017 23684
rect 22051 23681 22063 23715
rect 22646 23712 22652 23724
rect 22607 23684 22652 23712
rect 22005 23675 22063 23681
rect 22646 23672 22652 23684
rect 22704 23672 22710 23724
rect 23569 23715 23627 23721
rect 23569 23681 23581 23715
rect 23615 23712 23627 23715
rect 24118 23712 24124 23724
rect 23615 23684 24124 23712
rect 23615 23681 23627 23684
rect 23569 23675 23627 23681
rect 24118 23672 24124 23684
rect 24176 23672 24182 23724
rect 27522 23712 27528 23724
rect 26436 23684 27528 23712
rect 21634 23644 21640 23656
rect 17420 23616 21640 23644
rect 16117 23607 16175 23613
rect 21634 23604 21640 23616
rect 21692 23604 21698 23656
rect 22097 23647 22155 23653
rect 22097 23613 22109 23647
rect 22143 23644 22155 23647
rect 26436 23644 26464 23684
rect 27522 23672 27528 23684
rect 27580 23672 27586 23724
rect 33226 23672 33232 23724
rect 33284 23712 33290 23724
rect 34241 23715 34299 23721
rect 34241 23712 34253 23715
rect 33284 23684 34253 23712
rect 33284 23672 33290 23684
rect 34241 23681 34253 23684
rect 34287 23681 34299 23715
rect 34241 23675 34299 23681
rect 22143 23616 26464 23644
rect 26605 23647 26663 23653
rect 22143 23613 22155 23616
rect 22097 23607 22155 23613
rect 26605 23613 26617 23647
rect 26651 23644 26663 23647
rect 26878 23644 26884 23656
rect 26651 23616 26884 23644
rect 26651 23613 26663 23616
rect 26605 23607 26663 23613
rect 26878 23604 26884 23616
rect 26936 23604 26942 23656
rect 27982 23644 27988 23656
rect 27943 23616 27988 23644
rect 27982 23604 27988 23616
rect 28040 23604 28046 23656
rect 29365 23647 29423 23653
rect 29365 23613 29377 23647
rect 29411 23644 29423 23647
rect 29822 23644 29828 23656
rect 29411 23616 29828 23644
rect 29411 23613 29423 23616
rect 29365 23607 29423 23613
rect 29822 23604 29828 23616
rect 29880 23604 29886 23656
rect 14734 23536 14740 23588
rect 14792 23576 14798 23588
rect 17218 23576 17224 23588
rect 14792 23548 17224 23576
rect 14792 23536 14798 23548
rect 17218 23536 17224 23548
rect 17276 23536 17282 23588
rect 20162 23536 20168 23588
rect 20220 23576 20226 23588
rect 22186 23576 22192 23588
rect 20220 23548 22192 23576
rect 20220 23536 20226 23548
rect 22186 23536 22192 23548
rect 22244 23576 22250 23588
rect 22462 23576 22468 23588
rect 22244 23548 22468 23576
rect 22244 23536 22250 23548
rect 22462 23536 22468 23548
rect 22520 23536 22526 23588
rect 22741 23579 22799 23585
rect 22741 23545 22753 23579
rect 22787 23576 22799 23579
rect 29914 23576 29920 23588
rect 22787 23548 29920 23576
rect 22787 23545 22799 23548
rect 22741 23539 22799 23545
rect 29914 23536 29920 23548
rect 29972 23536 29978 23588
rect 9677 23511 9735 23517
rect 9677 23508 9689 23511
rect 6886 23480 9689 23508
rect 9677 23477 9689 23480
rect 9723 23477 9735 23511
rect 9677 23471 9735 23477
rect 13906 23468 13912 23520
rect 13964 23508 13970 23520
rect 20346 23508 20352 23520
rect 13964 23480 20352 23508
rect 13964 23468 13970 23480
rect 20346 23468 20352 23480
rect 20404 23468 20410 23520
rect 24394 23508 24400 23520
rect 24355 23480 24400 23508
rect 24394 23468 24400 23480
rect 24452 23468 24458 23520
rect 34333 23511 34391 23517
rect 34333 23477 34345 23511
rect 34379 23508 34391 23511
rect 34422 23508 34428 23520
rect 34379 23480 34428 23508
rect 34379 23477 34391 23480
rect 34333 23471 34391 23477
rect 34422 23468 34428 23480
rect 34480 23468 34486 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 15194 23304 15200 23316
rect 10612 23276 15200 23304
rect 4614 23128 4620 23180
rect 4672 23168 4678 23180
rect 5074 23168 5080 23180
rect 4672 23140 5080 23168
rect 4672 23128 4678 23140
rect 5074 23128 5080 23140
rect 5132 23168 5138 23180
rect 5721 23171 5779 23177
rect 5721 23168 5733 23171
rect 5132 23140 5733 23168
rect 5132 23128 5138 23140
rect 5721 23137 5733 23140
rect 5767 23137 5779 23171
rect 5721 23131 5779 23137
rect 5997 23171 6055 23177
rect 5997 23137 6009 23171
rect 6043 23168 6055 23171
rect 10612 23168 10640 23276
rect 15194 23264 15200 23276
rect 15252 23264 15258 23316
rect 20714 23304 20720 23316
rect 15304 23276 20720 23304
rect 12986 23236 12992 23248
rect 11808 23208 12992 23236
rect 6043 23140 10640 23168
rect 10781 23171 10839 23177
rect 6043 23137 6055 23140
rect 5997 23131 6055 23137
rect 10781 23137 10793 23171
rect 10827 23168 10839 23171
rect 11808 23168 11836 23208
rect 12986 23196 12992 23208
rect 13044 23196 13050 23248
rect 15304 23236 15332 23276
rect 20714 23264 20720 23276
rect 20772 23264 20778 23316
rect 28442 23264 28448 23316
rect 28500 23304 28506 23316
rect 28537 23307 28595 23313
rect 28537 23304 28549 23307
rect 28500 23276 28549 23304
rect 28500 23264 28506 23276
rect 28537 23273 28549 23276
rect 28583 23273 28595 23307
rect 28537 23267 28595 23273
rect 14752 23208 15332 23236
rect 14752 23168 14780 23208
rect 16942 23196 16948 23248
rect 17000 23236 17006 23248
rect 20530 23236 20536 23248
rect 17000 23208 20536 23236
rect 17000 23196 17006 23208
rect 20530 23196 20536 23208
rect 20588 23196 20594 23248
rect 10827 23140 11836 23168
rect 11900 23140 14780 23168
rect 10827 23137 10839 23140
rect 10781 23131 10839 23137
rect 1578 23060 1584 23112
rect 1636 23100 1642 23112
rect 1673 23103 1731 23109
rect 1673 23100 1685 23103
rect 1636 23072 1685 23100
rect 1636 23060 1642 23072
rect 1673 23069 1685 23072
rect 1719 23069 1731 23103
rect 1673 23063 1731 23069
rect 9306 23060 9312 23112
rect 9364 23100 9370 23112
rect 10505 23103 10563 23109
rect 10505 23100 10517 23103
rect 9364 23072 10517 23100
rect 9364 23060 9370 23072
rect 10505 23069 10517 23072
rect 10551 23069 10563 23103
rect 11900 23086 11928 23140
rect 14826 23128 14832 23180
rect 14884 23168 14890 23180
rect 17497 23171 17555 23177
rect 17497 23168 17509 23171
rect 14884 23140 17509 23168
rect 14884 23128 14890 23140
rect 17497 23137 17509 23140
rect 17543 23137 17555 23171
rect 17497 23131 17555 23137
rect 25590 23128 25596 23180
rect 25648 23168 25654 23180
rect 25961 23171 26019 23177
rect 25961 23168 25973 23171
rect 25648 23140 25973 23168
rect 25648 23128 25654 23140
rect 25961 23137 25973 23140
rect 26007 23137 26019 23171
rect 29822 23168 29828 23180
rect 29783 23140 29828 23168
rect 25961 23131 26019 23137
rect 29822 23128 29828 23140
rect 29880 23128 29886 23180
rect 10505 23063 10563 23069
rect 12342 23060 12348 23112
rect 12400 23100 12406 23112
rect 12802 23100 12808 23112
rect 12400 23072 12808 23100
rect 12400 23060 12406 23072
rect 12802 23060 12808 23072
rect 12860 23060 12866 23112
rect 12894 23060 12900 23112
rect 12952 23100 12958 23112
rect 15286 23100 15292 23112
rect 12952 23072 15292 23100
rect 12952 23060 12958 23072
rect 15286 23060 15292 23072
rect 15344 23060 15350 23112
rect 15470 23100 15476 23112
rect 15431 23072 15476 23100
rect 15470 23060 15476 23072
rect 15528 23060 15534 23112
rect 18230 23100 18236 23112
rect 16882 23072 18236 23100
rect 18230 23060 18236 23072
rect 18288 23060 18294 23112
rect 18966 23060 18972 23112
rect 19024 23100 19030 23112
rect 19429 23103 19487 23109
rect 19429 23100 19441 23103
rect 19024 23072 19441 23100
rect 19024 23060 19030 23072
rect 19429 23069 19441 23072
rect 19475 23069 19487 23103
rect 19429 23063 19487 23069
rect 20346 23060 20352 23112
rect 20404 23100 20410 23112
rect 20993 23103 21051 23109
rect 20993 23100 21005 23103
rect 20404 23072 21005 23100
rect 20404 23060 20410 23072
rect 20993 23069 21005 23072
rect 21039 23100 21051 23103
rect 21542 23100 21548 23112
rect 21039 23072 21548 23100
rect 21039 23069 21051 23072
rect 20993 23063 21051 23069
rect 21542 23060 21548 23072
rect 21600 23060 21606 23112
rect 26142 23100 26148 23112
rect 26103 23072 26148 23100
rect 26142 23060 26148 23072
rect 26200 23060 26206 23112
rect 28166 23100 28172 23112
rect 28127 23072 28172 23100
rect 28166 23060 28172 23072
rect 28224 23060 28230 23112
rect 28353 23103 28411 23109
rect 28353 23069 28365 23103
rect 28399 23100 28411 23103
rect 28718 23100 28724 23112
rect 28399 23072 28724 23100
rect 28399 23069 28411 23072
rect 28353 23063 28411 23069
rect 28718 23060 28724 23072
rect 28776 23060 28782 23112
rect 1949 23035 2007 23041
rect 1949 23001 1961 23035
rect 1995 23032 2007 23035
rect 2038 23032 2044 23044
rect 1995 23004 2044 23032
rect 1995 23001 2007 23004
rect 1949 22995 2007 23001
rect 2038 22992 2044 23004
rect 2096 22992 2102 23044
rect 3786 23032 3792 23044
rect 3174 23004 3792 23032
rect 3786 22992 3792 23004
rect 3844 22992 3850 23044
rect 6730 22992 6736 23044
rect 6788 22992 6794 23044
rect 12710 22992 12716 23044
rect 12768 23032 12774 23044
rect 13538 23032 13544 23044
rect 12768 23004 13544 23032
rect 12768 22992 12774 23004
rect 13538 22992 13544 23004
rect 13596 22992 13602 23044
rect 15746 23032 15752 23044
rect 15707 23004 15752 23032
rect 15746 22992 15752 23004
rect 15804 22992 15810 23044
rect 17402 22992 17408 23044
rect 17460 23032 17466 23044
rect 18506 23032 18512 23044
rect 17460 23004 18512 23032
rect 17460 22992 17466 23004
rect 18506 22992 18512 23004
rect 18564 23032 18570 23044
rect 19705 23035 19763 23041
rect 19705 23032 19717 23035
rect 18564 23004 19717 23032
rect 18564 22992 18570 23004
rect 19705 23001 19717 23004
rect 19751 23001 19763 23035
rect 29914 23032 29920 23044
rect 29875 23004 29920 23032
rect 19705 22995 19763 23001
rect 29914 22992 29920 23004
rect 29972 22992 29978 23044
rect 30837 23035 30895 23041
rect 30837 23001 30849 23035
rect 30883 23032 30895 23035
rect 32950 23032 32956 23044
rect 30883 23004 32956 23032
rect 30883 23001 30895 23004
rect 30837 22995 30895 23001
rect 32950 22992 32956 23004
rect 33008 23032 33014 23044
rect 35986 23032 35992 23044
rect 33008 23004 35992 23032
rect 33008 22992 33014 23004
rect 35986 22992 35992 23004
rect 36044 22992 36050 23044
rect 3418 22964 3424 22976
rect 3379 22936 3424 22964
rect 3418 22924 3424 22936
rect 3476 22924 3482 22976
rect 7469 22967 7527 22973
rect 7469 22933 7481 22967
rect 7515 22964 7527 22967
rect 7558 22964 7564 22976
rect 7515 22936 7564 22964
rect 7515 22933 7527 22936
rect 7469 22927 7527 22933
rect 7558 22924 7564 22936
rect 7616 22924 7622 22976
rect 12250 22964 12256 22976
rect 12163 22936 12256 22964
rect 12250 22924 12256 22936
rect 12308 22964 12314 22976
rect 17218 22964 17224 22976
rect 12308 22936 17224 22964
rect 12308 22924 12314 22936
rect 17218 22924 17224 22936
rect 17276 22924 17282 22976
rect 17678 22924 17684 22976
rect 17736 22964 17742 22976
rect 21085 22967 21143 22973
rect 21085 22964 21097 22967
rect 17736 22936 21097 22964
rect 17736 22924 17742 22936
rect 21085 22933 21097 22936
rect 21131 22933 21143 22967
rect 21085 22927 21143 22933
rect 26605 22967 26663 22973
rect 26605 22933 26617 22967
rect 26651 22964 26663 22967
rect 28442 22964 28448 22976
rect 26651 22936 28448 22964
rect 26651 22933 26663 22936
rect 26605 22927 26663 22933
rect 28442 22924 28448 22936
rect 28500 22924 28506 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 3329 22763 3387 22769
rect 3329 22729 3341 22763
rect 3375 22760 3387 22763
rect 7466 22760 7472 22772
rect 3375 22732 7472 22760
rect 3375 22729 3387 22732
rect 3329 22723 3387 22729
rect 7466 22720 7472 22732
rect 7524 22760 7530 22772
rect 11054 22760 11060 22772
rect 7524 22732 8708 22760
rect 7524 22720 7530 22732
rect 1394 22652 1400 22704
rect 1452 22692 1458 22704
rect 1857 22695 1915 22701
rect 1857 22692 1869 22695
rect 1452 22664 1869 22692
rect 1452 22652 1458 22664
rect 1857 22661 1869 22664
rect 1903 22661 1915 22695
rect 3142 22692 3148 22704
rect 3082 22664 3148 22692
rect 1857 22655 1915 22661
rect 3142 22652 3148 22664
rect 3200 22652 3206 22704
rect 5534 22652 5540 22704
rect 5592 22652 5598 22704
rect 1578 22556 1584 22568
rect 1539 22528 1584 22556
rect 1578 22516 1584 22528
rect 1636 22516 1642 22568
rect 4249 22559 4307 22565
rect 4249 22525 4261 22559
rect 4295 22525 4307 22559
rect 4249 22519 4307 22525
rect 4525 22559 4583 22565
rect 4525 22525 4537 22559
rect 4571 22556 4583 22559
rect 6822 22556 6828 22568
rect 4571 22528 6828 22556
rect 4571 22525 4583 22528
rect 4525 22519 4583 22525
rect 4264 22420 4292 22519
rect 6822 22516 6828 22528
rect 6880 22516 6886 22568
rect 4706 22420 4712 22432
rect 4264 22392 4712 22420
rect 4706 22380 4712 22392
rect 4764 22380 4770 22432
rect 5994 22420 6000 22432
rect 5955 22392 6000 22420
rect 5994 22380 6000 22392
rect 6052 22380 6058 22432
rect 8680 22420 8708 22732
rect 9600 22732 11060 22760
rect 9600 22701 9628 22732
rect 11054 22720 11060 22732
rect 11112 22720 11118 22772
rect 15470 22760 15476 22772
rect 13280 22732 15476 22760
rect 9585 22695 9643 22701
rect 9585 22661 9597 22695
rect 9631 22661 9643 22695
rect 9585 22655 9643 22661
rect 13280 22633 13308 22732
rect 15470 22720 15476 22732
rect 15528 22720 15534 22772
rect 17218 22720 17224 22772
rect 17276 22760 17282 22772
rect 24578 22760 24584 22772
rect 17276 22732 24584 22760
rect 17276 22720 17282 22732
rect 24578 22720 24584 22732
rect 24636 22720 24642 22772
rect 25777 22763 25835 22769
rect 25777 22729 25789 22763
rect 25823 22760 25835 22763
rect 26142 22760 26148 22772
rect 25823 22732 26148 22760
rect 25823 22729 25835 22732
rect 25777 22723 25835 22729
rect 26142 22720 26148 22732
rect 26200 22720 26206 22772
rect 28718 22760 28724 22772
rect 28679 22732 28724 22760
rect 28718 22720 28724 22732
rect 28776 22720 28782 22772
rect 31113 22763 31171 22769
rect 31113 22729 31125 22763
rect 31159 22760 31171 22763
rect 34698 22760 34704 22772
rect 31159 22732 34704 22760
rect 31159 22729 31171 22732
rect 31113 22723 31171 22729
rect 34698 22720 34704 22732
rect 34756 22720 34762 22772
rect 15286 22692 15292 22704
rect 15199 22664 15292 22692
rect 15286 22652 15292 22664
rect 15344 22692 15350 22704
rect 16574 22692 16580 22704
rect 15344 22664 16580 22692
rect 15344 22652 15350 22664
rect 16574 22652 16580 22664
rect 16632 22692 16638 22704
rect 16632 22664 19564 22692
rect 16632 22652 16638 22664
rect 13265 22627 13323 22633
rect 9122 22516 9128 22568
rect 9180 22556 9186 22568
rect 9309 22559 9367 22565
rect 9309 22556 9321 22559
rect 9180 22528 9321 22556
rect 9180 22516 9186 22528
rect 9309 22525 9321 22528
rect 9355 22525 9367 22559
rect 10704 22556 10732 22610
rect 13265 22593 13277 22627
rect 13311 22593 13323 22627
rect 13265 22587 13323 22593
rect 14642 22584 14648 22636
rect 14700 22584 14706 22636
rect 15212 22596 15516 22624
rect 10704 22528 13400 22556
rect 9309 22519 9367 22525
rect 11057 22491 11115 22497
rect 11057 22457 11069 22491
rect 11103 22488 11115 22491
rect 11882 22488 11888 22500
rect 11103 22460 11888 22488
rect 11103 22457 11115 22460
rect 11057 22451 11115 22457
rect 11882 22448 11888 22460
rect 11940 22488 11946 22500
rect 13262 22488 13268 22500
rect 11940 22460 13268 22488
rect 11940 22448 11946 22460
rect 13262 22448 13268 22460
rect 13320 22448 13326 22500
rect 11422 22420 11428 22432
rect 8680 22392 11428 22420
rect 11422 22380 11428 22392
rect 11480 22380 11486 22432
rect 11514 22380 11520 22432
rect 11572 22420 11578 22432
rect 13170 22420 13176 22432
rect 11572 22392 13176 22420
rect 11572 22380 11578 22392
rect 13170 22380 13176 22392
rect 13228 22380 13234 22432
rect 13372 22420 13400 22528
rect 13538 22516 13544 22568
rect 13596 22556 13602 22568
rect 15212 22556 15240 22596
rect 13596 22528 15240 22556
rect 15488 22556 15516 22596
rect 17034 22584 17040 22636
rect 17092 22624 17098 22636
rect 17865 22627 17923 22633
rect 17865 22624 17877 22627
rect 17092 22596 17877 22624
rect 17092 22584 17098 22596
rect 17865 22593 17877 22596
rect 17911 22593 17923 22627
rect 18506 22624 18512 22636
rect 18467 22596 18512 22624
rect 17865 22587 17923 22593
rect 18506 22584 18512 22596
rect 18564 22584 18570 22636
rect 18966 22584 18972 22636
rect 19024 22624 19030 22636
rect 19429 22627 19487 22633
rect 19429 22624 19441 22627
rect 19024 22596 19441 22624
rect 19024 22584 19030 22596
rect 19429 22593 19441 22596
rect 19475 22593 19487 22627
rect 19536 22624 19564 22664
rect 20622 22652 20628 22704
rect 20680 22692 20686 22704
rect 21177 22695 21235 22701
rect 21177 22692 21189 22695
rect 20680 22664 21189 22692
rect 20680 22652 20686 22664
rect 21177 22661 21189 22664
rect 21223 22661 21235 22695
rect 22186 22692 22192 22704
rect 22147 22664 22192 22692
rect 21177 22655 21235 22661
rect 22186 22652 22192 22664
rect 22244 22652 22250 22704
rect 26513 22695 26571 22701
rect 26513 22661 26525 22695
rect 26559 22692 26571 22695
rect 27341 22695 27399 22701
rect 27341 22692 27353 22695
rect 26559 22664 27353 22692
rect 26559 22661 26571 22664
rect 26513 22655 26571 22661
rect 27341 22661 27353 22664
rect 27387 22661 27399 22695
rect 27341 22655 27399 22661
rect 27798 22652 27804 22704
rect 27856 22692 27862 22704
rect 28074 22692 28080 22704
rect 27856 22664 28080 22692
rect 27856 22652 27862 22664
rect 28074 22652 28080 22664
rect 28132 22692 28138 22704
rect 28261 22695 28319 22701
rect 28261 22692 28273 22695
rect 28132 22664 28273 22692
rect 28132 22652 28138 22664
rect 28261 22661 28273 22664
rect 28307 22661 28319 22695
rect 28261 22655 28319 22661
rect 20806 22624 20812 22636
rect 19536 22596 20812 22624
rect 19429 22587 19487 22593
rect 20806 22584 20812 22596
rect 20864 22584 20870 22636
rect 21085 22627 21143 22633
rect 21085 22624 21097 22627
rect 20916 22596 21097 22624
rect 17770 22556 17776 22568
rect 15488 22528 17776 22556
rect 13596 22516 13602 22528
rect 17770 22516 17776 22528
rect 17828 22516 17834 22568
rect 18414 22516 18420 22568
rect 18472 22556 18478 22568
rect 18785 22559 18843 22565
rect 18785 22556 18797 22559
rect 18472 22528 18797 22556
rect 18472 22516 18478 22528
rect 18785 22525 18797 22528
rect 18831 22556 18843 22559
rect 19150 22556 19156 22568
rect 18831 22528 19156 22556
rect 18831 22525 18843 22528
rect 18785 22519 18843 22525
rect 19150 22516 19156 22528
rect 19208 22516 19214 22568
rect 19610 22556 19616 22568
rect 19571 22528 19616 22556
rect 19610 22516 19616 22528
rect 19668 22516 19674 22568
rect 20530 22516 20536 22568
rect 20588 22556 20594 22568
rect 20916 22556 20944 22596
rect 21085 22593 21097 22596
rect 21131 22593 21143 22627
rect 25958 22624 25964 22636
rect 25919 22596 25964 22624
rect 21085 22587 21143 22593
rect 25958 22584 25964 22596
rect 26016 22584 26022 22636
rect 26421 22627 26479 22633
rect 26421 22593 26433 22627
rect 26467 22593 26479 22627
rect 28902 22624 28908 22636
rect 28863 22596 28908 22624
rect 26421 22587 26479 22593
rect 20588 22528 20944 22556
rect 20588 22516 20594 22528
rect 19978 22488 19984 22500
rect 14568 22460 19984 22488
rect 14568 22420 14596 22460
rect 19978 22448 19984 22460
rect 20036 22448 20042 22500
rect 20916 22488 20944 22528
rect 20990 22516 20996 22568
rect 21048 22556 21054 22568
rect 22097 22559 22155 22565
rect 22097 22556 22109 22559
rect 21048 22528 22109 22556
rect 21048 22516 21054 22528
rect 22097 22525 22109 22528
rect 22143 22525 22155 22559
rect 22097 22519 22155 22525
rect 25774 22516 25780 22568
rect 25832 22556 25838 22568
rect 26436 22556 26464 22587
rect 28902 22584 28908 22596
rect 28960 22584 28966 22636
rect 31294 22624 31300 22636
rect 31255 22596 31300 22624
rect 31294 22584 31300 22596
rect 31352 22584 31358 22636
rect 34422 22624 34428 22636
rect 34383 22596 34428 22624
rect 34422 22584 34428 22596
rect 34480 22584 34486 22636
rect 38013 22627 38071 22633
rect 38013 22593 38025 22627
rect 38059 22593 38071 22627
rect 38013 22587 38071 22593
rect 25832 22528 26464 22556
rect 27249 22559 27307 22565
rect 25832 22516 25838 22528
rect 27249 22525 27261 22559
rect 27295 22556 27307 22559
rect 28074 22556 28080 22568
rect 27295 22528 28080 22556
rect 27295 22525 27307 22528
rect 27249 22519 27307 22525
rect 28074 22516 28080 22528
rect 28132 22516 28138 22568
rect 38028 22556 38056 22587
rect 34256 22528 38056 22556
rect 22462 22488 22468 22500
rect 20916 22460 22468 22488
rect 22462 22448 22468 22460
rect 22520 22448 22526 22500
rect 22646 22488 22652 22500
rect 22607 22460 22652 22488
rect 22646 22448 22652 22460
rect 22704 22448 22710 22500
rect 34256 22497 34284 22528
rect 34241 22491 34299 22497
rect 34241 22457 34253 22491
rect 34287 22457 34299 22491
rect 38194 22488 38200 22500
rect 38155 22460 38200 22488
rect 34241 22451 34299 22457
rect 38194 22448 38200 22460
rect 38252 22448 38258 22500
rect 13372 22392 14596 22420
rect 15838 22380 15844 22432
rect 15896 22420 15902 22432
rect 16482 22420 16488 22432
rect 15896 22392 16488 22420
rect 15896 22380 15902 22392
rect 16482 22380 16488 22392
rect 16540 22380 16546 22432
rect 17957 22423 18015 22429
rect 17957 22389 17969 22423
rect 18003 22420 18015 22423
rect 19334 22420 19340 22432
rect 18003 22392 19340 22420
rect 18003 22389 18015 22392
rect 17957 22383 18015 22389
rect 19334 22380 19340 22392
rect 19392 22380 19398 22432
rect 20162 22380 20168 22432
rect 20220 22420 20226 22432
rect 22094 22420 22100 22432
rect 20220 22392 22100 22420
rect 20220 22380 20226 22392
rect 22094 22380 22100 22392
rect 22152 22380 22158 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 5340 22219 5398 22225
rect 5340 22185 5352 22219
rect 5386 22216 5398 22219
rect 8294 22216 8300 22228
rect 5386 22188 8300 22216
rect 5386 22185 5398 22188
rect 5340 22179 5398 22185
rect 8294 22176 8300 22188
rect 8352 22176 8358 22228
rect 9388 22219 9446 22225
rect 9388 22185 9400 22219
rect 9434 22216 9446 22219
rect 11514 22216 11520 22228
rect 9434 22188 11520 22216
rect 9434 22185 9446 22188
rect 9388 22179 9446 22185
rect 11514 22176 11520 22188
rect 11572 22176 11578 22228
rect 12148 22219 12206 22225
rect 12148 22185 12160 22219
rect 12194 22216 12206 22219
rect 12894 22216 12900 22228
rect 12194 22188 12900 22216
rect 12194 22185 12206 22188
rect 12148 22179 12206 22185
rect 12894 22176 12900 22188
rect 12952 22176 12958 22228
rect 13262 22176 13268 22228
rect 13320 22216 13326 22228
rect 25130 22216 25136 22228
rect 13320 22188 25136 22216
rect 13320 22176 13326 22188
rect 25130 22176 25136 22188
rect 25188 22216 25194 22228
rect 25774 22216 25780 22228
rect 25188 22188 25780 22216
rect 25188 22176 25194 22188
rect 25774 22176 25780 22188
rect 25832 22176 25838 22228
rect 25958 22176 25964 22228
rect 26016 22216 26022 22228
rect 26145 22219 26203 22225
rect 26145 22216 26157 22219
rect 26016 22188 26157 22216
rect 26016 22176 26022 22188
rect 26145 22185 26157 22188
rect 26191 22185 26203 22219
rect 26145 22179 26203 22185
rect 11716 22120 12020 22148
rect 5074 22080 5080 22092
rect 5035 22052 5080 22080
rect 5074 22040 5080 22052
rect 5132 22040 5138 22092
rect 6822 22080 6828 22092
rect 6735 22052 6828 22080
rect 6822 22040 6828 22052
rect 6880 22080 6886 22092
rect 10778 22080 10784 22092
rect 6880 22052 10784 22080
rect 6880 22040 6886 22052
rect 10778 22040 10784 22052
rect 10836 22040 10842 22092
rect 11716 22080 11744 22120
rect 10888 22052 11744 22080
rect 9125 22015 9183 22021
rect 9125 21981 9137 22015
rect 9171 21981 9183 22015
rect 9125 21975 9183 21981
rect 1670 21944 1676 21956
rect 1631 21916 1676 21944
rect 1670 21904 1676 21916
rect 1728 21904 1734 21956
rect 1857 21947 1915 21953
rect 1857 21913 1869 21947
rect 1903 21944 1915 21947
rect 3326 21944 3332 21956
rect 1903 21916 3332 21944
rect 1903 21913 1915 21916
rect 1857 21907 1915 21913
rect 3326 21904 3332 21916
rect 3384 21904 3390 21956
rect 5258 21904 5264 21956
rect 5316 21944 5322 21956
rect 9140 21944 9168 21975
rect 9306 21944 9312 21956
rect 5316 21916 5842 21944
rect 9140 21916 9312 21944
rect 5316 21904 5322 21916
rect 9306 21904 9312 21916
rect 9364 21904 9370 21956
rect 9674 21904 9680 21956
rect 9732 21944 9738 21956
rect 9732 21916 9890 21944
rect 9732 21904 9738 21916
rect 4890 21836 4896 21888
rect 4948 21876 4954 21888
rect 5074 21876 5080 21888
rect 4948 21848 5080 21876
rect 4948 21836 4954 21848
rect 5074 21836 5080 21848
rect 5132 21836 5138 21888
rect 7742 21836 7748 21888
rect 7800 21876 7806 21888
rect 10888 21885 10916 22052
rect 11790 22040 11796 22092
rect 11848 22080 11854 22092
rect 11885 22083 11943 22089
rect 11885 22080 11897 22083
rect 11848 22052 11897 22080
rect 11848 22040 11854 22052
rect 11885 22049 11897 22052
rect 11931 22049 11943 22083
rect 11992 22080 12020 22120
rect 13170 22108 13176 22160
rect 13228 22148 13234 22160
rect 16298 22148 16304 22160
rect 13228 22120 16304 22148
rect 13228 22108 13234 22120
rect 16298 22108 16304 22120
rect 16356 22108 16362 22160
rect 16482 22108 16488 22160
rect 16540 22148 16546 22160
rect 19610 22148 19616 22160
rect 16540 22120 19616 22148
rect 16540 22108 16546 22120
rect 19610 22108 19616 22120
rect 19668 22108 19674 22160
rect 22094 22108 22100 22160
rect 22152 22148 22158 22160
rect 22278 22148 22284 22160
rect 22152 22120 22284 22148
rect 22152 22108 22158 22120
rect 22278 22108 22284 22120
rect 22336 22108 22342 22160
rect 13630 22080 13636 22092
rect 11992 22052 13492 22080
rect 13591 22052 13636 22080
rect 11885 22043 11943 22049
rect 13464 22012 13492 22052
rect 13630 22040 13636 22052
rect 13688 22040 13694 22092
rect 17310 22040 17316 22092
rect 17368 22080 17374 22092
rect 19058 22080 19064 22092
rect 17368 22052 19064 22080
rect 17368 22040 17374 22052
rect 19058 22040 19064 22052
rect 19116 22040 19122 22092
rect 20346 22080 20352 22092
rect 19444 22052 20352 22080
rect 13814 22012 13820 22024
rect 13464 21984 13820 22012
rect 13814 21972 13820 21984
rect 13872 21972 13878 22024
rect 18417 22015 18475 22021
rect 18417 21981 18429 22015
rect 18463 22012 18475 22015
rect 18506 22012 18512 22024
rect 18463 21984 18512 22012
rect 18463 21981 18475 21984
rect 18417 21975 18475 21981
rect 18506 21972 18512 21984
rect 18564 22012 18570 22024
rect 18966 22012 18972 22024
rect 18564 21984 18972 22012
rect 18564 21972 18570 21984
rect 18966 21972 18972 21984
rect 19024 21972 19030 22024
rect 19444 22021 19472 22052
rect 20346 22040 20352 22052
rect 20404 22040 20410 22092
rect 20806 22040 20812 22092
rect 20864 22080 20870 22092
rect 21358 22080 21364 22092
rect 20864 22052 21364 22080
rect 20864 22040 20870 22052
rect 21358 22040 21364 22052
rect 21416 22040 21422 22092
rect 23750 22040 23756 22092
rect 23808 22080 23814 22092
rect 29825 22083 29883 22089
rect 23808 22052 29776 22080
rect 23808 22040 23814 22052
rect 19429 22015 19487 22021
rect 19429 21981 19441 22015
rect 19475 21981 19487 22015
rect 19429 21975 19487 21981
rect 20073 22015 20131 22021
rect 20073 21981 20085 22015
rect 20119 22012 20131 22015
rect 20530 22012 20536 22024
rect 20119 21984 20536 22012
rect 20119 21981 20131 21984
rect 20073 21975 20131 21981
rect 12618 21904 12624 21956
rect 12676 21904 12682 21956
rect 18693 21947 18751 21953
rect 18693 21944 18705 21947
rect 17880 21916 18705 21944
rect 10873 21879 10931 21885
rect 10873 21876 10885 21879
rect 7800 21848 10885 21876
rect 7800 21836 7806 21848
rect 10873 21845 10885 21848
rect 10919 21845 10931 21879
rect 10873 21839 10931 21845
rect 11790 21836 11796 21888
rect 11848 21876 11854 21888
rect 17880 21876 17908 21916
rect 18693 21913 18705 21916
rect 18739 21944 18751 21947
rect 20088 21944 20116 21975
rect 20530 21972 20536 21984
rect 20588 21972 20594 22024
rect 22462 21972 22468 22024
rect 22520 22012 22526 22024
rect 22557 22015 22615 22021
rect 22557 22012 22569 22015
rect 22520 21984 22569 22012
rect 22520 21972 22526 21984
rect 22557 21981 22569 21984
rect 22603 21981 22615 22015
rect 23198 22012 23204 22024
rect 23159 21984 23204 22012
rect 22557 21975 22615 21981
rect 23198 21972 23204 21984
rect 23256 21972 23262 22024
rect 23842 22012 23848 22024
rect 23803 21984 23848 22012
rect 23842 21972 23848 21984
rect 23900 21972 23906 22024
rect 26326 22012 26332 22024
rect 26287 21984 26332 22012
rect 26326 21972 26332 21984
rect 26384 21972 26390 22024
rect 29748 22021 29776 22052
rect 29825 22049 29837 22083
rect 29871 22080 29883 22083
rect 31294 22080 31300 22092
rect 29871 22052 31300 22080
rect 29871 22049 29883 22052
rect 29825 22043 29883 22049
rect 31294 22040 31300 22052
rect 31352 22040 31358 22092
rect 29733 22015 29791 22021
rect 29733 21981 29745 22015
rect 29779 21981 29791 22015
rect 29733 21975 29791 21981
rect 18739 21916 20116 21944
rect 18739 21913 18751 21916
rect 18693 21907 18751 21913
rect 20254 21904 20260 21956
rect 20312 21944 20318 21956
rect 20349 21947 20407 21953
rect 20349 21944 20361 21947
rect 20312 21916 20361 21944
rect 20312 21904 20318 21916
rect 20349 21913 20361 21916
rect 20395 21913 20407 21947
rect 21082 21944 21088 21956
rect 21043 21916 21088 21944
rect 20349 21907 20407 21913
rect 21082 21904 21088 21916
rect 21140 21904 21146 21956
rect 21177 21947 21235 21953
rect 21177 21913 21189 21947
rect 21223 21944 21235 21947
rect 23293 21947 23351 21953
rect 23293 21944 23305 21947
rect 21223 21916 23305 21944
rect 21223 21913 21235 21916
rect 21177 21907 21235 21913
rect 23293 21913 23305 21916
rect 23339 21913 23351 21947
rect 24670 21944 24676 21956
rect 24631 21916 24676 21944
rect 23293 21907 23351 21913
rect 24670 21904 24676 21916
rect 24728 21904 24734 21956
rect 24765 21947 24823 21953
rect 24765 21913 24777 21947
rect 24811 21913 24823 21947
rect 24765 21907 24823 21913
rect 11848 21848 17908 21876
rect 11848 21836 11854 21848
rect 17954 21836 17960 21888
rect 18012 21876 18018 21888
rect 19521 21879 19579 21885
rect 19521 21876 19533 21879
rect 18012 21848 19533 21876
rect 18012 21836 18018 21848
rect 19521 21845 19533 21848
rect 19567 21845 19579 21879
rect 19521 21839 19579 21845
rect 20622 21836 20628 21888
rect 20680 21876 20686 21888
rect 22649 21879 22707 21885
rect 22649 21876 22661 21879
rect 20680 21848 22661 21876
rect 20680 21836 20686 21848
rect 22649 21845 22661 21848
rect 22695 21845 22707 21879
rect 22649 21839 22707 21845
rect 23937 21879 23995 21885
rect 23937 21845 23949 21879
rect 23983 21876 23995 21879
rect 24780 21876 24808 21907
rect 25314 21904 25320 21956
rect 25372 21944 25378 21956
rect 25685 21947 25743 21953
rect 25685 21944 25697 21947
rect 25372 21916 25697 21944
rect 25372 21904 25378 21916
rect 25685 21913 25697 21916
rect 25731 21913 25743 21947
rect 25685 21907 25743 21913
rect 23983 21848 24808 21876
rect 23983 21845 23995 21848
rect 23937 21839 23995 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 5810 21632 5816 21684
rect 5868 21672 5874 21684
rect 5868 21644 7880 21672
rect 5868 21632 5874 21644
rect 5077 21607 5135 21613
rect 5077 21573 5089 21607
rect 5123 21604 5135 21607
rect 6914 21604 6920 21616
rect 5123 21576 6920 21604
rect 5123 21573 5135 21576
rect 5077 21567 5135 21573
rect 6914 21564 6920 21576
rect 6972 21564 6978 21616
rect 7742 21604 7748 21616
rect 7703 21576 7748 21604
rect 7742 21564 7748 21576
rect 7800 21564 7806 21616
rect 7852 21604 7880 21644
rect 10134 21632 10140 21684
rect 10192 21672 10198 21684
rect 16206 21672 16212 21684
rect 10192 21644 16212 21672
rect 10192 21632 10198 21644
rect 16206 21632 16212 21644
rect 16264 21632 16270 21684
rect 20806 21672 20812 21684
rect 16316 21644 20812 21672
rect 7852 21576 8234 21604
rect 16114 21564 16120 21616
rect 16172 21604 16178 21616
rect 16316 21604 16344 21644
rect 20806 21632 20812 21644
rect 20864 21632 20870 21684
rect 21082 21632 21088 21684
rect 21140 21672 21146 21684
rect 21269 21675 21327 21681
rect 21269 21672 21281 21675
rect 21140 21644 21281 21672
rect 21140 21632 21146 21644
rect 21269 21641 21281 21644
rect 21315 21641 21327 21675
rect 21269 21635 21327 21641
rect 21358 21632 21364 21684
rect 21416 21672 21422 21684
rect 23750 21672 23756 21684
rect 21416 21644 23756 21672
rect 21416 21632 21422 21644
rect 23750 21632 23756 21644
rect 23808 21632 23814 21684
rect 24026 21672 24032 21684
rect 23987 21644 24032 21672
rect 24026 21632 24032 21644
rect 24084 21632 24090 21684
rect 31481 21675 31539 21681
rect 31481 21641 31493 21675
rect 31527 21672 31539 21675
rect 38010 21672 38016 21684
rect 31527 21644 38016 21672
rect 31527 21641 31539 21644
rect 31481 21635 31539 21641
rect 38010 21632 38016 21644
rect 38068 21632 38074 21684
rect 16172 21576 16344 21604
rect 16172 21564 16178 21576
rect 16390 21564 16396 21616
rect 16448 21604 16454 21616
rect 23198 21604 23204 21616
rect 16448 21576 23204 21604
rect 16448 21564 16454 21576
rect 23198 21564 23204 21576
rect 23256 21564 23262 21616
rect 35894 21604 35900 21616
rect 29196 21576 35900 21604
rect 15838 21496 15844 21548
rect 15896 21496 15902 21548
rect 18322 21536 18328 21548
rect 18283 21508 18328 21536
rect 18322 21496 18328 21508
rect 18380 21496 18386 21548
rect 18966 21536 18972 21548
rect 18879 21508 18972 21536
rect 18966 21496 18972 21508
rect 19024 21536 19030 21548
rect 19889 21539 19947 21545
rect 19889 21536 19901 21539
rect 19024 21508 19901 21536
rect 19024 21496 19030 21508
rect 19889 21505 19901 21508
rect 19935 21536 19947 21539
rect 20346 21536 20352 21548
rect 19935 21508 20352 21536
rect 19935 21505 19947 21508
rect 19889 21499 19947 21505
rect 20346 21496 20352 21508
rect 20404 21496 20410 21548
rect 20530 21496 20536 21548
rect 20588 21536 20594 21548
rect 22005 21539 22063 21545
rect 22005 21536 22017 21539
rect 20588 21508 22017 21536
rect 20588 21496 20594 21508
rect 22005 21505 22017 21508
rect 22051 21505 22063 21539
rect 23290 21536 23296 21548
rect 22005 21499 22063 21505
rect 22112 21508 23296 21536
rect 4798 21428 4804 21480
rect 4856 21468 4862 21480
rect 5813 21471 5871 21477
rect 5813 21468 5825 21471
rect 4856 21440 5825 21468
rect 4856 21428 4862 21440
rect 5813 21437 5825 21440
rect 5859 21437 5871 21471
rect 5813 21431 5871 21437
rect 6546 21428 6552 21480
rect 6604 21468 6610 21480
rect 7469 21471 7527 21477
rect 7469 21468 7481 21471
rect 6604 21440 7481 21468
rect 6604 21428 6610 21440
rect 7469 21437 7481 21440
rect 7515 21468 7527 21471
rect 9122 21468 9128 21480
rect 7515 21440 9128 21468
rect 7515 21437 7527 21440
rect 7469 21431 7527 21437
rect 9122 21428 9128 21440
rect 9180 21428 9186 21480
rect 14458 21468 14464 21480
rect 14419 21440 14464 21468
rect 14458 21428 14464 21440
rect 14516 21428 14522 21480
rect 15194 21428 15200 21480
rect 15252 21468 15258 21480
rect 15252 21440 16252 21468
rect 15252 21428 15258 21440
rect 16224 21409 16252 21440
rect 18874 21428 18880 21480
rect 18932 21468 18938 21480
rect 19058 21468 19064 21480
rect 18932 21440 19064 21468
rect 18932 21428 18938 21440
rect 19058 21428 19064 21440
rect 19116 21468 19122 21480
rect 19153 21471 19211 21477
rect 19153 21468 19165 21471
rect 19116 21440 19165 21468
rect 19116 21428 19122 21440
rect 19153 21437 19165 21440
rect 19199 21437 19211 21471
rect 19153 21431 19211 21437
rect 19242 21428 19248 21480
rect 19300 21468 19306 21480
rect 20625 21471 20683 21477
rect 20625 21468 20637 21471
rect 19300 21440 20637 21468
rect 19300 21428 19306 21440
rect 20625 21437 20637 21440
rect 20671 21437 20683 21471
rect 20625 21431 20683 21437
rect 20714 21428 20720 21480
rect 20772 21468 20778 21480
rect 22112 21468 22140 21508
rect 23290 21496 23296 21508
rect 23348 21496 23354 21548
rect 23937 21539 23995 21545
rect 23937 21505 23949 21539
rect 23983 21505 23995 21539
rect 24578 21536 24584 21548
rect 24539 21508 24584 21536
rect 23937 21499 23995 21505
rect 22278 21468 22284 21480
rect 20772 21440 22140 21468
rect 22239 21440 22284 21468
rect 20772 21428 20778 21440
rect 22278 21428 22284 21440
rect 22336 21428 22342 21480
rect 23952 21468 23980 21499
rect 24578 21496 24584 21508
rect 24636 21496 24642 21548
rect 28074 21536 28080 21548
rect 28035 21508 28080 21536
rect 28074 21496 28080 21508
rect 28132 21496 28138 21548
rect 29196 21545 29224 21576
rect 35894 21564 35900 21576
rect 35952 21564 35958 21616
rect 29181 21539 29239 21545
rect 29181 21505 29193 21539
rect 29227 21505 29239 21539
rect 31662 21536 31668 21548
rect 31623 21508 31668 21536
rect 29181 21499 29239 21505
rect 31662 21496 31668 21508
rect 31720 21496 31726 21548
rect 37826 21496 37832 21548
rect 37884 21536 37890 21548
rect 38013 21539 38071 21545
rect 38013 21536 38025 21539
rect 37884 21508 38025 21536
rect 37884 21496 37890 21508
rect 38013 21505 38025 21508
rect 38059 21505 38071 21539
rect 38013 21499 38071 21505
rect 22756 21440 23980 21468
rect 22756 21412 22784 21440
rect 26234 21428 26240 21480
rect 26292 21468 26298 21480
rect 28261 21471 28319 21477
rect 28261 21468 28273 21471
rect 26292 21440 28273 21468
rect 26292 21428 26298 21440
rect 28261 21437 28273 21440
rect 28307 21437 28319 21471
rect 28261 21431 28319 21437
rect 16209 21403 16267 21409
rect 16209 21369 16221 21403
rect 16255 21400 16267 21403
rect 22738 21400 22744 21412
rect 16255 21372 22744 21400
rect 16255 21369 16267 21372
rect 16209 21363 16267 21369
rect 22738 21360 22744 21372
rect 22796 21360 22802 21412
rect 28442 21400 28448 21412
rect 28403 21372 28448 21400
rect 28442 21360 28448 21372
rect 28500 21360 28506 21412
rect 9217 21335 9275 21341
rect 9217 21301 9229 21335
rect 9263 21332 9275 21335
rect 9766 21332 9772 21344
rect 9263 21304 9772 21332
rect 9263 21301 9275 21304
rect 9217 21295 9275 21301
rect 9766 21292 9772 21304
rect 9824 21292 9830 21344
rect 14724 21335 14782 21341
rect 14724 21301 14736 21335
rect 14770 21332 14782 21335
rect 17126 21332 17132 21344
rect 14770 21304 17132 21332
rect 14770 21301 14782 21304
rect 14724 21295 14782 21301
rect 17126 21292 17132 21304
rect 17184 21292 17190 21344
rect 18414 21332 18420 21344
rect 18375 21304 18420 21332
rect 18414 21292 18420 21304
rect 18472 21292 18478 21344
rect 19702 21292 19708 21344
rect 19760 21332 19766 21344
rect 20806 21332 20812 21344
rect 19760 21304 20812 21332
rect 19760 21292 19766 21304
rect 20806 21292 20812 21304
rect 20864 21292 20870 21344
rect 20898 21292 20904 21344
rect 20956 21332 20962 21344
rect 23385 21335 23443 21341
rect 23385 21332 23397 21335
rect 20956 21304 23397 21332
rect 20956 21292 20962 21304
rect 23385 21301 23397 21304
rect 23431 21301 23443 21335
rect 23385 21295 23443 21301
rect 23658 21292 23664 21344
rect 23716 21332 23722 21344
rect 24673 21335 24731 21341
rect 24673 21332 24685 21335
rect 23716 21304 24685 21332
rect 23716 21292 23722 21304
rect 24673 21301 24685 21304
rect 24719 21301 24731 21335
rect 24673 21295 24731 21301
rect 27430 21292 27436 21344
rect 27488 21332 27494 21344
rect 29273 21335 29331 21341
rect 29273 21332 29285 21335
rect 27488 21304 29285 21332
rect 27488 21292 27494 21304
rect 29273 21301 29285 21304
rect 29319 21301 29331 21335
rect 38194 21332 38200 21344
rect 38155 21304 38200 21332
rect 29273 21295 29331 21301
rect 38194 21292 38200 21304
rect 38252 21292 38258 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 5340 21131 5398 21137
rect 5340 21097 5352 21131
rect 5386 21128 5398 21131
rect 8202 21128 8208 21140
rect 5386 21100 8208 21128
rect 5386 21097 5398 21100
rect 5340 21091 5398 21097
rect 8202 21088 8208 21100
rect 8260 21128 8266 21140
rect 12434 21128 12440 21140
rect 8260 21100 12440 21128
rect 8260 21088 8266 21100
rect 12434 21088 12440 21100
rect 12492 21088 12498 21140
rect 15838 21088 15844 21140
rect 15896 21128 15902 21140
rect 21269 21131 21327 21137
rect 21269 21128 21281 21131
rect 15896 21100 21281 21128
rect 15896 21088 15902 21100
rect 21269 21097 21281 21100
rect 21315 21097 21327 21131
rect 21269 21091 21327 21097
rect 28074 21088 28080 21140
rect 28132 21128 28138 21140
rect 28353 21131 28411 21137
rect 28353 21128 28365 21131
rect 28132 21100 28365 21128
rect 28132 21088 28138 21100
rect 28353 21097 28365 21100
rect 28399 21097 28411 21131
rect 29086 21128 29092 21140
rect 29047 21100 29092 21128
rect 28353 21091 28411 21097
rect 29086 21088 29092 21100
rect 29144 21088 29150 21140
rect 14826 21060 14832 21072
rect 12406 21032 14832 21060
rect 5077 20995 5135 21001
rect 5077 20961 5089 20995
rect 5123 20992 5135 20995
rect 6546 20992 6552 21004
rect 5123 20964 6552 20992
rect 5123 20961 5135 20964
rect 5077 20955 5135 20961
rect 6546 20952 6552 20964
rect 6604 20952 6610 21004
rect 6638 20952 6644 21004
rect 6696 20992 6702 21004
rect 6825 20995 6883 21001
rect 6825 20992 6837 20995
rect 6696 20964 6837 20992
rect 6696 20952 6702 20964
rect 6825 20961 6837 20964
rect 6871 20961 6883 20995
rect 9122 20992 9128 21004
rect 9083 20964 9128 20992
rect 6825 20955 6883 20961
rect 9122 20952 9128 20964
rect 9180 20952 9186 21004
rect 9401 20995 9459 21001
rect 9401 20961 9413 20995
rect 9447 20992 9459 20995
rect 12406 20992 12434 21032
rect 14826 21020 14832 21032
rect 14884 21020 14890 21072
rect 16669 21063 16727 21069
rect 16669 21029 16681 21063
rect 16715 21060 16727 21063
rect 16758 21060 16764 21072
rect 16715 21032 16764 21060
rect 16715 21029 16727 21032
rect 16669 21023 16727 21029
rect 16758 21020 16764 21032
rect 16816 21060 16822 21072
rect 20714 21060 20720 21072
rect 16816 21032 20720 21060
rect 16816 21020 16822 21032
rect 20714 21020 20720 21032
rect 20772 21020 20778 21072
rect 27338 21060 27344 21072
rect 23676 21032 27344 21060
rect 20162 20992 20168 21004
rect 9447 20964 12434 20992
rect 14384 20964 20168 20992
rect 9447 20961 9459 20964
rect 9401 20955 9459 20961
rect 9030 20924 9036 20936
rect 6486 20896 9036 20924
rect 9030 20884 9036 20896
rect 9088 20884 9094 20936
rect 1670 20856 1676 20868
rect 1631 20828 1676 20856
rect 1670 20816 1676 20828
rect 1728 20816 1734 20868
rect 6748 20828 7144 20856
rect 1765 20791 1823 20797
rect 1765 20757 1777 20791
rect 1811 20788 1823 20791
rect 6748 20788 6776 20828
rect 1811 20760 6776 20788
rect 7116 20788 7144 20828
rect 10410 20816 10416 20868
rect 10468 20816 10474 20868
rect 10704 20828 12434 20856
rect 10704 20788 10732 20828
rect 7116 20760 10732 20788
rect 10873 20791 10931 20797
rect 1811 20757 1823 20760
rect 1765 20751 1823 20757
rect 10873 20757 10885 20791
rect 10919 20788 10931 20791
rect 12158 20788 12164 20800
rect 10919 20760 12164 20788
rect 10919 20757 10931 20760
rect 10873 20751 10931 20757
rect 12158 20748 12164 20760
rect 12216 20748 12222 20800
rect 12406 20788 12434 20828
rect 14384 20788 14412 20964
rect 20162 20952 20168 20964
rect 20220 20952 20226 21004
rect 20530 20992 20536 21004
rect 20491 20964 20536 20992
rect 20530 20952 20536 20964
rect 20588 20992 20594 21004
rect 23676 20992 23704 21032
rect 27338 21020 27344 21032
rect 27396 21020 27402 21072
rect 38102 21060 38108 21072
rect 29012 21032 38108 21060
rect 20588 20964 23704 20992
rect 20588 20952 20594 20964
rect 23750 20952 23756 21004
rect 23808 20992 23814 21004
rect 24670 20992 24676 21004
rect 23808 20964 24676 20992
rect 23808 20952 23814 20964
rect 24670 20952 24676 20964
rect 24728 20952 24734 21004
rect 25869 20995 25927 21001
rect 25869 20961 25881 20995
rect 25915 20992 25927 20995
rect 27430 20992 27436 21004
rect 25915 20964 27436 20992
rect 25915 20961 25927 20964
rect 25869 20955 25927 20961
rect 27430 20952 27436 20964
rect 27488 20952 27494 21004
rect 14458 20884 14464 20936
rect 14516 20924 14522 20936
rect 14921 20927 14979 20933
rect 14921 20924 14933 20927
rect 14516 20896 14933 20924
rect 14516 20884 14522 20896
rect 14921 20893 14933 20896
rect 14967 20893 14979 20927
rect 14921 20887 14979 20893
rect 14936 20856 14964 20887
rect 17770 20884 17776 20936
rect 17828 20924 17834 20936
rect 18509 20927 18567 20933
rect 18509 20924 18521 20927
rect 17828 20896 18521 20924
rect 17828 20884 17834 20896
rect 18509 20893 18521 20896
rect 18555 20893 18567 20927
rect 21174 20924 21180 20936
rect 21135 20896 21180 20924
rect 18509 20887 18567 20893
rect 21174 20884 21180 20896
rect 21232 20884 21238 20936
rect 28261 20927 28319 20933
rect 28261 20893 28273 20927
rect 28307 20924 28319 20927
rect 28626 20924 28632 20936
rect 28307 20896 28632 20924
rect 28307 20893 28319 20896
rect 28261 20887 28319 20893
rect 28626 20884 28632 20896
rect 28684 20884 28690 20936
rect 29012 20933 29040 21032
rect 38102 21020 38108 21032
rect 38160 21020 38166 21072
rect 30009 20995 30067 21001
rect 30009 20961 30021 20995
rect 30055 20992 30067 20995
rect 31021 20995 31079 21001
rect 31021 20992 31033 20995
rect 30055 20964 31033 20992
rect 30055 20961 30067 20964
rect 30009 20955 30067 20961
rect 31021 20961 31033 20964
rect 31067 20961 31079 20995
rect 31021 20955 31079 20961
rect 28997 20927 29055 20933
rect 28997 20893 29009 20927
rect 29043 20893 29055 20927
rect 28997 20887 29055 20893
rect 29825 20927 29883 20933
rect 29825 20893 29837 20927
rect 29871 20893 29883 20927
rect 30926 20924 30932 20936
rect 30887 20896 30932 20924
rect 29825 20887 29883 20893
rect 15102 20856 15108 20868
rect 14936 20828 15108 20856
rect 15102 20816 15108 20828
rect 15160 20816 15166 20868
rect 15197 20859 15255 20865
rect 15197 20825 15209 20859
rect 15243 20825 15255 20859
rect 17678 20856 17684 20868
rect 16422 20828 17684 20856
rect 15197 20819 15255 20825
rect 12406 20760 14412 20788
rect 15212 20788 15240 20819
rect 17678 20816 17684 20828
rect 17736 20816 17742 20868
rect 19702 20856 19708 20868
rect 17788 20828 18736 20856
rect 19663 20828 19708 20856
rect 17034 20788 17040 20800
rect 15212 20760 17040 20788
rect 17034 20748 17040 20760
rect 17092 20748 17098 20800
rect 17126 20748 17132 20800
rect 17184 20788 17190 20800
rect 17788 20788 17816 20828
rect 17184 20760 17816 20788
rect 17184 20748 17190 20760
rect 18322 20748 18328 20800
rect 18380 20788 18386 20800
rect 18601 20791 18659 20797
rect 18601 20788 18613 20791
rect 18380 20760 18613 20788
rect 18380 20748 18386 20760
rect 18601 20757 18613 20760
rect 18647 20757 18659 20791
rect 18708 20788 18736 20828
rect 19702 20816 19708 20828
rect 19760 20816 19766 20868
rect 19797 20859 19855 20865
rect 19797 20825 19809 20859
rect 19843 20856 19855 20859
rect 20622 20856 20628 20868
rect 19843 20828 20628 20856
rect 19843 20825 19855 20828
rect 19797 20819 19855 20825
rect 20622 20816 20628 20828
rect 20680 20816 20686 20868
rect 23014 20856 23020 20868
rect 21100 20828 23020 20856
rect 21100 20788 21128 20828
rect 23014 20816 23020 20828
rect 23072 20816 23078 20868
rect 23106 20816 23112 20868
rect 23164 20856 23170 20868
rect 25961 20859 26019 20865
rect 23164 20828 24992 20856
rect 23164 20816 23170 20828
rect 18708 20760 21128 20788
rect 18601 20751 18659 20757
rect 21174 20748 21180 20800
rect 21232 20788 21238 20800
rect 22278 20788 22284 20800
rect 21232 20760 22284 20788
rect 21232 20748 21238 20760
rect 22278 20748 22284 20760
rect 22336 20748 22342 20800
rect 23566 20748 23572 20800
rect 23624 20788 23630 20800
rect 24854 20788 24860 20800
rect 23624 20760 24860 20788
rect 23624 20748 23630 20760
rect 24854 20748 24860 20760
rect 24912 20748 24918 20800
rect 24964 20788 24992 20828
rect 25961 20825 25973 20859
rect 26007 20856 26019 20859
rect 26786 20856 26792 20868
rect 26007 20828 26792 20856
rect 26007 20825 26019 20828
rect 25961 20819 26019 20825
rect 26786 20816 26792 20828
rect 26844 20816 26850 20868
rect 26881 20859 26939 20865
rect 26881 20825 26893 20859
rect 26927 20825 26939 20859
rect 26881 20819 26939 20825
rect 26896 20788 26924 20819
rect 28442 20816 28448 20868
rect 28500 20856 28506 20868
rect 29840 20856 29868 20887
rect 30926 20884 30932 20896
rect 30984 20884 30990 20936
rect 31754 20924 31760 20936
rect 31715 20896 31760 20924
rect 31754 20884 31760 20896
rect 31812 20884 31818 20936
rect 37182 20884 37188 20936
rect 37240 20924 37246 20936
rect 37461 20927 37519 20933
rect 37461 20924 37473 20927
rect 37240 20896 37473 20924
rect 37240 20884 37246 20896
rect 37461 20893 37473 20896
rect 37507 20893 37519 20927
rect 37734 20924 37740 20936
rect 37695 20896 37740 20924
rect 37461 20887 37519 20893
rect 37734 20884 37740 20896
rect 37792 20884 37798 20936
rect 28500 20828 29868 20856
rect 30469 20859 30527 20865
rect 28500 20816 28506 20828
rect 30469 20825 30481 20859
rect 30515 20856 30527 20859
rect 31846 20856 31852 20868
rect 30515 20828 31852 20856
rect 30515 20825 30527 20828
rect 30469 20819 30527 20825
rect 31846 20816 31852 20828
rect 31904 20816 31910 20868
rect 31570 20788 31576 20800
rect 24964 20760 26924 20788
rect 31531 20760 31576 20788
rect 31570 20748 31576 20760
rect 31628 20748 31634 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 10686 20544 10692 20596
rect 10744 20584 10750 20596
rect 17954 20584 17960 20596
rect 10744 20556 17960 20584
rect 10744 20544 10750 20556
rect 17954 20544 17960 20556
rect 18012 20544 18018 20596
rect 20438 20544 20444 20596
rect 20496 20584 20502 20596
rect 20622 20584 20628 20596
rect 20496 20556 20628 20584
rect 20496 20544 20502 20556
rect 20622 20544 20628 20556
rect 20680 20544 20686 20596
rect 22097 20587 22155 20593
rect 22097 20553 22109 20587
rect 22143 20584 22155 20587
rect 22186 20584 22192 20596
rect 22143 20556 22192 20584
rect 22143 20553 22155 20556
rect 22097 20547 22155 20553
rect 22186 20544 22192 20556
rect 22244 20544 22250 20596
rect 25777 20587 25835 20593
rect 25777 20553 25789 20587
rect 25823 20584 25835 20587
rect 26234 20584 26240 20596
rect 25823 20556 26240 20584
rect 25823 20553 25835 20556
rect 25777 20547 25835 20553
rect 26234 20544 26240 20556
rect 26292 20544 26298 20596
rect 26786 20544 26792 20596
rect 26844 20584 26850 20596
rect 27985 20587 28043 20593
rect 27985 20584 27997 20587
rect 26844 20556 27997 20584
rect 26844 20544 26850 20556
rect 27985 20553 27997 20556
rect 28031 20553 28043 20587
rect 27985 20547 28043 20553
rect 30469 20587 30527 20593
rect 30469 20553 30481 20587
rect 30515 20584 30527 20587
rect 31754 20584 31760 20596
rect 30515 20556 31760 20584
rect 30515 20553 30527 20556
rect 30469 20547 30527 20553
rect 31754 20544 31760 20556
rect 31812 20544 31818 20596
rect 6914 20476 6920 20528
rect 6972 20516 6978 20528
rect 8205 20519 8263 20525
rect 8205 20516 8217 20519
rect 6972 20488 8217 20516
rect 6972 20476 6978 20488
rect 8205 20485 8217 20488
rect 8251 20485 8263 20519
rect 8205 20479 8263 20485
rect 9033 20519 9091 20525
rect 9033 20485 9045 20519
rect 9079 20516 9091 20519
rect 9122 20516 9128 20528
rect 9079 20488 9128 20516
rect 9079 20485 9091 20488
rect 9033 20479 9091 20485
rect 1762 20448 1768 20460
rect 1723 20420 1768 20448
rect 1762 20408 1768 20420
rect 1820 20408 1826 20460
rect 7466 20448 7472 20460
rect 4094 20420 7472 20448
rect 7466 20408 7472 20420
rect 7524 20408 7530 20460
rect 8220 20448 8248 20479
rect 9122 20476 9128 20488
rect 9180 20476 9186 20528
rect 13725 20519 13783 20525
rect 13725 20516 13737 20519
rect 11716 20488 13737 20516
rect 11716 20457 11744 20488
rect 13725 20485 13737 20488
rect 13771 20485 13783 20519
rect 13725 20479 13783 20485
rect 17402 20476 17408 20528
rect 17460 20516 17466 20528
rect 17460 20488 27292 20516
rect 17460 20476 17466 20488
rect 27264 20460 27292 20488
rect 11701 20451 11759 20457
rect 11701 20448 11713 20451
rect 8220 20420 11713 20448
rect 11701 20417 11713 20420
rect 11747 20417 11759 20451
rect 11701 20411 11759 20417
rect 17034 20408 17040 20460
rect 17092 20448 17098 20460
rect 18138 20448 18144 20460
rect 17092 20420 18144 20448
rect 17092 20408 17098 20420
rect 18138 20408 18144 20420
rect 18196 20408 18202 20460
rect 20346 20448 20352 20460
rect 20307 20420 20352 20448
rect 20346 20408 20352 20420
rect 20404 20408 20410 20460
rect 22005 20451 22063 20457
rect 22005 20448 22017 20451
rect 20456 20420 22017 20448
rect 1578 20340 1584 20392
rect 1636 20380 1642 20392
rect 2685 20383 2743 20389
rect 2685 20380 2697 20383
rect 1636 20352 2697 20380
rect 1636 20340 1642 20352
rect 2685 20349 2697 20352
rect 2731 20349 2743 20383
rect 2685 20343 2743 20349
rect 2961 20383 3019 20389
rect 2961 20349 2973 20383
rect 3007 20380 3019 20383
rect 3050 20380 3056 20392
rect 3007 20352 3056 20380
rect 3007 20349 3019 20352
rect 2961 20343 3019 20349
rect 3050 20340 3056 20352
rect 3108 20340 3114 20392
rect 11974 20340 11980 20392
rect 12032 20380 12038 20392
rect 12437 20383 12495 20389
rect 12437 20380 12449 20383
rect 12032 20352 12449 20380
rect 12032 20340 12038 20352
rect 12437 20349 12449 20352
rect 12483 20349 12495 20383
rect 12437 20343 12495 20349
rect 14553 20383 14611 20389
rect 14553 20349 14565 20383
rect 14599 20380 14611 20383
rect 15102 20380 15108 20392
rect 14599 20352 15108 20380
rect 14599 20349 14611 20352
rect 14553 20343 14611 20349
rect 15102 20340 15108 20352
rect 15160 20340 15166 20392
rect 17494 20340 17500 20392
rect 17552 20380 17558 20392
rect 20456 20380 20484 20420
rect 22005 20417 22017 20420
rect 22051 20417 22063 20451
rect 22005 20411 22063 20417
rect 25685 20451 25743 20457
rect 25685 20417 25697 20451
rect 25731 20448 25743 20451
rect 26326 20448 26332 20460
rect 25731 20420 26332 20448
rect 25731 20417 25743 20420
rect 25685 20411 25743 20417
rect 20622 20380 20628 20392
rect 17552 20352 20484 20380
rect 20583 20352 20628 20380
rect 17552 20340 17558 20352
rect 20622 20340 20628 20352
rect 20680 20340 20686 20392
rect 21910 20340 21916 20392
rect 21968 20380 21974 20392
rect 25700 20380 25728 20411
rect 26326 20408 26332 20420
rect 26384 20408 26390 20460
rect 27246 20448 27252 20460
rect 27159 20420 27252 20448
rect 27246 20408 27252 20420
rect 27304 20408 27310 20460
rect 27890 20457 27896 20460
rect 27885 20448 27896 20457
rect 27851 20420 27896 20448
rect 27885 20411 27896 20420
rect 27890 20408 27896 20411
rect 27948 20408 27954 20460
rect 28626 20448 28632 20460
rect 28587 20420 28632 20448
rect 28626 20408 28632 20420
rect 28684 20408 28690 20460
rect 30653 20451 30711 20457
rect 30653 20417 30665 20451
rect 30699 20448 30711 20451
rect 30926 20448 30932 20460
rect 30699 20420 30932 20448
rect 30699 20417 30711 20420
rect 30653 20411 30711 20417
rect 30926 20408 30932 20420
rect 30984 20408 30990 20460
rect 31297 20451 31355 20457
rect 31297 20417 31309 20451
rect 31343 20448 31355 20451
rect 31570 20448 31576 20460
rect 31343 20420 31576 20448
rect 31343 20417 31355 20420
rect 31297 20411 31355 20417
rect 31570 20408 31576 20420
rect 31628 20408 31634 20460
rect 31757 20451 31815 20457
rect 31757 20417 31769 20451
rect 31803 20448 31815 20451
rect 31846 20448 31852 20460
rect 31803 20420 31852 20448
rect 31803 20417 31815 20420
rect 31757 20411 31815 20417
rect 31846 20408 31852 20420
rect 31904 20408 31910 20460
rect 31110 20380 31116 20392
rect 21968 20352 25728 20380
rect 31071 20352 31116 20380
rect 21968 20340 21974 20352
rect 31110 20340 31116 20352
rect 31168 20340 31174 20392
rect 9398 20272 9404 20324
rect 9456 20312 9462 20324
rect 28813 20315 28871 20321
rect 28813 20312 28825 20315
rect 9456 20284 28825 20312
rect 9456 20272 9462 20284
rect 28813 20281 28825 20284
rect 28859 20281 28871 20315
rect 28813 20275 28871 20281
rect 1581 20247 1639 20253
rect 1581 20213 1593 20247
rect 1627 20244 1639 20247
rect 2130 20244 2136 20256
rect 1627 20216 2136 20244
rect 1627 20213 1639 20216
rect 1581 20207 1639 20213
rect 2130 20204 2136 20216
rect 2188 20204 2194 20256
rect 4433 20247 4491 20253
rect 4433 20213 4445 20247
rect 4479 20244 4491 20247
rect 5350 20244 5356 20256
rect 4479 20216 5356 20244
rect 4479 20213 4491 20216
rect 4433 20207 4491 20213
rect 5350 20204 5356 20216
rect 5408 20204 5414 20256
rect 5626 20204 5632 20256
rect 5684 20244 5690 20256
rect 8478 20244 8484 20256
rect 5684 20216 8484 20244
rect 5684 20204 5690 20216
rect 8478 20204 8484 20216
rect 8536 20204 8542 20256
rect 27341 20247 27399 20253
rect 27341 20213 27353 20247
rect 27387 20244 27399 20247
rect 27522 20244 27528 20256
rect 27387 20216 27528 20244
rect 27387 20213 27399 20216
rect 27341 20207 27399 20213
rect 27522 20204 27528 20216
rect 27580 20204 27586 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 3326 20000 3332 20052
rect 3384 20040 3390 20052
rect 19978 20040 19984 20052
rect 3384 20012 19984 20040
rect 3384 20000 3390 20012
rect 19978 20000 19984 20012
rect 20036 20000 20042 20052
rect 26878 20040 26884 20052
rect 22204 20012 26884 20040
rect 3421 19975 3479 19981
rect 3421 19941 3433 19975
rect 3467 19972 3479 19975
rect 14550 19972 14556 19984
rect 3467 19944 5672 19972
rect 3467 19941 3479 19944
rect 3421 19935 3479 19941
rect 1949 19907 2007 19913
rect 1949 19873 1961 19907
rect 1995 19904 2007 19907
rect 3970 19904 3976 19916
rect 1995 19876 3976 19904
rect 1995 19873 2007 19876
rect 1949 19867 2007 19873
rect 3970 19864 3976 19876
rect 4028 19864 4034 19916
rect 1578 19796 1584 19848
rect 1636 19836 1642 19848
rect 1673 19839 1731 19845
rect 1673 19836 1685 19839
rect 1636 19808 1685 19836
rect 1636 19796 1642 19808
rect 1673 19805 1685 19808
rect 1719 19805 1731 19839
rect 1673 19799 1731 19805
rect 5534 19768 5540 19780
rect 3174 19740 5540 19768
rect 5534 19728 5540 19740
rect 5592 19728 5598 19780
rect 5644 19768 5672 19944
rect 13004 19944 14556 19972
rect 5905 19907 5963 19913
rect 5905 19873 5917 19907
rect 5951 19904 5963 19907
rect 6546 19904 6552 19916
rect 5951 19876 6552 19904
rect 5951 19873 5963 19876
rect 5905 19867 5963 19873
rect 6546 19864 6552 19876
rect 6604 19864 6610 19916
rect 11609 19907 11667 19913
rect 11609 19904 11621 19907
rect 9324 19876 11621 19904
rect 9324 19848 9352 19876
rect 11609 19873 11621 19876
rect 11655 19904 11667 19907
rect 11974 19904 11980 19916
rect 11655 19876 11980 19904
rect 11655 19873 11667 19876
rect 11609 19867 11667 19873
rect 11974 19864 11980 19876
rect 12032 19864 12038 19916
rect 9306 19836 9312 19848
rect 9267 19808 9312 19836
rect 9306 19796 9312 19808
rect 9364 19796 9370 19848
rect 10686 19796 10692 19848
rect 10744 19796 10750 19848
rect 13004 19822 13032 19944
rect 14550 19932 14556 19944
rect 14608 19932 14614 19984
rect 21910 19972 21916 19984
rect 16408 19944 21916 19972
rect 13357 19907 13415 19913
rect 13357 19873 13369 19907
rect 13403 19904 13415 19907
rect 16408 19904 16436 19944
rect 21910 19932 21916 19944
rect 21968 19932 21974 19984
rect 13403 19876 16436 19904
rect 20533 19907 20591 19913
rect 13403 19873 13415 19876
rect 13357 19867 13415 19873
rect 20533 19873 20545 19907
rect 20579 19904 20591 19907
rect 22204 19904 22232 20012
rect 26878 20000 26884 20012
rect 26936 20000 26942 20052
rect 27706 19972 27712 19984
rect 25792 19944 27712 19972
rect 25792 19904 25820 19944
rect 27706 19932 27712 19944
rect 27764 19932 27770 19984
rect 27430 19904 27436 19916
rect 20579 19876 22232 19904
rect 22296 19876 25820 19904
rect 27391 19876 27436 19904
rect 20579 19873 20591 19876
rect 20533 19867 20591 19873
rect 6086 19768 6092 19780
rect 5644 19740 6092 19768
rect 6086 19728 6092 19740
rect 6144 19768 6150 19780
rect 6181 19771 6239 19777
rect 6181 19768 6193 19771
rect 6144 19740 6193 19768
rect 6144 19728 6150 19740
rect 6181 19737 6193 19740
rect 6227 19737 6239 19771
rect 6181 19731 6239 19737
rect 6914 19728 6920 19780
rect 6972 19728 6978 19780
rect 7742 19768 7748 19780
rect 7484 19740 7748 19768
rect 4154 19660 4160 19712
rect 4212 19700 4218 19712
rect 7484 19700 7512 19740
rect 7742 19728 7748 19740
rect 7800 19728 7806 19780
rect 9582 19768 9588 19780
rect 9543 19740 9588 19768
rect 9582 19728 9588 19740
rect 9640 19728 9646 19780
rect 10962 19728 10968 19780
rect 11020 19768 11026 19780
rect 11885 19771 11943 19777
rect 11020 19740 11284 19768
rect 11020 19728 11026 19740
rect 7650 19700 7656 19712
rect 4212 19672 7512 19700
rect 7611 19672 7656 19700
rect 4212 19660 4218 19672
rect 7650 19660 7656 19672
rect 7708 19700 7714 19712
rect 8110 19700 8116 19712
rect 7708 19672 8116 19700
rect 7708 19660 7714 19672
rect 8110 19660 8116 19672
rect 8168 19660 8174 19712
rect 11054 19700 11060 19712
rect 11015 19672 11060 19700
rect 11054 19660 11060 19672
rect 11112 19660 11118 19712
rect 11256 19700 11284 19740
rect 11885 19737 11897 19771
rect 11931 19768 11943 19771
rect 12158 19768 12164 19780
rect 11931 19740 12164 19768
rect 11931 19737 11943 19740
rect 11885 19731 11943 19737
rect 12158 19728 12164 19740
rect 12216 19728 12222 19780
rect 13372 19700 13400 19867
rect 15102 19836 15108 19848
rect 15063 19808 15108 19836
rect 15102 19796 15108 19808
rect 15160 19796 15166 19848
rect 22097 19839 22155 19845
rect 22097 19836 22109 19839
rect 21376 19808 22109 19836
rect 15378 19768 15384 19780
rect 15339 19740 15384 19768
rect 15378 19728 15384 19740
rect 15436 19728 15442 19780
rect 16758 19768 16764 19780
rect 16606 19740 16764 19768
rect 16758 19728 16764 19740
rect 16816 19728 16822 19780
rect 17954 19728 17960 19780
rect 18012 19768 18018 19780
rect 20625 19771 20683 19777
rect 20625 19768 20637 19771
rect 18012 19740 20637 19768
rect 18012 19728 18018 19740
rect 20625 19737 20637 19740
rect 20671 19737 20683 19771
rect 20625 19731 20683 19737
rect 16850 19700 16856 19712
rect 11256 19672 13400 19700
rect 16811 19672 16856 19700
rect 16850 19660 16856 19672
rect 16908 19660 16914 19712
rect 20346 19660 20352 19712
rect 20404 19700 20410 19712
rect 21376 19700 21404 19808
rect 22097 19805 22109 19808
rect 22143 19836 22155 19839
rect 22296 19836 22324 19876
rect 27430 19864 27436 19876
rect 27488 19864 27494 19916
rect 27798 19904 27804 19916
rect 27759 19876 27804 19904
rect 27798 19864 27804 19876
rect 27856 19864 27862 19916
rect 31110 19864 31116 19916
rect 31168 19904 31174 19916
rect 31297 19907 31355 19913
rect 31297 19904 31309 19907
rect 31168 19876 31309 19904
rect 31168 19864 31174 19876
rect 31297 19873 31309 19876
rect 31343 19873 31355 19907
rect 31297 19867 31355 19873
rect 23198 19836 23204 19848
rect 22143 19808 22324 19836
rect 22388 19808 23204 19836
rect 22143 19805 22155 19808
rect 22097 19799 22155 19805
rect 21545 19771 21603 19777
rect 21545 19737 21557 19771
rect 21591 19768 21603 19771
rect 22388 19768 22416 19808
rect 23198 19796 23204 19808
rect 23256 19796 23262 19848
rect 22554 19768 22560 19780
rect 21591 19740 22416 19768
rect 22515 19740 22560 19768
rect 21591 19737 21603 19740
rect 21545 19731 21603 19737
rect 22554 19728 22560 19740
rect 22612 19728 22618 19780
rect 27522 19728 27528 19780
rect 27580 19768 27586 19780
rect 27580 19740 27625 19768
rect 27580 19728 27586 19740
rect 20404 19672 21404 19700
rect 20404 19660 20410 19672
rect 21634 19660 21640 19712
rect 21692 19700 21698 19712
rect 23566 19700 23572 19712
rect 21692 19672 23572 19700
rect 21692 19660 21698 19672
rect 23566 19660 23572 19672
rect 23624 19660 23630 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 3234 19456 3240 19508
rect 3292 19496 3298 19508
rect 3329 19499 3387 19505
rect 3329 19496 3341 19499
rect 3292 19468 3341 19496
rect 3292 19456 3298 19468
rect 3329 19465 3341 19468
rect 3375 19465 3387 19499
rect 3329 19459 3387 19465
rect 4246 19456 4252 19508
rect 4304 19496 4310 19508
rect 5350 19496 5356 19508
rect 4304 19468 5356 19496
rect 4304 19456 4310 19468
rect 5350 19456 5356 19468
rect 5408 19456 5414 19508
rect 8202 19496 8208 19508
rect 7208 19468 8208 19496
rect 4154 19428 4160 19440
rect 3082 19400 4160 19428
rect 4154 19388 4160 19400
rect 4212 19388 4218 19440
rect 4798 19428 4804 19440
rect 4264 19400 4804 19428
rect 4062 19320 4068 19372
rect 4120 19360 4126 19372
rect 4264 19369 4292 19400
rect 4798 19388 4804 19400
rect 4856 19388 4862 19440
rect 7208 19428 7236 19468
rect 8202 19456 8208 19468
rect 8260 19456 8266 19508
rect 9582 19456 9588 19508
rect 9640 19496 9646 19508
rect 11149 19499 11207 19505
rect 11149 19496 11161 19499
rect 9640 19468 11161 19496
rect 9640 19456 9646 19468
rect 11149 19465 11161 19468
rect 11195 19496 11207 19499
rect 11514 19496 11520 19508
rect 11195 19468 11520 19496
rect 11195 19465 11207 19468
rect 11149 19459 11207 19465
rect 11514 19456 11520 19468
rect 11572 19456 11578 19508
rect 11698 19456 11704 19508
rect 11756 19496 11762 19508
rect 11793 19499 11851 19505
rect 11793 19496 11805 19499
rect 11756 19468 11805 19496
rect 11756 19456 11762 19468
rect 11793 19465 11805 19468
rect 11839 19465 11851 19499
rect 11793 19459 11851 19465
rect 16758 19456 16764 19508
rect 16816 19496 16822 19508
rect 23661 19499 23719 19505
rect 23661 19496 23673 19499
rect 16816 19468 23673 19496
rect 16816 19456 16822 19468
rect 23661 19465 23673 19468
rect 23707 19465 23719 19499
rect 23661 19459 23719 19465
rect 30929 19499 30987 19505
rect 30929 19465 30941 19499
rect 30975 19496 30987 19499
rect 31662 19496 31668 19508
rect 30975 19468 31668 19496
rect 30975 19465 30987 19468
rect 30929 19459 30987 19465
rect 31662 19456 31668 19468
rect 31720 19456 31726 19508
rect 38102 19496 38108 19508
rect 38063 19468 38108 19496
rect 38102 19456 38108 19468
rect 38160 19456 38166 19508
rect 5750 19400 7236 19428
rect 7374 19388 7380 19440
rect 7432 19388 7438 19440
rect 9677 19431 9735 19437
rect 9677 19397 9689 19431
rect 9723 19428 9735 19431
rect 9766 19428 9772 19440
rect 9723 19400 9772 19428
rect 9723 19397 9735 19400
rect 9677 19391 9735 19397
rect 9766 19388 9772 19400
rect 9824 19388 9830 19440
rect 9950 19388 9956 19440
rect 10008 19428 10014 19440
rect 10008 19400 10166 19428
rect 10008 19388 10014 19400
rect 11054 19388 11060 19440
rect 11112 19428 11118 19440
rect 12342 19428 12348 19440
rect 11112 19400 12348 19428
rect 11112 19388 11118 19400
rect 12342 19388 12348 19400
rect 12400 19388 12406 19440
rect 15102 19428 15108 19440
rect 14568 19400 15108 19428
rect 4249 19363 4307 19369
rect 4249 19360 4261 19363
rect 4120 19332 4261 19360
rect 4120 19320 4126 19332
rect 4249 19329 4261 19332
rect 4295 19329 4307 19363
rect 6546 19360 6552 19372
rect 6507 19332 6552 19360
rect 4249 19323 4307 19329
rect 6546 19320 6552 19332
rect 6604 19320 6610 19372
rect 8110 19320 8116 19372
rect 8168 19360 8174 19372
rect 8168 19332 8524 19360
rect 8168 19320 8174 19332
rect 1578 19292 1584 19304
rect 1539 19264 1584 19292
rect 1578 19252 1584 19264
rect 1636 19252 1642 19304
rect 1857 19295 1915 19301
rect 1857 19261 1869 19295
rect 1903 19292 1915 19295
rect 4154 19292 4160 19304
rect 1903 19264 4160 19292
rect 1903 19261 1915 19264
rect 1857 19255 1915 19261
rect 4154 19252 4160 19264
rect 4212 19252 4218 19304
rect 4525 19295 4583 19301
rect 4525 19261 4537 19295
rect 4571 19292 4583 19295
rect 5718 19292 5724 19304
rect 4571 19264 5724 19292
rect 4571 19261 4583 19264
rect 4525 19255 4583 19261
rect 5718 19252 5724 19264
rect 5776 19252 5782 19304
rect 7190 19252 7196 19304
rect 7248 19292 7254 19304
rect 8496 19292 8524 19332
rect 9122 19320 9128 19372
rect 9180 19360 9186 19372
rect 9401 19363 9459 19369
rect 9401 19360 9413 19363
rect 9180 19332 9413 19360
rect 9180 19320 9186 19332
rect 9401 19329 9413 19332
rect 9447 19329 9459 19363
rect 11701 19363 11759 19369
rect 11701 19360 11713 19363
rect 9401 19323 9459 19329
rect 11072 19332 11713 19360
rect 11072 19304 11100 19332
rect 11701 19329 11713 19332
rect 11747 19360 11759 19363
rect 12250 19360 12256 19372
rect 11747 19332 12256 19360
rect 11747 19329 11759 19332
rect 11701 19323 11759 19329
rect 12250 19320 12256 19332
rect 12308 19320 12314 19372
rect 14568 19369 14596 19400
rect 15102 19388 15108 19400
rect 15160 19388 15166 19440
rect 16482 19428 16488 19440
rect 16054 19400 16488 19428
rect 16482 19388 16488 19400
rect 16540 19388 16546 19440
rect 22186 19428 22192 19440
rect 22147 19400 22192 19428
rect 22186 19388 22192 19400
rect 22244 19388 22250 19440
rect 23014 19388 23020 19440
rect 23072 19428 23078 19440
rect 27890 19428 27896 19440
rect 23072 19400 27896 19428
rect 23072 19388 23078 19400
rect 27890 19388 27896 19400
rect 27948 19388 27954 19440
rect 14553 19363 14611 19369
rect 14553 19329 14565 19363
rect 14599 19329 14611 19363
rect 14553 19323 14611 19329
rect 19889 19363 19947 19369
rect 19889 19329 19901 19363
rect 19935 19360 19947 19363
rect 19978 19360 19984 19372
rect 19935 19332 19984 19360
rect 19935 19329 19947 19332
rect 19889 19323 19947 19329
rect 19978 19320 19984 19332
rect 20036 19320 20042 19372
rect 21910 19320 21916 19372
rect 21968 19320 21974 19372
rect 23566 19360 23572 19372
rect 23527 19332 23572 19360
rect 23566 19320 23572 19332
rect 23624 19320 23630 19372
rect 30834 19360 30840 19372
rect 30795 19332 30840 19360
rect 30834 19320 30840 19332
rect 30892 19320 30898 19372
rect 31846 19320 31852 19372
rect 31904 19360 31910 19372
rect 32585 19363 32643 19369
rect 32585 19360 32597 19363
rect 31904 19332 32597 19360
rect 31904 19320 31910 19332
rect 32585 19329 32597 19332
rect 32631 19329 32643 19363
rect 32585 19323 32643 19329
rect 32677 19363 32735 19369
rect 32677 19329 32689 19363
rect 32723 19360 32735 19363
rect 33318 19360 33324 19372
rect 32723 19332 33324 19360
rect 32723 19329 32735 19332
rect 32677 19323 32735 19329
rect 33318 19320 33324 19332
rect 33376 19320 33382 19372
rect 38286 19360 38292 19372
rect 38247 19332 38292 19360
rect 38286 19320 38292 19332
rect 38344 19320 38350 19372
rect 10134 19292 10140 19304
rect 7248 19264 7880 19292
rect 8496 19264 10140 19292
rect 7248 19252 7254 19264
rect 7852 19224 7880 19264
rect 10134 19252 10140 19264
rect 10192 19252 10198 19304
rect 11054 19252 11060 19304
rect 11112 19252 11118 19304
rect 14829 19295 14887 19301
rect 14829 19261 14841 19295
rect 14875 19292 14887 19295
rect 17586 19292 17592 19304
rect 14875 19264 17592 19292
rect 14875 19261 14887 19264
rect 14829 19255 14887 19261
rect 17586 19252 17592 19264
rect 17644 19252 17650 19304
rect 21928 19292 21956 19320
rect 22097 19295 22155 19301
rect 22097 19292 22109 19295
rect 21928 19264 22109 19292
rect 22097 19261 22109 19264
rect 22143 19261 22155 19295
rect 22097 19255 22155 19261
rect 22373 19295 22431 19301
rect 22373 19261 22385 19295
rect 22419 19261 22431 19295
rect 22373 19255 22431 19261
rect 7852 19196 8432 19224
rect 4706 19116 4712 19168
rect 4764 19156 4770 19168
rect 5997 19159 6055 19165
rect 5997 19156 6009 19159
rect 4764 19128 6009 19156
rect 4764 19116 4770 19128
rect 5997 19125 6009 19128
rect 6043 19125 6055 19159
rect 5997 19119 6055 19125
rect 6812 19159 6870 19165
rect 6812 19125 6824 19159
rect 6858 19156 6870 19159
rect 7558 19156 7564 19168
rect 6858 19128 7564 19156
rect 6858 19125 6870 19128
rect 6812 19119 6870 19125
rect 7558 19116 7564 19128
rect 7616 19156 7622 19168
rect 8110 19156 8116 19168
rect 7616 19128 8116 19156
rect 7616 19116 7622 19128
rect 8110 19116 8116 19128
rect 8168 19116 8174 19168
rect 8294 19156 8300 19168
rect 8255 19128 8300 19156
rect 8294 19116 8300 19128
rect 8352 19116 8358 19168
rect 8404 19156 8432 19196
rect 16206 19184 16212 19236
rect 16264 19224 16270 19236
rect 19702 19224 19708 19236
rect 16264 19196 19708 19224
rect 16264 19184 16270 19196
rect 19702 19184 19708 19196
rect 19760 19184 19766 19236
rect 20714 19184 20720 19236
rect 20772 19224 20778 19236
rect 22388 19224 22416 19255
rect 20772 19196 22416 19224
rect 20772 19184 20778 19196
rect 22066 19168 22094 19196
rect 14458 19156 14464 19168
rect 8404 19128 14464 19156
rect 14458 19116 14464 19128
rect 14516 19116 14522 19168
rect 16301 19159 16359 19165
rect 16301 19125 16313 19159
rect 16347 19156 16359 19159
rect 16390 19156 16396 19168
rect 16347 19128 16396 19156
rect 16347 19125 16359 19128
rect 16301 19119 16359 19125
rect 16390 19116 16396 19128
rect 16448 19116 16454 19168
rect 19518 19116 19524 19168
rect 19576 19156 19582 19168
rect 19981 19159 20039 19165
rect 19981 19156 19993 19159
rect 19576 19128 19993 19156
rect 19576 19116 19582 19128
rect 19981 19125 19993 19128
rect 20027 19156 20039 19159
rect 20254 19156 20260 19168
rect 20027 19128 20260 19156
rect 20027 19125 20039 19128
rect 19981 19119 20039 19125
rect 20254 19116 20260 19128
rect 20312 19116 20318 19168
rect 22066 19128 22100 19168
rect 22094 19116 22100 19128
rect 22152 19116 22158 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 1302 18912 1308 18964
rect 1360 18952 1366 18964
rect 6181 18955 6239 18961
rect 6181 18952 6193 18955
rect 1360 18924 6193 18952
rect 1360 18912 1366 18924
rect 6181 18921 6193 18924
rect 6227 18921 6239 18955
rect 6181 18915 6239 18921
rect 6638 18912 6644 18964
rect 6696 18952 6702 18964
rect 10318 18952 10324 18964
rect 6696 18924 10324 18952
rect 6696 18912 6702 18924
rect 10318 18912 10324 18924
rect 10376 18912 10382 18964
rect 18046 18952 18052 18964
rect 10888 18924 18052 18952
rect 4430 18884 4436 18896
rect 2976 18856 4436 18884
rect 1857 18819 1915 18825
rect 1857 18785 1869 18819
rect 1903 18816 1915 18819
rect 2976 18816 3004 18856
rect 4430 18844 4436 18856
rect 4488 18844 4494 18896
rect 5718 18844 5724 18896
rect 5776 18884 5782 18896
rect 6454 18884 6460 18896
rect 5776 18856 6460 18884
rect 5776 18844 5782 18856
rect 6454 18844 6460 18856
rect 6512 18884 6518 18896
rect 6512 18856 6960 18884
rect 6512 18844 6518 18856
rect 1903 18788 3004 18816
rect 1903 18785 1915 18788
rect 1857 18779 1915 18785
rect 3050 18776 3056 18828
rect 3108 18816 3114 18828
rect 3329 18819 3387 18825
rect 3329 18816 3341 18819
rect 3108 18788 3341 18816
rect 3108 18776 3114 18788
rect 3329 18785 3341 18788
rect 3375 18816 3387 18819
rect 4798 18816 4804 18828
rect 3375 18788 4804 18816
rect 3375 18785 3387 18788
rect 3329 18779 3387 18785
rect 4798 18776 4804 18788
rect 4856 18776 4862 18828
rect 6546 18776 6552 18828
rect 6604 18816 6610 18828
rect 6825 18819 6883 18825
rect 6825 18816 6837 18819
rect 6604 18788 6837 18816
rect 6604 18776 6610 18788
rect 6825 18785 6837 18788
rect 6871 18785 6883 18819
rect 6932 18816 6960 18856
rect 8478 18844 8484 18896
rect 8536 18884 8542 18896
rect 8573 18887 8631 18893
rect 8573 18884 8585 18887
rect 8536 18856 8585 18884
rect 8536 18844 8542 18856
rect 8573 18853 8585 18856
rect 8619 18853 8631 18887
rect 8573 18847 8631 18853
rect 8386 18816 8392 18828
rect 6932 18788 8392 18816
rect 6825 18779 6883 18785
rect 8386 18776 8392 18788
rect 8444 18776 8450 18828
rect 8588 18816 8616 18847
rect 10888 18816 10916 18924
rect 18046 18912 18052 18924
rect 18104 18912 18110 18964
rect 19978 18912 19984 18964
rect 20036 18952 20042 18964
rect 20036 18924 22094 18952
rect 20036 18912 20042 18924
rect 17678 18844 17684 18896
rect 17736 18884 17742 18896
rect 21634 18884 21640 18896
rect 17736 18856 21640 18884
rect 17736 18844 17742 18856
rect 21634 18844 21640 18856
rect 21692 18844 21698 18896
rect 22066 18884 22094 18924
rect 22186 18912 22192 18964
rect 22244 18952 22250 18964
rect 22281 18955 22339 18961
rect 22281 18952 22293 18955
rect 22244 18924 22293 18952
rect 22244 18912 22250 18924
rect 22281 18921 22293 18924
rect 22327 18921 22339 18955
rect 22281 18915 22339 18921
rect 23017 18887 23075 18893
rect 23017 18884 23029 18887
rect 22066 18856 23029 18884
rect 23017 18853 23029 18856
rect 23063 18853 23075 18887
rect 23017 18847 23075 18853
rect 11974 18816 11980 18828
rect 8588 18788 10916 18816
rect 11935 18788 11980 18816
rect 11974 18776 11980 18788
rect 12032 18776 12038 18828
rect 12253 18819 12311 18825
rect 12253 18785 12265 18819
rect 12299 18816 12311 18819
rect 12299 18788 14412 18816
rect 12299 18785 12311 18788
rect 12253 18779 12311 18785
rect 1578 18748 1584 18760
rect 1539 18720 1584 18748
rect 1578 18708 1584 18720
rect 1636 18708 1642 18760
rect 4154 18708 4160 18760
rect 4212 18748 4218 18760
rect 4433 18751 4491 18757
rect 4433 18748 4445 18751
rect 4212 18720 4445 18748
rect 4212 18708 4218 18720
rect 4433 18717 4445 18720
rect 4479 18717 4491 18751
rect 4433 18711 4491 18717
rect 8754 18708 8760 18760
rect 8812 18748 8818 18760
rect 9306 18748 9312 18760
rect 8812 18720 9312 18748
rect 8812 18708 8818 18720
rect 9306 18708 9312 18720
rect 9364 18748 9370 18760
rect 9585 18751 9643 18757
rect 9585 18748 9597 18751
rect 9364 18720 9597 18748
rect 9364 18708 9370 18720
rect 9585 18717 9597 18720
rect 9631 18717 9643 18751
rect 14384 18748 14412 18788
rect 14458 18776 14464 18828
rect 14516 18816 14522 18828
rect 14516 18788 22094 18816
rect 14516 18776 14522 18788
rect 14384 18720 14504 18748
rect 9585 18711 9643 18717
rect 3082 18652 4660 18680
rect 4632 18612 4660 18652
rect 4706 18640 4712 18692
rect 4764 18680 4770 18692
rect 4764 18652 4809 18680
rect 4764 18640 4770 18652
rect 5718 18640 5724 18692
rect 5776 18640 5782 18692
rect 7101 18683 7159 18689
rect 7101 18649 7113 18683
rect 7147 18680 7159 18683
rect 7147 18652 7328 18680
rect 7147 18649 7159 18652
rect 7101 18643 7159 18649
rect 7300 18624 7328 18652
rect 7558 18640 7564 18692
rect 7616 18640 7622 18692
rect 9398 18680 9404 18692
rect 8496 18652 9404 18680
rect 6638 18612 6644 18624
rect 4632 18584 6644 18612
rect 6638 18572 6644 18584
rect 6696 18572 6702 18624
rect 7282 18572 7288 18624
rect 7340 18612 7346 18624
rect 8496 18612 8524 18652
rect 9398 18640 9404 18652
rect 9456 18640 9462 18692
rect 9858 18680 9864 18692
rect 9819 18652 9864 18680
rect 9858 18640 9864 18652
rect 9916 18640 9922 18692
rect 14366 18680 14372 18692
rect 9968 18652 10350 18680
rect 13478 18652 14372 18680
rect 7340 18584 8524 18612
rect 7340 18572 7346 18584
rect 8846 18572 8852 18624
rect 8904 18612 8910 18624
rect 9968 18612 9996 18652
rect 14366 18640 14372 18652
rect 14424 18640 14430 18692
rect 14476 18680 14504 18720
rect 15102 18708 15108 18760
rect 15160 18748 15166 18760
rect 15381 18751 15439 18757
rect 15381 18748 15393 18751
rect 15160 18720 15393 18748
rect 15160 18708 15166 18720
rect 15381 18717 15393 18720
rect 15427 18717 15439 18751
rect 15381 18711 15439 18717
rect 17405 18751 17463 18757
rect 17405 18717 17417 18751
rect 17451 18748 17463 18751
rect 17494 18748 17500 18760
rect 17451 18720 17500 18748
rect 17451 18717 17463 18720
rect 17405 18711 17463 18717
rect 17494 18708 17500 18720
rect 17552 18708 17558 18760
rect 22066 18748 22094 18788
rect 22189 18751 22247 18757
rect 22189 18748 22201 18751
rect 22066 18720 22201 18748
rect 22189 18717 22201 18720
rect 22235 18717 22247 18751
rect 22922 18748 22928 18760
rect 22883 18720 22928 18748
rect 22189 18711 22247 18717
rect 22922 18708 22928 18720
rect 22980 18748 22986 18760
rect 23382 18748 23388 18760
rect 22980 18720 23388 18748
rect 22980 18708 22986 18720
rect 23382 18708 23388 18720
rect 23440 18708 23446 18760
rect 27246 18708 27252 18760
rect 27304 18748 27310 18760
rect 30285 18751 30343 18757
rect 30285 18748 30297 18751
rect 27304 18720 30297 18748
rect 27304 18708 27310 18720
rect 30285 18717 30297 18720
rect 30331 18717 30343 18751
rect 30285 18711 30343 18717
rect 15562 18680 15568 18692
rect 14476 18652 15568 18680
rect 15562 18640 15568 18652
rect 15620 18640 15626 18692
rect 15657 18683 15715 18689
rect 15657 18649 15669 18683
rect 15703 18649 15715 18683
rect 17678 18680 17684 18692
rect 16882 18652 17684 18680
rect 15657 18643 15715 18649
rect 11330 18612 11336 18624
rect 8904 18584 9996 18612
rect 11291 18584 11336 18612
rect 8904 18572 8910 18584
rect 11330 18572 11336 18584
rect 11388 18572 11394 18624
rect 13170 18572 13176 18624
rect 13228 18612 13234 18624
rect 13725 18615 13783 18621
rect 13725 18612 13737 18615
rect 13228 18584 13737 18612
rect 13228 18572 13234 18584
rect 13725 18581 13737 18584
rect 13771 18581 13783 18615
rect 15672 18612 15700 18643
rect 17678 18640 17684 18652
rect 17736 18640 17742 18692
rect 19518 18680 19524 18692
rect 19479 18652 19524 18680
rect 19518 18640 19524 18652
rect 19576 18640 19582 18692
rect 19613 18683 19671 18689
rect 19613 18649 19625 18683
rect 19659 18649 19671 18683
rect 19613 18643 19671 18649
rect 16390 18612 16396 18624
rect 15672 18584 16396 18612
rect 13725 18575 13783 18581
rect 16390 18572 16396 18584
rect 16448 18572 16454 18624
rect 19334 18572 19340 18624
rect 19392 18612 19398 18624
rect 19628 18612 19656 18643
rect 20070 18640 20076 18692
rect 20128 18680 20134 18692
rect 20530 18680 20536 18692
rect 20128 18652 20536 18680
rect 20128 18640 20134 18652
rect 20530 18640 20536 18652
rect 20588 18640 20594 18692
rect 21082 18680 21088 18692
rect 21043 18652 21088 18680
rect 21082 18640 21088 18652
rect 21140 18640 21146 18692
rect 19392 18584 19656 18612
rect 19392 18572 19398 18584
rect 19702 18572 19708 18624
rect 19760 18612 19766 18624
rect 21177 18615 21235 18621
rect 21177 18612 21189 18615
rect 19760 18584 21189 18612
rect 19760 18572 19766 18584
rect 21177 18581 21189 18584
rect 21223 18581 21235 18615
rect 30374 18612 30380 18624
rect 30335 18584 30380 18612
rect 21177 18575 21235 18581
rect 30374 18572 30380 18584
rect 30432 18572 30438 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 3694 18368 3700 18420
rect 3752 18408 3758 18420
rect 4706 18408 4712 18420
rect 3752 18380 4712 18408
rect 3752 18368 3758 18380
rect 4706 18368 4712 18380
rect 4764 18368 4770 18420
rect 7190 18368 7196 18420
rect 7248 18408 7254 18420
rect 7248 18380 8892 18408
rect 7248 18368 7254 18380
rect 1670 18340 1676 18352
rect 1631 18312 1676 18340
rect 1670 18300 1676 18312
rect 1728 18300 1734 18352
rect 3326 18300 3332 18352
rect 3384 18300 3390 18352
rect 4430 18300 4436 18352
rect 4488 18340 4494 18352
rect 6546 18340 6552 18352
rect 4488 18312 6552 18340
rect 4488 18300 4494 18312
rect 6546 18300 6552 18312
rect 6604 18300 6610 18352
rect 8754 18340 8760 18352
rect 8220 18312 8760 18340
rect 7558 18272 7564 18284
rect 4080 18244 7564 18272
rect 2590 18204 2596 18216
rect 2551 18176 2596 18204
rect 2590 18164 2596 18176
rect 2648 18164 2654 18216
rect 2866 18204 2872 18216
rect 2827 18176 2872 18204
rect 2866 18164 2872 18176
rect 2924 18164 2930 18216
rect 3418 18164 3424 18216
rect 3476 18204 3482 18216
rect 4080 18204 4108 18244
rect 7558 18232 7564 18244
rect 7616 18232 7622 18284
rect 7834 18232 7840 18284
rect 7892 18232 7898 18284
rect 8220 18281 8248 18312
rect 8754 18300 8760 18312
rect 8812 18300 8818 18352
rect 8864 18340 8892 18380
rect 9398 18368 9404 18420
rect 9456 18408 9462 18420
rect 9953 18411 10011 18417
rect 9953 18408 9965 18411
rect 9456 18380 9965 18408
rect 9456 18368 9462 18380
rect 9953 18377 9965 18380
rect 9999 18377 10011 18411
rect 9953 18371 10011 18377
rect 11330 18368 11336 18420
rect 11388 18408 11394 18420
rect 25682 18408 25688 18420
rect 11388 18380 25688 18408
rect 11388 18368 11394 18380
rect 25682 18368 25688 18380
rect 25740 18368 25746 18420
rect 29454 18368 29460 18420
rect 29512 18408 29518 18420
rect 29733 18411 29791 18417
rect 29733 18408 29745 18411
rect 29512 18380 29745 18408
rect 29512 18368 29518 18380
rect 29733 18377 29745 18380
rect 29779 18377 29791 18411
rect 29733 18371 29791 18377
rect 33137 18411 33195 18417
rect 33137 18377 33149 18411
rect 33183 18408 33195 18411
rect 33183 18380 35894 18408
rect 33183 18377 33195 18380
rect 33137 18371 33195 18377
rect 8864 18312 8970 18340
rect 10318 18300 10324 18352
rect 10376 18340 10382 18352
rect 12802 18340 12808 18352
rect 10376 18312 12808 18340
rect 10376 18300 10382 18312
rect 12802 18300 12808 18312
rect 12860 18300 12866 18352
rect 15470 18340 15476 18352
rect 14398 18312 15476 18340
rect 15470 18300 15476 18312
rect 15528 18300 15534 18352
rect 16758 18300 16764 18352
rect 16816 18340 16822 18352
rect 16816 18312 17618 18340
rect 16816 18300 16822 18312
rect 18690 18300 18696 18352
rect 18748 18340 18754 18352
rect 19886 18340 19892 18352
rect 18748 18312 19892 18340
rect 18748 18300 18754 18312
rect 19886 18300 19892 18312
rect 19944 18300 19950 18352
rect 19981 18343 20039 18349
rect 19981 18309 19993 18343
rect 20027 18340 20039 18343
rect 20990 18340 20996 18352
rect 20027 18312 20996 18340
rect 20027 18309 20039 18312
rect 19981 18303 20039 18309
rect 20990 18300 20996 18312
rect 21048 18300 21054 18352
rect 23842 18340 23848 18352
rect 23803 18312 23848 18340
rect 23842 18300 23848 18312
rect 23900 18300 23906 18352
rect 8205 18275 8263 18281
rect 8205 18241 8217 18275
rect 8251 18241 8263 18275
rect 8205 18235 8263 18241
rect 15102 18232 15108 18284
rect 15160 18272 15166 18284
rect 16853 18275 16911 18281
rect 16853 18272 16865 18275
rect 15160 18244 16865 18272
rect 15160 18232 15166 18244
rect 16853 18241 16865 18244
rect 16899 18241 16911 18275
rect 16853 18235 16911 18241
rect 29641 18275 29699 18281
rect 29641 18241 29653 18275
rect 29687 18272 29699 18275
rect 33318 18272 33324 18284
rect 29687 18244 30236 18272
rect 33279 18244 33324 18272
rect 29687 18241 29699 18244
rect 29641 18235 29699 18241
rect 3476 18176 4108 18204
rect 4617 18207 4675 18213
rect 3476 18164 3482 18176
rect 4617 18173 4629 18207
rect 4663 18204 4675 18207
rect 4706 18204 4712 18216
rect 4663 18176 4712 18204
rect 4663 18173 4675 18176
rect 4617 18167 4675 18173
rect 4706 18164 4712 18176
rect 4764 18204 4770 18216
rect 7852 18204 7880 18232
rect 30208 18216 30236 18244
rect 33318 18232 33324 18244
rect 33376 18232 33382 18284
rect 35866 18272 35894 18380
rect 38013 18275 38071 18281
rect 38013 18272 38025 18275
rect 35866 18244 38025 18272
rect 38013 18241 38025 18244
rect 38059 18241 38071 18275
rect 38013 18235 38071 18241
rect 4764 18176 7880 18204
rect 8481 18207 8539 18213
rect 4764 18164 4770 18176
rect 8481 18173 8493 18207
rect 8527 18204 8539 18207
rect 11330 18204 11336 18216
rect 8527 18176 11336 18204
rect 8527 18173 8539 18176
rect 8481 18167 8539 18173
rect 11330 18164 11336 18176
rect 11388 18164 11394 18216
rect 12894 18204 12900 18216
rect 12855 18176 12900 18204
rect 12894 18164 12900 18176
rect 12952 18164 12958 18216
rect 13170 18204 13176 18216
rect 13131 18176 13176 18204
rect 13170 18164 13176 18176
rect 13228 18164 13234 18216
rect 14921 18207 14979 18213
rect 14921 18173 14933 18207
rect 14967 18204 14979 18207
rect 15378 18204 15384 18216
rect 14967 18176 15384 18204
rect 14967 18173 14979 18176
rect 14921 18167 14979 18173
rect 15378 18164 15384 18176
rect 15436 18164 15442 18216
rect 15562 18164 15568 18216
rect 15620 18204 15626 18216
rect 16206 18204 16212 18216
rect 15620 18176 16212 18204
rect 15620 18164 15626 18176
rect 16206 18164 16212 18176
rect 16264 18164 16270 18216
rect 17126 18204 17132 18216
rect 17039 18176 17132 18204
rect 17126 18164 17132 18176
rect 17184 18204 17190 18216
rect 17494 18204 17500 18216
rect 17184 18176 17500 18204
rect 17184 18164 17190 18176
rect 17494 18164 17500 18176
rect 17552 18164 17558 18216
rect 18138 18164 18144 18216
rect 18196 18204 18202 18216
rect 18598 18204 18604 18216
rect 18196 18176 18604 18204
rect 18196 18164 18202 18176
rect 18598 18164 18604 18176
rect 18656 18164 18662 18216
rect 20257 18207 20315 18213
rect 20257 18173 20269 18207
rect 20303 18173 20315 18207
rect 23750 18204 23756 18216
rect 23711 18176 23756 18204
rect 20257 18167 20315 18173
rect 5350 18096 5356 18148
rect 5408 18136 5414 18148
rect 7558 18136 7564 18148
rect 5408 18108 7564 18136
rect 5408 18096 5414 18108
rect 7558 18096 7564 18108
rect 7616 18096 7622 18148
rect 19886 18136 19892 18148
rect 9508 18108 12434 18136
rect 1765 18071 1823 18077
rect 1765 18037 1777 18071
rect 1811 18068 1823 18071
rect 9508 18068 9536 18108
rect 1811 18040 9536 18068
rect 12406 18068 12434 18108
rect 18156 18108 19892 18136
rect 18156 18068 18184 18108
rect 19886 18096 19892 18108
rect 19944 18096 19950 18148
rect 12406 18040 18184 18068
rect 1811 18037 1823 18040
rect 1765 18031 1823 18037
rect 19150 18028 19156 18080
rect 19208 18068 19214 18080
rect 20272 18068 20300 18167
rect 23750 18164 23756 18176
rect 23808 18164 23814 18216
rect 24029 18207 24087 18213
rect 24029 18173 24041 18207
rect 24075 18173 24087 18207
rect 24029 18167 24087 18173
rect 21450 18096 21456 18148
rect 21508 18136 21514 18148
rect 22002 18136 22008 18148
rect 21508 18108 22008 18136
rect 21508 18096 21514 18108
rect 22002 18096 22008 18108
rect 22060 18136 22066 18148
rect 24044 18136 24072 18167
rect 30190 18164 30196 18216
rect 30248 18204 30254 18216
rect 37918 18204 37924 18216
rect 30248 18176 37924 18204
rect 30248 18164 30254 18176
rect 37918 18164 37924 18176
rect 37976 18164 37982 18216
rect 22060 18108 24072 18136
rect 22060 18096 22066 18108
rect 38194 18068 38200 18080
rect 19208 18040 20300 18068
rect 38155 18040 38200 18068
rect 19208 18028 19214 18040
rect 38194 18028 38200 18040
rect 38252 18028 38258 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 9214 17864 9220 17876
rect 9175 17836 9220 17864
rect 9214 17824 9220 17836
rect 9272 17824 9278 17876
rect 10321 17867 10379 17873
rect 10321 17833 10333 17867
rect 10367 17864 10379 17867
rect 10410 17864 10416 17876
rect 10367 17836 10416 17864
rect 10367 17833 10379 17836
rect 10321 17827 10379 17833
rect 10410 17824 10416 17836
rect 10468 17824 10474 17876
rect 11504 17867 11562 17873
rect 11504 17833 11516 17867
rect 11550 17864 11562 17867
rect 15930 17864 15936 17876
rect 11550 17836 15936 17864
rect 11550 17833 11562 17836
rect 11504 17827 11562 17833
rect 15930 17824 15936 17836
rect 15988 17824 15994 17876
rect 16666 17824 16672 17876
rect 16724 17864 16730 17876
rect 17862 17864 17868 17876
rect 16724 17836 17868 17864
rect 16724 17824 16730 17836
rect 17862 17824 17868 17836
rect 17920 17824 17926 17876
rect 17972 17836 20852 17864
rect 17678 17756 17684 17808
rect 17736 17796 17742 17808
rect 17972 17796 18000 17836
rect 19886 17796 19892 17808
rect 17736 17768 18000 17796
rect 18064 17768 19892 17796
rect 17736 17756 17742 17768
rect 1578 17728 1584 17740
rect 1491 17700 1584 17728
rect 1578 17688 1584 17700
rect 1636 17728 1642 17740
rect 2590 17728 2596 17740
rect 1636 17700 2596 17728
rect 1636 17688 1642 17700
rect 2590 17688 2596 17700
rect 2648 17728 2654 17740
rect 4062 17728 4068 17740
rect 2648 17700 4068 17728
rect 2648 17688 2654 17700
rect 4062 17688 4068 17700
rect 4120 17728 4126 17740
rect 6089 17731 6147 17737
rect 6089 17728 6101 17731
rect 4120 17700 6101 17728
rect 4120 17688 4126 17700
rect 6089 17697 6101 17700
rect 6135 17697 6147 17731
rect 6089 17691 6147 17697
rect 11241 17731 11299 17737
rect 11241 17697 11253 17731
rect 11287 17728 11299 17731
rect 12894 17728 12900 17740
rect 11287 17700 12900 17728
rect 11287 17697 11299 17700
rect 11241 17691 11299 17697
rect 12894 17688 12900 17700
rect 12952 17728 12958 17740
rect 15102 17728 15108 17740
rect 12952 17700 15108 17728
rect 12952 17688 12958 17700
rect 15102 17688 15108 17700
rect 15160 17688 15166 17740
rect 15381 17731 15439 17737
rect 15381 17697 15393 17731
rect 15427 17728 15439 17731
rect 16850 17728 16856 17740
rect 15427 17700 16856 17728
rect 15427 17697 15439 17700
rect 15381 17691 15439 17697
rect 16850 17688 16856 17700
rect 16908 17728 16914 17740
rect 18064 17728 18092 17768
rect 19886 17756 19892 17768
rect 19944 17756 19950 17808
rect 16908 17700 18092 17728
rect 19797 17731 19855 17737
rect 16908 17688 16914 17700
rect 19797 17697 19809 17731
rect 19843 17728 19855 17731
rect 19978 17728 19984 17740
rect 19843 17700 19984 17728
rect 19843 17697 19855 17700
rect 19797 17691 19855 17697
rect 19978 17688 19984 17700
rect 20036 17688 20042 17740
rect 20824 17737 20852 17836
rect 23750 17756 23756 17808
rect 23808 17796 23814 17808
rect 27522 17796 27528 17808
rect 23808 17768 27528 17796
rect 23808 17756 23814 17768
rect 27522 17756 27528 17768
rect 27580 17756 27586 17808
rect 27798 17756 27804 17808
rect 27856 17756 27862 17808
rect 20809 17731 20867 17737
rect 20809 17697 20821 17731
rect 20855 17728 20867 17731
rect 27816 17728 27844 17756
rect 20855 17700 27844 17728
rect 20855 17697 20867 17700
rect 20809 17691 20867 17697
rect 9122 17660 9128 17672
rect 9083 17632 9128 17660
rect 9122 17620 9128 17632
rect 9180 17620 9186 17672
rect 10229 17663 10287 17669
rect 10229 17660 10241 17663
rect 9646 17632 10241 17660
rect 1857 17595 1915 17601
rect 1857 17561 1869 17595
rect 1903 17561 1915 17595
rect 5074 17592 5080 17604
rect 3082 17564 5080 17592
rect 1857 17555 1915 17561
rect 1872 17524 1900 17555
rect 5074 17552 5080 17564
rect 5132 17552 5138 17604
rect 6365 17595 6423 17601
rect 6365 17561 6377 17595
rect 6411 17561 6423 17595
rect 6365 17555 6423 17561
rect 3234 17524 3240 17536
rect 1872 17496 3240 17524
rect 3234 17484 3240 17496
rect 3292 17484 3298 17536
rect 3329 17527 3387 17533
rect 3329 17493 3341 17527
rect 3375 17524 3387 17527
rect 3510 17524 3516 17536
rect 3375 17496 3516 17524
rect 3375 17493 3387 17496
rect 3329 17487 3387 17493
rect 3510 17484 3516 17496
rect 3568 17524 3574 17536
rect 6380 17524 6408 17555
rect 7006 17552 7012 17604
rect 7064 17552 7070 17604
rect 8110 17552 8116 17604
rect 8168 17592 8174 17604
rect 9646 17592 9674 17632
rect 10229 17629 10241 17632
rect 10275 17629 10287 17663
rect 21542 17660 21548 17672
rect 21503 17632 21548 17660
rect 10229 17623 10287 17629
rect 21542 17620 21548 17632
rect 21600 17620 21606 17672
rect 24578 17660 24584 17672
rect 24539 17632 24584 17660
rect 24578 17620 24584 17632
rect 24636 17660 24642 17672
rect 25501 17663 25559 17669
rect 25501 17660 25513 17663
rect 24636 17632 25513 17660
rect 24636 17620 24642 17632
rect 25501 17629 25513 17632
rect 25547 17629 25559 17663
rect 25501 17623 25559 17629
rect 26329 17663 26387 17669
rect 26329 17629 26341 17663
rect 26375 17629 26387 17663
rect 26329 17623 26387 17629
rect 8168 17564 9674 17592
rect 8168 17552 8174 17564
rect 12526 17552 12532 17604
rect 12584 17552 12590 17604
rect 13998 17592 14004 17604
rect 12820 17564 14004 17592
rect 3568 17496 6408 17524
rect 7837 17527 7895 17533
rect 3568 17484 3574 17496
rect 7837 17493 7849 17527
rect 7883 17524 7895 17527
rect 9858 17524 9864 17536
rect 7883 17496 9864 17524
rect 7883 17493 7895 17496
rect 7837 17487 7895 17493
rect 9858 17484 9864 17496
rect 9916 17524 9922 17536
rect 12820 17524 12848 17564
rect 13998 17552 14004 17564
rect 14056 17552 14062 17604
rect 17034 17592 17040 17604
rect 16606 17564 17040 17592
rect 17034 17552 17040 17564
rect 17092 17552 17098 17604
rect 17129 17595 17187 17601
rect 17129 17561 17141 17595
rect 17175 17592 17187 17595
rect 17586 17592 17592 17604
rect 17175 17564 17592 17592
rect 17175 17561 17187 17564
rect 17129 17555 17187 17561
rect 17586 17552 17592 17564
rect 17644 17552 17650 17604
rect 19610 17592 19616 17604
rect 18340 17564 19616 17592
rect 12986 17524 12992 17536
rect 9916 17496 12848 17524
rect 12947 17496 12992 17524
rect 9916 17484 9922 17496
rect 12986 17484 12992 17496
rect 13044 17484 13050 17536
rect 13354 17484 13360 17536
rect 13412 17524 13418 17536
rect 18340 17524 18368 17564
rect 19610 17552 19616 17564
rect 19668 17552 19674 17604
rect 19886 17552 19892 17604
rect 19944 17592 19950 17604
rect 19944 17564 19989 17592
rect 19944 17552 19950 17564
rect 20438 17552 20444 17604
rect 20496 17592 20502 17604
rect 21560 17592 21588 17620
rect 20496 17564 21588 17592
rect 20496 17552 20502 17564
rect 21634 17552 21640 17604
rect 21692 17592 21698 17604
rect 22278 17592 22284 17604
rect 21692 17564 21737 17592
rect 22239 17564 22284 17592
rect 21692 17552 21698 17564
rect 22278 17552 22284 17564
rect 22336 17552 22342 17604
rect 22370 17552 22376 17604
rect 22428 17592 22434 17604
rect 22428 17564 22473 17592
rect 22428 17552 22434 17564
rect 23198 17552 23204 17604
rect 23256 17592 23262 17604
rect 23293 17595 23351 17601
rect 23293 17592 23305 17595
rect 23256 17564 23305 17592
rect 23256 17552 23262 17564
rect 23293 17561 23305 17564
rect 23339 17561 23351 17595
rect 26344 17592 26372 17623
rect 27154 17620 27160 17672
rect 27212 17660 27218 17672
rect 27801 17663 27859 17669
rect 27801 17660 27813 17663
rect 27212 17632 27813 17660
rect 27212 17620 27218 17632
rect 27801 17629 27813 17632
rect 27847 17629 27859 17663
rect 27801 17623 27859 17629
rect 28258 17620 28264 17672
rect 28316 17660 28322 17672
rect 28997 17663 29055 17669
rect 28997 17660 29009 17663
rect 28316 17632 29009 17660
rect 28316 17620 28322 17632
rect 28997 17629 29009 17632
rect 29043 17660 29055 17663
rect 29362 17660 29368 17672
rect 29043 17632 29368 17660
rect 29043 17629 29055 17632
rect 28997 17623 29055 17629
rect 29362 17620 29368 17632
rect 29420 17620 29426 17672
rect 30190 17660 30196 17672
rect 30151 17632 30196 17660
rect 30190 17620 30196 17632
rect 30248 17620 30254 17672
rect 23293 17555 23351 17561
rect 25332 17564 26372 17592
rect 30377 17595 30435 17601
rect 13412 17496 18368 17524
rect 13412 17484 13418 17496
rect 18414 17484 18420 17536
rect 18472 17524 18478 17536
rect 19702 17524 19708 17536
rect 18472 17496 19708 17524
rect 18472 17484 18478 17496
rect 19702 17484 19708 17496
rect 19760 17484 19766 17536
rect 23474 17484 23480 17536
rect 23532 17524 23538 17536
rect 25332 17533 25360 17564
rect 30377 17561 30389 17595
rect 30423 17592 30435 17595
rect 30558 17592 30564 17604
rect 30423 17564 30564 17592
rect 30423 17561 30435 17564
rect 30377 17555 30435 17561
rect 30558 17552 30564 17564
rect 30616 17552 30622 17604
rect 24673 17527 24731 17533
rect 24673 17524 24685 17527
rect 23532 17496 24685 17524
rect 23532 17484 23538 17496
rect 24673 17493 24685 17496
rect 24719 17493 24731 17527
rect 24673 17487 24731 17493
rect 25317 17527 25375 17533
rect 25317 17493 25329 17527
rect 25363 17493 25375 17527
rect 25317 17487 25375 17493
rect 26145 17527 26203 17533
rect 26145 17493 26157 17527
rect 26191 17524 26203 17527
rect 27246 17524 27252 17536
rect 26191 17496 27252 17524
rect 26191 17493 26203 17496
rect 26145 17487 26203 17493
rect 27246 17484 27252 17496
rect 27304 17484 27310 17536
rect 27893 17527 27951 17533
rect 27893 17493 27905 17527
rect 27939 17524 27951 17527
rect 28074 17524 28080 17536
rect 27939 17496 28080 17524
rect 27939 17493 27951 17496
rect 27893 17487 27951 17493
rect 28074 17484 28080 17496
rect 28132 17484 28138 17536
rect 29089 17527 29147 17533
rect 29089 17493 29101 17527
rect 29135 17524 29147 17527
rect 29914 17524 29920 17536
rect 29135 17496 29920 17524
rect 29135 17493 29147 17496
rect 29089 17487 29147 17493
rect 29914 17484 29920 17496
rect 29972 17484 29978 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 8294 17280 8300 17332
rect 8352 17320 8358 17332
rect 16945 17323 17003 17329
rect 8352 17292 14412 17320
rect 8352 17280 8358 17292
rect 3234 17212 3240 17264
rect 3292 17252 3298 17264
rect 10410 17252 10416 17264
rect 3292 17224 10416 17252
rect 3292 17212 3298 17224
rect 10410 17212 10416 17224
rect 10468 17212 10474 17264
rect 11974 17252 11980 17264
rect 10704 17224 11980 17252
rect 1670 17184 1676 17196
rect 1631 17156 1676 17184
rect 1670 17144 1676 17156
rect 1728 17144 1734 17196
rect 2498 17184 2504 17196
rect 2459 17156 2504 17184
rect 2498 17144 2504 17156
rect 2556 17144 2562 17196
rect 7834 17144 7840 17196
rect 7892 17184 7898 17196
rect 10704 17184 10732 17224
rect 11974 17212 11980 17224
rect 12032 17212 12038 17264
rect 7892 17156 10732 17184
rect 7892 17144 7898 17156
rect 10778 17144 10784 17196
rect 10836 17184 10842 17196
rect 14093 17187 14151 17193
rect 14093 17184 14105 17187
rect 10836 17156 14105 17184
rect 10836 17144 10842 17156
rect 14093 17153 14105 17156
rect 14139 17153 14151 17187
rect 14093 17147 14151 17153
rect 14182 17144 14188 17196
rect 14240 17184 14246 17196
rect 14384 17184 14412 17292
rect 16945 17289 16957 17323
rect 16991 17320 17003 17323
rect 17954 17320 17960 17332
rect 16991 17292 17960 17320
rect 16991 17289 17003 17292
rect 16945 17283 17003 17289
rect 17954 17280 17960 17292
rect 18012 17280 18018 17332
rect 20990 17320 20996 17332
rect 20951 17292 20996 17320
rect 20990 17280 20996 17292
rect 21048 17280 21054 17332
rect 28350 17280 28356 17332
rect 28408 17320 28414 17332
rect 28408 17292 30880 17320
rect 28408 17280 28414 17292
rect 17218 17212 17224 17264
rect 17276 17252 17282 17264
rect 22370 17252 22376 17264
rect 17276 17224 22376 17252
rect 17276 17212 17282 17224
rect 22370 17212 22376 17224
rect 22428 17212 22434 17264
rect 25222 17252 25228 17264
rect 23676 17224 25228 17252
rect 16853 17187 16911 17193
rect 16853 17184 16865 17187
rect 14240 17156 14285 17184
rect 14384 17156 16865 17184
rect 14240 17144 14246 17156
rect 16853 17153 16865 17156
rect 16899 17153 16911 17187
rect 17770 17184 17776 17196
rect 17731 17156 17776 17184
rect 16853 17147 16911 17153
rect 17770 17144 17776 17156
rect 17828 17144 17834 17196
rect 17862 17144 17868 17196
rect 17920 17184 17926 17196
rect 20901 17187 20959 17193
rect 20901 17184 20913 17187
rect 17920 17156 20913 17184
rect 17920 17144 17926 17156
rect 20901 17153 20913 17156
rect 20947 17153 20959 17187
rect 20901 17147 20959 17153
rect 9214 17076 9220 17128
rect 9272 17116 9278 17128
rect 23676 17116 23704 17224
rect 25222 17212 25228 17224
rect 25280 17212 25286 17264
rect 27614 17212 27620 17264
rect 27672 17252 27678 17264
rect 30852 17261 30880 17292
rect 29917 17255 29975 17261
rect 29917 17252 29929 17255
rect 27672 17224 29929 17252
rect 27672 17212 27678 17224
rect 29917 17221 29929 17224
rect 29963 17221 29975 17255
rect 29917 17215 29975 17221
rect 30837 17255 30895 17261
rect 30837 17221 30849 17255
rect 30883 17221 30895 17255
rect 30837 17215 30895 17221
rect 24673 17187 24731 17193
rect 24673 17153 24685 17187
rect 24719 17153 24731 17187
rect 27338 17184 27344 17196
rect 27299 17156 27344 17184
rect 24673 17147 24731 17153
rect 9272 17088 23704 17116
rect 9272 17076 9278 17088
rect 1854 17048 1860 17060
rect 1815 17020 1860 17048
rect 1854 17008 1860 17020
rect 1912 17008 1918 17060
rect 1946 17008 1952 17060
rect 2004 17048 2010 17060
rect 8478 17048 8484 17060
rect 2004 17020 8484 17048
rect 2004 17008 2010 17020
rect 8478 17008 8484 17020
rect 8536 17008 8542 17060
rect 8754 17008 8760 17060
rect 8812 17048 8818 17060
rect 11882 17048 11888 17060
rect 8812 17020 11888 17048
rect 8812 17008 8818 17020
rect 11882 17008 11888 17020
rect 11940 17008 11946 17060
rect 11974 17008 11980 17060
rect 12032 17048 12038 17060
rect 17218 17048 17224 17060
rect 12032 17020 17224 17048
rect 12032 17008 12038 17020
rect 17218 17008 17224 17020
rect 17276 17008 17282 17060
rect 24688 17048 24716 17147
rect 27338 17144 27344 17156
rect 27396 17144 27402 17196
rect 28074 17184 28080 17196
rect 28035 17156 28080 17184
rect 28074 17144 28080 17156
rect 28132 17144 28138 17196
rect 25317 17119 25375 17125
rect 25317 17085 25329 17119
rect 25363 17116 25375 17119
rect 25961 17119 26019 17125
rect 25961 17116 25973 17119
rect 25363 17088 25973 17116
rect 25363 17085 25375 17088
rect 25317 17079 25375 17085
rect 25961 17085 25973 17088
rect 26007 17085 26019 17119
rect 26142 17116 26148 17128
rect 26103 17088 26148 17116
rect 25961 17079 26019 17085
rect 26142 17076 26148 17088
rect 26200 17076 26206 17128
rect 27893 17119 27951 17125
rect 27893 17085 27905 17119
rect 27939 17116 27951 17119
rect 29454 17116 29460 17128
rect 27939 17088 29460 17116
rect 27939 17085 27951 17088
rect 27893 17079 27951 17085
rect 29454 17076 29460 17088
rect 29512 17076 29518 17128
rect 29825 17119 29883 17125
rect 29825 17085 29837 17119
rect 29871 17085 29883 17119
rect 29825 17079 29883 17085
rect 26234 17048 26240 17060
rect 17328 17020 26240 17048
rect 2317 16983 2375 16989
rect 2317 16949 2329 16983
rect 2363 16980 2375 16983
rect 3234 16980 3240 16992
rect 2363 16952 3240 16980
rect 2363 16949 2375 16952
rect 2317 16943 2375 16949
rect 3234 16940 3240 16952
rect 3292 16940 3298 16992
rect 8294 16940 8300 16992
rect 8352 16980 8358 16992
rect 9122 16980 9128 16992
rect 8352 16952 9128 16980
rect 8352 16940 8358 16952
rect 9122 16940 9128 16952
rect 9180 16980 9186 16992
rect 15746 16980 15752 16992
rect 9180 16952 15752 16980
rect 9180 16940 9186 16952
rect 15746 16940 15752 16952
rect 15804 16940 15810 16992
rect 16390 16940 16396 16992
rect 16448 16980 16454 16992
rect 17328 16980 17356 17020
rect 26234 17008 26240 17020
rect 26292 17008 26298 17060
rect 29730 17008 29736 17060
rect 29788 17048 29794 17060
rect 29840 17048 29868 17079
rect 29788 17020 29868 17048
rect 29788 17008 29794 17020
rect 16448 16952 17356 16980
rect 16448 16940 16454 16952
rect 17770 16940 17776 16992
rect 17828 16980 17834 16992
rect 17865 16983 17923 16989
rect 17865 16980 17877 16983
rect 17828 16952 17877 16980
rect 17828 16940 17834 16952
rect 17865 16949 17877 16952
rect 17911 16949 17923 16983
rect 17865 16943 17923 16949
rect 17954 16940 17960 16992
rect 18012 16980 18018 16992
rect 20438 16980 20444 16992
rect 18012 16952 20444 16980
rect 18012 16940 18018 16952
rect 20438 16940 20444 16952
rect 20496 16940 20502 16992
rect 24762 16980 24768 16992
rect 24723 16952 24768 16980
rect 24762 16940 24768 16952
rect 24820 16940 24826 16992
rect 26326 16980 26332 16992
rect 26287 16952 26332 16980
rect 26326 16940 26332 16952
rect 26384 16940 26390 16992
rect 26970 16940 26976 16992
rect 27028 16980 27034 16992
rect 27157 16983 27215 16989
rect 27157 16980 27169 16983
rect 27028 16952 27169 16980
rect 27028 16940 27034 16952
rect 27157 16949 27169 16952
rect 27203 16949 27215 16983
rect 28534 16980 28540 16992
rect 28495 16952 28540 16980
rect 27157 16943 27215 16949
rect 28534 16940 28540 16952
rect 28592 16940 28598 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 2774 16736 2780 16788
rect 2832 16776 2838 16788
rect 3602 16776 3608 16788
rect 2832 16748 3608 16776
rect 2832 16736 2838 16748
rect 3602 16736 3608 16748
rect 3660 16736 3666 16788
rect 8110 16736 8116 16788
rect 8168 16776 8174 16788
rect 8168 16748 14320 16776
rect 8168 16736 8174 16748
rect 14292 16720 14320 16748
rect 17218 16736 17224 16788
rect 17276 16776 17282 16788
rect 27982 16776 27988 16788
rect 17276 16748 27988 16776
rect 17276 16736 17282 16748
rect 27982 16736 27988 16748
rect 28040 16736 28046 16788
rect 2130 16668 2136 16720
rect 2188 16708 2194 16720
rect 2188 16680 2912 16708
rect 2188 16668 2194 16680
rect 1946 16640 1952 16652
rect 1907 16612 1952 16640
rect 1946 16600 1952 16612
rect 2004 16600 2010 16652
rect 2317 16643 2375 16649
rect 2317 16609 2329 16643
rect 2363 16640 2375 16643
rect 2774 16640 2780 16652
rect 2363 16612 2780 16640
rect 2363 16609 2375 16612
rect 2317 16603 2375 16609
rect 2774 16600 2780 16612
rect 2832 16600 2838 16652
rect 2884 16581 2912 16680
rect 8478 16668 8484 16720
rect 8536 16708 8542 16720
rect 9769 16711 9827 16717
rect 9769 16708 9781 16711
rect 8536 16680 9781 16708
rect 8536 16668 8542 16680
rect 9769 16677 9781 16680
rect 9815 16677 9827 16711
rect 13354 16708 13360 16720
rect 9769 16671 9827 16677
rect 9876 16680 13360 16708
rect 8294 16640 8300 16652
rect 6748 16612 8300 16640
rect 2869 16575 2927 16581
rect 2869 16541 2881 16575
rect 2915 16541 2927 16575
rect 2869 16535 2927 16541
rect 4062 16532 4068 16584
rect 4120 16572 4126 16584
rect 4157 16575 4215 16581
rect 4157 16572 4169 16575
rect 4120 16544 4169 16572
rect 4120 16532 4126 16544
rect 4157 16541 4169 16544
rect 4203 16541 4215 16575
rect 4157 16535 4215 16541
rect 5537 16575 5595 16581
rect 5537 16541 5549 16575
rect 5583 16572 5595 16575
rect 6178 16572 6184 16584
rect 5583 16544 6184 16572
rect 5583 16541 5595 16544
rect 5537 16535 5595 16541
rect 6178 16532 6184 16544
rect 6236 16532 6242 16584
rect 6748 16581 6776 16612
rect 7392 16581 7420 16612
rect 8294 16600 8300 16612
rect 8352 16600 8358 16652
rect 8386 16600 8392 16652
rect 8444 16640 8450 16652
rect 9876 16640 9904 16680
rect 13354 16668 13360 16680
rect 13412 16668 13418 16720
rect 13464 16680 14228 16708
rect 11790 16640 11796 16652
rect 8444 16612 9904 16640
rect 10888 16612 11796 16640
rect 8444 16600 8450 16612
rect 6733 16575 6791 16581
rect 6733 16541 6745 16575
rect 6779 16541 6791 16575
rect 6733 16535 6791 16541
rect 7377 16575 7435 16581
rect 7377 16541 7389 16575
rect 7423 16541 7435 16575
rect 7377 16535 7435 16541
rect 7466 16532 7472 16584
rect 7524 16572 7530 16584
rect 8110 16572 8116 16584
rect 7524 16544 7569 16572
rect 8071 16544 8116 16572
rect 7524 16532 7530 16544
rect 8110 16532 8116 16544
rect 8168 16532 8174 16584
rect 10318 16532 10324 16584
rect 10376 16572 10382 16584
rect 10888 16581 10916 16612
rect 11532 16581 11560 16612
rect 11790 16600 11796 16612
rect 11848 16600 11854 16652
rect 11882 16600 11888 16652
rect 11940 16640 11946 16652
rect 13464 16640 13492 16680
rect 13722 16640 13728 16652
rect 11940 16612 13492 16640
rect 13556 16612 13728 16640
rect 11940 16600 11946 16612
rect 12176 16581 12204 16612
rect 10873 16575 10931 16581
rect 10873 16572 10885 16575
rect 10376 16544 10885 16572
rect 10376 16532 10382 16544
rect 10873 16541 10885 16544
rect 10919 16541 10931 16575
rect 10873 16535 10931 16541
rect 11517 16575 11575 16581
rect 11517 16541 11529 16575
rect 11563 16541 11575 16575
rect 11517 16535 11575 16541
rect 12161 16575 12219 16581
rect 12161 16541 12173 16575
rect 12207 16541 12219 16575
rect 12161 16535 12219 16541
rect 12253 16575 12311 16581
rect 12253 16541 12265 16575
rect 12299 16572 12311 16575
rect 12526 16572 12532 16584
rect 12299 16544 12532 16572
rect 12299 16541 12311 16544
rect 12253 16535 12311 16541
rect 12526 16532 12532 16544
rect 12584 16532 12590 16584
rect 13556 16581 13584 16612
rect 13722 16600 13728 16612
rect 13780 16600 13786 16652
rect 14200 16640 14228 16680
rect 14274 16668 14280 16720
rect 14332 16708 14338 16720
rect 19058 16708 19064 16720
rect 14332 16680 19064 16708
rect 14332 16668 14338 16680
rect 19058 16668 19064 16680
rect 19116 16668 19122 16720
rect 20622 16640 20628 16652
rect 14200 16612 20628 16640
rect 20622 16600 20628 16612
rect 20680 16600 20686 16652
rect 21082 16600 21088 16652
rect 21140 16640 21146 16652
rect 21726 16640 21732 16652
rect 21140 16612 21732 16640
rect 21140 16600 21146 16612
rect 13541 16575 13599 16581
rect 13541 16541 13553 16575
rect 13587 16541 13599 16575
rect 14274 16572 14280 16584
rect 14235 16544 14280 16572
rect 13541 16535 13599 16541
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 14366 16532 14372 16584
rect 14424 16572 14430 16584
rect 14424 16544 14469 16572
rect 14424 16532 14430 16544
rect 16298 16532 16304 16584
rect 16356 16572 16362 16584
rect 17494 16572 17500 16584
rect 16356 16544 17500 16572
rect 16356 16532 16362 16544
rect 17494 16532 17500 16544
rect 17552 16532 17558 16584
rect 20073 16575 20131 16581
rect 20073 16541 20085 16575
rect 20119 16572 20131 16575
rect 20438 16572 20444 16584
rect 20119 16544 20444 16572
rect 20119 16541 20131 16544
rect 20073 16535 20131 16541
rect 20438 16532 20444 16544
rect 20496 16532 20502 16584
rect 21192 16581 21220 16612
rect 21726 16600 21732 16612
rect 21784 16600 21790 16652
rect 22370 16640 22376 16652
rect 22331 16612 22376 16640
rect 22370 16600 22376 16612
rect 22428 16600 22434 16652
rect 23566 16640 23572 16652
rect 23492 16612 23572 16640
rect 21177 16575 21235 16581
rect 21177 16541 21189 16575
rect 21223 16541 21235 16575
rect 22554 16572 22560 16584
rect 22515 16544 22560 16572
rect 21177 16535 21235 16541
rect 22554 16532 22560 16544
rect 22612 16532 22618 16584
rect 23492 16581 23520 16612
rect 23566 16600 23572 16612
rect 23624 16600 23630 16652
rect 24486 16600 24492 16652
rect 24544 16640 24550 16652
rect 28994 16640 29000 16652
rect 24544 16612 29000 16640
rect 24544 16600 24550 16612
rect 24596 16581 24624 16612
rect 28994 16600 29000 16612
rect 29052 16600 29058 16652
rect 29914 16640 29920 16652
rect 29875 16612 29920 16640
rect 29914 16600 29920 16612
rect 29972 16600 29978 16652
rect 23477 16575 23535 16581
rect 23477 16541 23489 16575
rect 23523 16541 23535 16575
rect 23477 16535 23535 16541
rect 24581 16575 24639 16581
rect 24581 16541 24593 16575
rect 24627 16541 24639 16575
rect 25406 16572 25412 16584
rect 25367 16544 25412 16572
rect 24581 16535 24639 16541
rect 25406 16532 25412 16544
rect 25464 16532 25470 16584
rect 26234 16572 26240 16584
rect 26195 16544 26240 16572
rect 26234 16532 26240 16544
rect 26292 16532 26298 16584
rect 27801 16575 27859 16581
rect 27801 16541 27813 16575
rect 27847 16572 27859 16575
rect 27890 16572 27896 16584
rect 27847 16544 27896 16572
rect 27847 16541 27859 16544
rect 27801 16535 27859 16541
rect 27890 16532 27896 16544
rect 27948 16532 27954 16584
rect 29730 16572 29736 16584
rect 29691 16544 29736 16572
rect 29730 16532 29736 16544
rect 29788 16532 29794 16584
rect 30377 16575 30435 16581
rect 30377 16541 30389 16575
rect 30423 16572 30435 16575
rect 30466 16572 30472 16584
rect 30423 16544 30472 16572
rect 30423 16541 30435 16544
rect 30377 16535 30435 16541
rect 30466 16532 30472 16544
rect 30524 16532 30530 16584
rect 38010 16572 38016 16584
rect 37971 16544 38016 16572
rect 38010 16532 38016 16544
rect 38068 16532 38074 16584
rect 2225 16507 2283 16513
rect 2225 16473 2237 16507
rect 2271 16504 2283 16507
rect 2590 16504 2596 16516
rect 2271 16476 2596 16504
rect 2271 16473 2283 16476
rect 2225 16467 2283 16473
rect 2590 16464 2596 16476
rect 2648 16464 2654 16516
rect 4614 16464 4620 16516
rect 4672 16504 4678 16516
rect 6270 16504 6276 16516
rect 4672 16476 6276 16504
rect 4672 16464 4678 16476
rect 6270 16464 6276 16476
rect 6328 16464 6334 16516
rect 6638 16464 6644 16516
rect 6696 16504 6702 16516
rect 6825 16507 6883 16513
rect 6825 16504 6837 16507
rect 6696 16476 6837 16504
rect 6696 16464 6702 16476
rect 6825 16473 6837 16476
rect 6871 16473 6883 16507
rect 6825 16467 6883 16473
rect 8202 16464 8208 16516
rect 8260 16504 8266 16516
rect 9214 16504 9220 16516
rect 8260 16476 8305 16504
rect 9175 16476 9220 16504
rect 8260 16464 8266 16476
rect 9214 16464 9220 16476
rect 9272 16464 9278 16516
rect 9318 16507 9376 16513
rect 9318 16473 9330 16507
rect 9364 16504 9376 16507
rect 9582 16504 9588 16516
rect 9364 16476 9588 16504
rect 9364 16473 9376 16476
rect 9318 16467 9376 16473
rect 9582 16464 9588 16476
rect 9640 16464 9646 16516
rect 11609 16507 11667 16513
rect 11609 16473 11621 16507
rect 11655 16504 11667 16507
rect 14642 16504 14648 16516
rect 11655 16476 14648 16504
rect 11655 16473 11667 16476
rect 11609 16467 11667 16473
rect 14642 16464 14648 16476
rect 14700 16464 14706 16516
rect 17034 16464 17040 16516
rect 17092 16504 17098 16516
rect 20165 16507 20223 16513
rect 20165 16504 20177 16507
rect 17092 16476 20177 16504
rect 17092 16464 17098 16476
rect 20165 16473 20177 16476
rect 20211 16473 20223 16507
rect 21818 16504 21824 16516
rect 20165 16467 20223 16473
rect 20732 16476 21824 16504
rect 2958 16436 2964 16448
rect 2919 16408 2964 16436
rect 2958 16396 2964 16408
rect 3016 16396 3022 16448
rect 3970 16436 3976 16448
rect 3931 16408 3976 16436
rect 3970 16396 3976 16408
rect 4028 16396 4034 16448
rect 5534 16396 5540 16448
rect 5592 16436 5598 16448
rect 5629 16439 5687 16445
rect 5629 16436 5641 16439
rect 5592 16408 5641 16436
rect 5592 16396 5598 16408
rect 5629 16405 5641 16408
rect 5675 16405 5687 16439
rect 5629 16399 5687 16405
rect 5902 16396 5908 16448
rect 5960 16436 5966 16448
rect 10594 16436 10600 16448
rect 5960 16408 10600 16436
rect 5960 16396 5966 16408
rect 10594 16396 10600 16408
rect 10652 16396 10658 16448
rect 10962 16436 10968 16448
rect 10923 16408 10968 16436
rect 10962 16396 10968 16408
rect 11020 16396 11026 16448
rect 13630 16436 13636 16448
rect 13591 16408 13636 16436
rect 13630 16396 13636 16408
rect 13688 16396 13694 16448
rect 16666 16396 16672 16448
rect 16724 16436 16730 16448
rect 20732 16436 20760 16476
rect 21818 16464 21824 16476
rect 21876 16464 21882 16516
rect 22002 16464 22008 16516
rect 22060 16504 22066 16516
rect 22922 16504 22928 16516
rect 22060 16476 22928 16504
rect 22060 16464 22066 16476
rect 22922 16464 22928 16476
rect 22980 16464 22986 16516
rect 23017 16507 23075 16513
rect 23017 16473 23029 16507
rect 23063 16504 23075 16507
rect 26326 16504 26332 16516
rect 23063 16476 26332 16504
rect 23063 16473 23075 16476
rect 23017 16467 23075 16473
rect 26326 16464 26332 16476
rect 26384 16464 26390 16516
rect 16724 16408 20760 16436
rect 16724 16396 16730 16408
rect 20806 16396 20812 16448
rect 20864 16436 20870 16448
rect 21266 16436 21272 16448
rect 20864 16408 21272 16436
rect 20864 16396 20870 16408
rect 21266 16396 21272 16408
rect 21324 16396 21330 16448
rect 23566 16436 23572 16448
rect 23527 16408 23572 16436
rect 23566 16396 23572 16408
rect 23624 16396 23630 16448
rect 24670 16436 24676 16448
rect 24631 16408 24676 16436
rect 24670 16396 24676 16408
rect 24728 16396 24734 16448
rect 25225 16439 25283 16445
rect 25225 16405 25237 16439
rect 25271 16436 25283 16439
rect 25774 16436 25780 16448
rect 25271 16408 25780 16436
rect 25271 16405 25283 16408
rect 25225 16399 25283 16405
rect 25774 16396 25780 16408
rect 25832 16396 25838 16448
rect 26053 16439 26111 16445
rect 26053 16405 26065 16439
rect 26099 16436 26111 16439
rect 27338 16436 27344 16448
rect 26099 16408 27344 16436
rect 26099 16405 26111 16408
rect 26053 16399 26111 16405
rect 27338 16396 27344 16408
rect 27396 16396 27402 16448
rect 27430 16396 27436 16448
rect 27488 16436 27494 16448
rect 27893 16439 27951 16445
rect 27893 16436 27905 16439
rect 27488 16408 27905 16436
rect 27488 16396 27494 16408
rect 27893 16405 27905 16408
rect 27939 16405 27951 16439
rect 38194 16436 38200 16448
rect 38155 16408 38200 16436
rect 27893 16399 27951 16405
rect 38194 16396 38200 16408
rect 38252 16396 38258 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 3970 16232 3976 16244
rect 1596 16204 3976 16232
rect 1596 16105 1624 16204
rect 3970 16192 3976 16204
rect 4028 16192 4034 16244
rect 5258 16232 5264 16244
rect 5219 16204 5264 16232
rect 5258 16192 5264 16204
rect 5316 16192 5322 16244
rect 5905 16235 5963 16241
rect 5905 16201 5917 16235
rect 5951 16232 5963 16235
rect 7374 16232 7380 16244
rect 5951 16204 7380 16232
rect 5951 16201 5963 16204
rect 5905 16195 5963 16201
rect 7374 16192 7380 16204
rect 7432 16192 7438 16244
rect 7742 16232 7748 16244
rect 7703 16204 7748 16232
rect 7742 16192 7748 16204
rect 7800 16192 7806 16244
rect 7926 16192 7932 16244
rect 7984 16232 7990 16244
rect 9490 16232 9496 16244
rect 7984 16204 9496 16232
rect 7984 16192 7990 16204
rect 9490 16192 9496 16204
rect 9548 16192 9554 16244
rect 10413 16235 10471 16241
rect 10413 16201 10425 16235
rect 10459 16232 10471 16235
rect 10502 16232 10508 16244
rect 10459 16204 10508 16232
rect 10459 16201 10471 16204
rect 10413 16195 10471 16201
rect 10502 16192 10508 16204
rect 10560 16192 10566 16244
rect 10962 16192 10968 16244
rect 11020 16232 11026 16244
rect 12618 16232 12624 16244
rect 11020 16204 12624 16232
rect 11020 16192 11026 16204
rect 12618 16192 12624 16204
rect 12676 16192 12682 16244
rect 16390 16192 16396 16244
rect 16448 16232 16454 16244
rect 16945 16235 17003 16241
rect 16945 16232 16957 16235
rect 16448 16204 16957 16232
rect 16448 16192 16454 16204
rect 16945 16201 16957 16204
rect 16991 16201 17003 16235
rect 20162 16232 20168 16244
rect 16945 16195 17003 16201
rect 17052 16204 20168 16232
rect 3053 16167 3111 16173
rect 3053 16133 3065 16167
rect 3099 16164 3111 16167
rect 4525 16167 4583 16173
rect 3099 16136 4292 16164
rect 3099 16133 3111 16136
rect 3053 16127 3111 16133
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16065 1639 16099
rect 1581 16059 1639 16065
rect 2958 16028 2964 16040
rect 2871 16000 2964 16028
rect 2958 15988 2964 16000
rect 3016 15988 3022 16040
rect 3602 16028 3608 16040
rect 3563 16000 3608 16028
rect 3602 15988 3608 16000
rect 3660 15988 3666 16040
rect 4264 16028 4292 16136
rect 4525 16133 4537 16167
rect 4571 16164 4583 16167
rect 5442 16164 5448 16176
rect 4571 16136 5448 16164
rect 4571 16133 4583 16136
rect 4525 16127 4583 16133
rect 5442 16124 5448 16136
rect 5500 16124 5506 16176
rect 6270 16124 6276 16176
rect 6328 16164 6334 16176
rect 7285 16167 7343 16173
rect 6328 16136 7236 16164
rect 6328 16124 6334 16136
rect 4433 16099 4491 16105
rect 4433 16065 4445 16099
rect 4479 16096 4491 16099
rect 5169 16099 5227 16105
rect 5169 16096 5181 16099
rect 4479 16068 5181 16096
rect 4479 16065 4491 16068
rect 4433 16059 4491 16065
rect 5169 16065 5181 16068
rect 5215 16096 5227 16099
rect 5258 16096 5264 16108
rect 5215 16068 5264 16096
rect 5215 16065 5227 16068
rect 5169 16059 5227 16065
rect 5258 16056 5264 16068
rect 5316 16056 5322 16108
rect 5626 16056 5632 16108
rect 5684 16096 5690 16108
rect 5813 16099 5871 16105
rect 5813 16096 5825 16099
rect 5684 16068 5825 16096
rect 5684 16056 5690 16068
rect 5813 16065 5825 16068
rect 5859 16096 5871 16099
rect 6178 16096 6184 16108
rect 5859 16068 6184 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 6178 16056 6184 16068
rect 6236 16056 6242 16108
rect 7208 16105 7236 16136
rect 7285 16133 7297 16167
rect 7331 16164 7343 16167
rect 9033 16167 9091 16173
rect 9033 16164 9045 16167
rect 7331 16136 9045 16164
rect 7331 16133 7343 16136
rect 7285 16127 7343 16133
rect 9033 16133 9045 16136
rect 9079 16133 9091 16167
rect 9033 16127 9091 16133
rect 9398 16124 9404 16176
rect 9456 16164 9462 16176
rect 11054 16164 11060 16176
rect 9456 16136 9628 16164
rect 9456 16124 9462 16136
rect 6549 16099 6607 16105
rect 6549 16065 6561 16099
rect 6595 16065 6607 16099
rect 6549 16059 6607 16065
rect 7193 16099 7251 16105
rect 7193 16065 7205 16099
rect 7239 16065 7251 16099
rect 7650 16096 7656 16108
rect 7611 16068 7656 16096
rect 7193 16059 7251 16065
rect 4706 16028 4712 16040
rect 4264 16000 4712 16028
rect 4706 15988 4712 16000
rect 4764 15988 4770 16040
rect 5074 15988 5080 16040
rect 5132 16028 5138 16040
rect 6564 16028 6592 16059
rect 7650 16056 7656 16068
rect 7708 16056 7714 16108
rect 8478 16096 8484 16108
rect 8439 16068 8484 16096
rect 8478 16056 8484 16068
rect 8536 16056 8542 16108
rect 9333 16086 9444 16096
rect 9490 16086 9496 16108
rect 9333 16068 9496 16086
rect 7926 16028 7932 16040
rect 5132 16000 6500 16028
rect 6564 16000 7932 16028
rect 5132 15988 5138 16000
rect 2976 15960 3004 15988
rect 6270 15960 6276 15972
rect 2976 15932 6276 15960
rect 6270 15920 6276 15932
rect 6328 15920 6334 15972
rect 6472 15960 6500 16000
rect 7926 15988 7932 16000
rect 7984 15988 7990 16040
rect 8205 16031 8263 16037
rect 8205 15997 8217 16031
rect 8251 16028 8263 16031
rect 9125 16031 9183 16037
rect 9125 16028 9137 16031
rect 8251 16000 9137 16028
rect 8251 15997 8263 16000
rect 8205 15991 8263 15997
rect 9125 15997 9137 16000
rect 9171 16028 9183 16031
rect 9333 16028 9361 16068
rect 9416 16058 9496 16068
rect 9490 16056 9496 16058
rect 9548 16056 9554 16108
rect 9600 16086 9628 16136
rect 9784 16136 11060 16164
rect 9677 16099 9735 16105
rect 9677 16086 9689 16099
rect 9600 16065 9689 16086
rect 9723 16086 9735 16099
rect 9784 16086 9812 16136
rect 11054 16124 11060 16136
rect 11112 16124 11118 16176
rect 11146 16124 11152 16176
rect 11204 16164 11210 16176
rect 16666 16164 16672 16176
rect 11204 16136 16672 16164
rect 11204 16124 11210 16136
rect 16666 16124 16672 16136
rect 16724 16124 16730 16176
rect 10318 16096 10324 16108
rect 9723 16065 9815 16086
rect 10279 16068 10324 16096
rect 9600 16058 9815 16065
rect 10318 16056 10324 16068
rect 10376 16056 10382 16108
rect 10410 16056 10416 16108
rect 10468 16096 10474 16108
rect 16853 16099 16911 16105
rect 16853 16096 16865 16099
rect 10468 16068 16865 16096
rect 10468 16056 10474 16068
rect 16853 16065 16865 16068
rect 16899 16065 16911 16099
rect 16853 16059 16911 16065
rect 9171 16000 9361 16028
rect 9171 15997 9183 16000
rect 9125 15991 9183 15997
rect 10594 15988 10600 16040
rect 10652 16028 10658 16040
rect 17052 16028 17080 16204
rect 20162 16192 20168 16204
rect 20220 16192 20226 16244
rect 22554 16192 22560 16244
rect 22612 16232 22618 16244
rect 23109 16235 23167 16241
rect 23109 16232 23121 16235
rect 22612 16204 23121 16232
rect 22612 16192 22618 16204
rect 23109 16201 23121 16204
rect 23155 16201 23167 16235
rect 23109 16195 23167 16201
rect 25593 16235 25651 16241
rect 25593 16201 25605 16235
rect 25639 16232 25651 16235
rect 26142 16232 26148 16244
rect 25639 16204 26148 16232
rect 25639 16201 25651 16204
rect 25593 16195 25651 16201
rect 26142 16192 26148 16204
rect 26200 16192 26206 16244
rect 27614 16232 27620 16244
rect 26252 16204 27620 16232
rect 17954 16124 17960 16176
rect 18012 16164 18018 16176
rect 18233 16167 18291 16173
rect 18233 16164 18245 16167
rect 18012 16136 18245 16164
rect 18012 16124 18018 16136
rect 18233 16133 18245 16136
rect 18279 16133 18291 16167
rect 18233 16127 18291 16133
rect 19153 16167 19211 16173
rect 19153 16133 19165 16167
rect 19199 16164 19211 16167
rect 20714 16164 20720 16176
rect 19199 16136 20720 16164
rect 19199 16133 19211 16136
rect 19153 16127 19211 16133
rect 20714 16124 20720 16136
rect 20772 16124 20778 16176
rect 23566 16124 23572 16176
rect 23624 16164 23630 16176
rect 26252 16164 26280 16204
rect 27614 16192 27620 16204
rect 27672 16192 27678 16244
rect 29730 16192 29736 16244
rect 29788 16232 29794 16244
rect 30101 16235 30159 16241
rect 30101 16232 30113 16235
rect 29788 16204 30113 16232
rect 29788 16192 29794 16204
rect 30101 16201 30113 16204
rect 30147 16201 30159 16235
rect 30101 16195 30159 16201
rect 23624 16136 26280 16164
rect 23624 16124 23630 16136
rect 27246 16124 27252 16176
rect 27304 16164 27310 16176
rect 27341 16167 27399 16173
rect 27341 16164 27353 16167
rect 27304 16136 27353 16164
rect 27304 16124 27310 16136
rect 27341 16133 27353 16136
rect 27387 16133 27399 16167
rect 27341 16127 27399 16133
rect 19978 16056 19984 16108
rect 20036 16096 20042 16108
rect 20073 16099 20131 16105
rect 20073 16096 20085 16099
rect 20036 16068 20085 16096
rect 20036 16056 20042 16068
rect 20073 16065 20085 16068
rect 20119 16065 20131 16099
rect 20073 16059 20131 16065
rect 21542 16056 21548 16108
rect 21600 16096 21606 16108
rect 23017 16099 23075 16105
rect 23017 16096 23029 16099
rect 21600 16068 23029 16096
rect 21600 16056 21606 16068
rect 23017 16065 23029 16068
rect 23063 16096 23075 16099
rect 25406 16096 25412 16108
rect 23063 16068 25412 16096
rect 23063 16065 23075 16068
rect 23017 16059 23075 16065
rect 25406 16056 25412 16068
rect 25464 16056 25470 16108
rect 25774 16096 25780 16108
rect 25735 16068 25780 16096
rect 25774 16056 25780 16068
rect 25832 16056 25838 16108
rect 28994 16096 29000 16108
rect 28955 16068 29000 16096
rect 28994 16056 29000 16068
rect 29052 16056 29058 16108
rect 30009 16099 30067 16105
rect 30009 16065 30021 16099
rect 30055 16096 30067 16099
rect 30055 16068 35894 16096
rect 30055 16065 30067 16068
rect 30009 16059 30067 16065
rect 10652 16000 17080 16028
rect 18141 16031 18199 16037
rect 10652 15988 10658 16000
rect 18141 15997 18153 16031
rect 18187 16028 18199 16031
rect 18414 16028 18420 16040
rect 18187 16000 18420 16028
rect 18187 15997 18199 16000
rect 18141 15991 18199 15997
rect 18414 15988 18420 16000
rect 18472 15988 18478 16040
rect 20257 16031 20315 16037
rect 20257 15997 20269 16031
rect 20303 16028 20315 16031
rect 20990 16028 20996 16040
rect 20303 16000 20996 16028
rect 20303 15997 20315 16000
rect 20257 15991 20315 15997
rect 20990 15988 20996 16000
rect 21048 15988 21054 16040
rect 26326 15988 26332 16040
rect 26384 16028 26390 16040
rect 27249 16031 27307 16037
rect 27249 16028 27261 16031
rect 26384 16000 27261 16028
rect 26384 15988 26390 16000
rect 27249 15997 27261 16000
rect 27295 15997 27307 16031
rect 27890 16028 27896 16040
rect 27851 16000 27896 16028
rect 27249 15991 27307 15997
rect 27890 15988 27896 16000
rect 27948 15988 27954 16040
rect 35866 16028 35894 16068
rect 36906 16056 36912 16108
rect 36964 16096 36970 16108
rect 38013 16099 38071 16105
rect 38013 16096 38025 16099
rect 36964 16068 38025 16096
rect 36964 16056 36970 16068
rect 38013 16065 38025 16068
rect 38059 16065 38071 16099
rect 38013 16059 38071 16065
rect 37734 16028 37740 16040
rect 35866 16000 37740 16028
rect 37734 15988 37740 16000
rect 37792 15988 37798 16040
rect 6472 15932 7880 15960
rect 1762 15892 1768 15904
rect 1723 15864 1768 15892
rect 1762 15852 1768 15864
rect 1820 15852 1826 15904
rect 6638 15892 6644 15904
rect 6599 15864 6644 15892
rect 6638 15852 6644 15864
rect 6696 15852 6702 15904
rect 7852 15892 7880 15932
rect 9490 15920 9496 15972
rect 9548 15960 9554 15972
rect 22830 15960 22836 15972
rect 9548 15932 22836 15960
rect 9548 15920 9554 15932
rect 22830 15920 22836 15932
rect 22888 15920 22894 15972
rect 24670 15920 24676 15972
rect 24728 15960 24734 15972
rect 28166 15960 28172 15972
rect 24728 15932 28172 15960
rect 24728 15920 24734 15932
rect 28166 15920 28172 15932
rect 28224 15920 28230 15972
rect 28813 15963 28871 15969
rect 28813 15929 28825 15963
rect 28859 15960 28871 15963
rect 28859 15932 35894 15960
rect 28859 15929 28871 15932
rect 28813 15923 28871 15929
rect 9769 15895 9827 15901
rect 9769 15892 9781 15895
rect 7852 15864 9781 15892
rect 9769 15861 9781 15864
rect 9815 15861 9827 15895
rect 9769 15855 9827 15861
rect 10226 15852 10232 15904
rect 10284 15892 10290 15904
rect 20346 15892 20352 15904
rect 10284 15864 20352 15892
rect 10284 15852 10290 15864
rect 20346 15852 20352 15864
rect 20404 15852 20410 15904
rect 20714 15892 20720 15904
rect 20675 15864 20720 15892
rect 20714 15852 20720 15864
rect 20772 15852 20778 15904
rect 35866 15892 35894 15932
rect 38010 15892 38016 15904
rect 35866 15864 38016 15892
rect 38010 15852 38016 15864
rect 38068 15852 38074 15904
rect 38194 15892 38200 15904
rect 38155 15864 38200 15892
rect 38194 15852 38200 15864
rect 38252 15852 38258 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 1854 15648 1860 15700
rect 1912 15688 1918 15700
rect 3326 15688 3332 15700
rect 1912 15660 3188 15688
rect 3287 15660 3332 15688
rect 1912 15648 1918 15660
rect 2774 15620 2780 15632
rect 2148 15592 2780 15620
rect 2148 15561 2176 15592
rect 2774 15580 2780 15592
rect 2832 15580 2838 15632
rect 3160 15620 3188 15660
rect 3326 15648 3332 15660
rect 3384 15648 3390 15700
rect 4062 15688 4068 15700
rect 4023 15660 4068 15688
rect 4062 15648 4068 15660
rect 4120 15648 4126 15700
rect 4801 15691 4859 15697
rect 4801 15657 4813 15691
rect 4847 15688 4859 15691
rect 5810 15688 5816 15700
rect 4847 15660 5816 15688
rect 4847 15657 4859 15660
rect 4801 15651 4859 15657
rect 5810 15648 5816 15660
rect 5868 15648 5874 15700
rect 6730 15688 6736 15700
rect 6691 15660 6736 15688
rect 6730 15648 6736 15660
rect 6788 15648 6794 15700
rect 7837 15691 7895 15697
rect 7837 15657 7849 15691
rect 7883 15688 7895 15691
rect 8662 15688 8668 15700
rect 7883 15660 8668 15688
rect 7883 15657 7895 15660
rect 7837 15651 7895 15657
rect 8662 15648 8668 15660
rect 8720 15648 8726 15700
rect 9030 15648 9036 15700
rect 9088 15688 9094 15700
rect 9217 15691 9275 15697
rect 9217 15688 9229 15691
rect 9088 15660 9229 15688
rect 9088 15648 9094 15660
rect 9217 15657 9229 15660
rect 9263 15657 9275 15691
rect 10594 15688 10600 15700
rect 10555 15660 10600 15688
rect 9217 15651 9275 15657
rect 10594 15648 10600 15660
rect 10652 15648 10658 15700
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 14550 15688 14556 15700
rect 12492 15660 12572 15688
rect 14511 15660 14556 15688
rect 12492 15648 12498 15660
rect 5258 15620 5264 15632
rect 3160 15592 5264 15620
rect 5258 15580 5264 15592
rect 5316 15580 5322 15632
rect 5445 15623 5503 15629
rect 5445 15589 5457 15623
rect 5491 15620 5503 15623
rect 6914 15620 6920 15632
rect 5491 15592 6920 15620
rect 5491 15589 5503 15592
rect 5445 15583 5503 15589
rect 6914 15580 6920 15592
rect 6972 15580 6978 15632
rect 8294 15580 8300 15632
rect 8352 15620 8358 15632
rect 8754 15620 8760 15632
rect 8352 15592 8760 15620
rect 8352 15580 8358 15592
rect 8754 15580 8760 15592
rect 8812 15580 8818 15632
rect 9306 15580 9312 15632
rect 9364 15620 9370 15632
rect 10226 15620 10232 15632
rect 9364 15592 10232 15620
rect 9364 15580 9370 15592
rect 10226 15580 10232 15592
rect 10284 15580 10290 15632
rect 12544 15620 12572 15660
rect 14550 15648 14556 15660
rect 14608 15648 14614 15700
rect 15470 15688 15476 15700
rect 15431 15660 15476 15688
rect 15470 15648 15476 15660
rect 15528 15648 15534 15700
rect 15838 15648 15844 15700
rect 15896 15688 15902 15700
rect 16298 15688 16304 15700
rect 15896 15660 16304 15688
rect 15896 15648 15902 15660
rect 16298 15648 16304 15660
rect 16356 15648 16362 15700
rect 16758 15688 16764 15700
rect 16719 15660 16764 15688
rect 16758 15648 16764 15660
rect 16816 15648 16822 15700
rect 17954 15648 17960 15700
rect 18012 15688 18018 15700
rect 18049 15691 18107 15697
rect 18049 15688 18061 15691
rect 18012 15660 18061 15688
rect 18012 15648 18018 15660
rect 18049 15657 18061 15660
rect 18095 15657 18107 15691
rect 18049 15651 18107 15657
rect 18138 15648 18144 15700
rect 18196 15688 18202 15700
rect 22002 15688 22008 15700
rect 18196 15660 22008 15688
rect 18196 15648 18202 15660
rect 22002 15648 22008 15660
rect 22060 15648 22066 15700
rect 23569 15691 23627 15697
rect 23569 15657 23581 15691
rect 23615 15688 23627 15691
rect 23842 15688 23848 15700
rect 23615 15660 23848 15688
rect 23615 15657 23627 15660
rect 23569 15651 23627 15657
rect 23842 15648 23848 15660
rect 23900 15648 23906 15700
rect 18782 15620 18788 15632
rect 12544 15592 18788 15620
rect 18782 15580 18788 15592
rect 18840 15580 18846 15632
rect 2133 15555 2191 15561
rect 2133 15521 2145 15555
rect 2179 15521 2191 15555
rect 2133 15515 2191 15521
rect 2314 15512 2320 15564
rect 2372 15552 2378 15564
rect 2409 15555 2467 15561
rect 2409 15552 2421 15555
rect 2372 15524 2421 15552
rect 2372 15512 2378 15524
rect 2409 15521 2421 15524
rect 2455 15521 2467 15555
rect 2409 15515 2467 15521
rect 6089 15555 6147 15561
rect 6089 15521 6101 15555
rect 6135 15552 6147 15555
rect 8846 15552 8852 15564
rect 6135 15524 8852 15552
rect 6135 15521 6147 15524
rect 6089 15515 6147 15521
rect 8846 15512 8852 15524
rect 8904 15512 8910 15564
rect 9398 15552 9404 15564
rect 8956 15524 9404 15552
rect 3237 15487 3295 15493
rect 3237 15453 3249 15487
rect 3283 15453 3295 15487
rect 3970 15484 3976 15496
rect 3931 15456 3976 15484
rect 3237 15447 3295 15453
rect 2225 15419 2283 15425
rect 2225 15385 2237 15419
rect 2271 15385 2283 15419
rect 3252 15416 3280 15447
rect 3970 15444 3976 15456
rect 4028 15444 4034 15496
rect 4709 15487 4767 15493
rect 4709 15453 4721 15487
rect 4755 15453 4767 15487
rect 4709 15447 4767 15453
rect 5353 15487 5411 15493
rect 5353 15453 5365 15487
rect 5399 15484 5411 15487
rect 5626 15484 5632 15496
rect 5399 15456 5632 15484
rect 5399 15453 5411 15456
rect 5353 15447 5411 15453
rect 4724 15416 4752 15447
rect 5626 15444 5632 15456
rect 5684 15444 5690 15496
rect 5902 15444 5908 15496
rect 5960 15484 5966 15496
rect 5997 15487 6055 15493
rect 5997 15484 6009 15487
rect 5960 15456 6009 15484
rect 5960 15444 5966 15456
rect 5997 15453 6009 15456
rect 6043 15453 6055 15487
rect 5997 15447 6055 15453
rect 6178 15444 6184 15496
rect 6236 15484 6242 15496
rect 6641 15487 6699 15493
rect 6641 15484 6653 15487
rect 6236 15456 6653 15484
rect 6236 15444 6242 15456
rect 6641 15453 6653 15456
rect 6687 15484 6699 15487
rect 6822 15484 6828 15496
rect 6687 15456 6828 15484
rect 6687 15453 6699 15456
rect 6641 15447 6699 15453
rect 6822 15444 6828 15456
rect 6880 15444 6886 15496
rect 6914 15444 6920 15496
rect 6972 15484 6978 15496
rect 7745 15487 7803 15493
rect 7745 15484 7757 15487
rect 6972 15456 7757 15484
rect 6972 15444 6978 15456
rect 7745 15453 7757 15456
rect 7791 15484 7803 15487
rect 8294 15484 8300 15496
rect 7791 15456 8300 15484
rect 7791 15453 7803 15456
rect 7745 15447 7803 15453
rect 8294 15444 8300 15456
rect 8352 15444 8358 15496
rect 8389 15487 8447 15493
rect 8389 15453 8401 15487
rect 8435 15484 8447 15487
rect 8956 15484 8984 15524
rect 9398 15512 9404 15524
rect 9456 15512 9462 15564
rect 9582 15512 9588 15564
rect 9640 15552 9646 15564
rect 12713 15555 12771 15561
rect 12713 15552 12725 15555
rect 9640 15524 12725 15552
rect 9640 15512 9646 15524
rect 12713 15521 12725 15524
rect 12759 15521 12771 15555
rect 12713 15515 12771 15521
rect 12802 15512 12808 15564
rect 12860 15552 12866 15564
rect 16132 15561 16252 15564
rect 16117 15555 16252 15561
rect 12860 15524 15608 15552
rect 12860 15512 12866 15524
rect 9122 15484 9128 15496
rect 8435 15456 8984 15484
rect 9083 15456 9128 15484
rect 8435 15453 8447 15456
rect 8389 15447 8447 15453
rect 3252 15388 4752 15416
rect 2225 15379 2283 15385
rect 1854 15308 1860 15360
rect 1912 15348 1918 15360
rect 2240 15348 2268 15379
rect 1912 15320 2268 15348
rect 4724 15348 4752 15388
rect 7650 15376 7656 15428
rect 7708 15416 7714 15428
rect 8404 15416 8432 15447
rect 9122 15444 9128 15456
rect 9180 15444 9186 15496
rect 10410 15444 10416 15496
rect 10468 15484 10474 15496
rect 10505 15487 10563 15493
rect 10505 15484 10517 15487
rect 10468 15456 10517 15484
rect 10468 15444 10474 15456
rect 10505 15453 10517 15456
rect 10551 15453 10563 15487
rect 10505 15447 10563 15453
rect 7708 15388 8432 15416
rect 10520 15416 10548 15447
rect 11606 15444 11612 15496
rect 11664 15484 11670 15496
rect 11977 15487 12035 15493
rect 11977 15484 11989 15487
rect 11664 15456 11989 15484
rect 11664 15444 11670 15456
rect 11977 15453 11989 15456
rect 12023 15453 12035 15487
rect 11977 15447 12035 15453
rect 14461 15487 14519 15493
rect 14461 15453 14473 15487
rect 14507 15484 14519 15487
rect 15381 15487 15439 15493
rect 15381 15484 15393 15487
rect 14507 15456 15393 15484
rect 14507 15453 14519 15456
rect 14461 15447 14519 15453
rect 15381 15453 15393 15456
rect 15427 15484 15439 15487
rect 15470 15484 15476 15496
rect 15427 15456 15476 15484
rect 15427 15453 15439 15456
rect 15381 15447 15439 15453
rect 15470 15444 15476 15456
rect 15528 15444 15534 15496
rect 15580 15484 15608 15524
rect 16117 15521 16129 15555
rect 16163 15552 16252 15555
rect 20533 15555 20591 15561
rect 16163 15536 20116 15552
rect 16163 15521 16175 15536
rect 16224 15524 20116 15536
rect 16117 15515 16175 15521
rect 16669 15487 16727 15493
rect 15580 15478 15976 15484
rect 16017 15481 16075 15487
rect 16017 15478 16029 15481
rect 15580 15456 16029 15478
rect 15948 15450 16029 15456
rect 16017 15447 16029 15450
rect 16063 15447 16075 15481
rect 16669 15453 16681 15487
rect 16715 15484 16727 15487
rect 17034 15484 17040 15496
rect 16715 15456 17040 15484
rect 16715 15453 16727 15456
rect 16669 15447 16727 15453
rect 16017 15441 16075 15447
rect 17034 15444 17040 15456
rect 17092 15484 17098 15496
rect 17862 15484 17868 15496
rect 17092 15456 17868 15484
rect 17092 15444 17098 15456
rect 17862 15444 17868 15456
rect 17920 15444 17926 15496
rect 17957 15487 18015 15493
rect 17957 15453 17969 15487
rect 18003 15484 18015 15487
rect 18046 15484 18052 15496
rect 18003 15456 18052 15484
rect 18003 15453 18015 15456
rect 17957 15447 18015 15453
rect 18046 15444 18052 15456
rect 18104 15444 18110 15496
rect 19886 15484 19892 15496
rect 19720 15456 19892 15484
rect 12805 15419 12863 15425
rect 10520 15388 12434 15416
rect 7708 15376 7714 15388
rect 5442 15348 5448 15360
rect 4724 15320 5448 15348
rect 1912 15308 1918 15320
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 5994 15308 6000 15360
rect 6052 15348 6058 15360
rect 8481 15351 8539 15357
rect 8481 15348 8493 15351
rect 6052 15320 8493 15348
rect 6052 15308 6058 15320
rect 8481 15317 8493 15320
rect 8527 15317 8539 15351
rect 8481 15311 8539 15317
rect 11974 15308 11980 15360
rect 12032 15348 12038 15360
rect 12069 15351 12127 15357
rect 12069 15348 12081 15351
rect 12032 15320 12081 15348
rect 12032 15308 12038 15320
rect 12069 15317 12081 15320
rect 12115 15317 12127 15351
rect 12406 15348 12434 15388
rect 12805 15385 12817 15419
rect 12851 15416 12863 15419
rect 13630 15416 13636 15428
rect 12851 15388 13636 15416
rect 12851 15385 12863 15388
rect 12805 15379 12863 15385
rect 13630 15376 13636 15388
rect 13688 15376 13694 15428
rect 13725 15419 13783 15425
rect 13725 15385 13737 15419
rect 13771 15416 13783 15419
rect 15838 15416 15844 15428
rect 13771 15388 15844 15416
rect 13771 15385 13783 15388
rect 13725 15379 13783 15385
rect 15838 15376 15844 15388
rect 15896 15376 15902 15428
rect 16298 15376 16304 15428
rect 16356 15416 16362 15428
rect 19720 15416 19748 15456
rect 19886 15444 19892 15456
rect 19944 15444 19950 15496
rect 16356 15388 19748 15416
rect 19797 15419 19855 15425
rect 16356 15376 16362 15388
rect 19797 15385 19809 15419
rect 19843 15416 19855 15419
rect 19978 15416 19984 15428
rect 19843 15388 19984 15416
rect 19843 15385 19855 15388
rect 19797 15379 19855 15385
rect 19978 15376 19984 15388
rect 20036 15376 20042 15428
rect 20088 15416 20116 15524
rect 20533 15521 20545 15555
rect 20579 15552 20591 15555
rect 24670 15552 24676 15564
rect 20579 15524 24676 15552
rect 20579 15521 20591 15524
rect 20533 15515 20591 15521
rect 24670 15512 24676 15524
rect 24728 15512 24734 15564
rect 26878 15512 26884 15564
rect 26936 15552 26942 15564
rect 27617 15555 27675 15561
rect 27617 15552 27629 15555
rect 26936 15524 27629 15552
rect 26936 15512 26942 15524
rect 27617 15521 27629 15524
rect 27663 15521 27675 15555
rect 27617 15515 27675 15521
rect 22922 15444 22928 15496
rect 22980 15484 22986 15496
rect 23382 15484 23388 15496
rect 22980 15456 23388 15484
rect 22980 15444 22986 15456
rect 23382 15444 23388 15456
rect 23440 15484 23446 15496
rect 23477 15487 23535 15493
rect 23477 15484 23489 15487
rect 23440 15456 23489 15484
rect 23440 15444 23446 15456
rect 23477 15453 23489 15456
rect 23523 15453 23535 15487
rect 23477 15447 23535 15453
rect 20625 15419 20683 15425
rect 20625 15416 20637 15419
rect 20088 15388 20637 15416
rect 20625 15385 20637 15388
rect 20671 15385 20683 15419
rect 21174 15416 21180 15428
rect 21135 15388 21180 15416
rect 20625 15379 20683 15385
rect 21174 15376 21180 15388
rect 21232 15376 21238 15428
rect 22066 15388 23704 15416
rect 13078 15348 13084 15360
rect 12406 15320 13084 15348
rect 12069 15311 12127 15317
rect 13078 15308 13084 15320
rect 13136 15308 13142 15360
rect 15930 15308 15936 15360
rect 15988 15348 15994 15360
rect 18138 15348 18144 15360
rect 15988 15320 18144 15348
rect 15988 15308 15994 15320
rect 18138 15308 18144 15320
rect 18196 15308 18202 15360
rect 19889 15351 19947 15357
rect 19889 15317 19901 15351
rect 19935 15348 19947 15351
rect 22066 15348 22094 15388
rect 19935 15320 22094 15348
rect 23676 15348 23704 15388
rect 26510 15376 26516 15428
rect 26568 15416 26574 15428
rect 27341 15419 27399 15425
rect 27341 15416 27353 15419
rect 26568 15388 27353 15416
rect 26568 15376 26574 15388
rect 27341 15385 27353 15388
rect 27387 15385 27399 15419
rect 27341 15379 27399 15385
rect 27430 15376 27436 15428
rect 27488 15416 27494 15428
rect 27488 15388 27533 15416
rect 27488 15376 27494 15388
rect 37274 15348 37280 15360
rect 23676 15320 37280 15348
rect 19935 15317 19947 15320
rect 19889 15311 19947 15317
rect 37274 15308 37280 15320
rect 37332 15308 37338 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 4614 15144 4620 15156
rect 1964 15116 4620 15144
rect 1964 15085 1992 15116
rect 4614 15104 4620 15116
rect 4672 15104 4678 15156
rect 4801 15147 4859 15153
rect 4801 15113 4813 15147
rect 4847 15144 4859 15147
rect 4890 15144 4896 15156
rect 4847 15116 4896 15144
rect 4847 15113 4859 15116
rect 4801 15107 4859 15113
rect 4890 15104 4896 15116
rect 4948 15104 4954 15156
rect 7190 15144 7196 15156
rect 6564 15116 7196 15144
rect 1949 15079 2007 15085
rect 1949 15045 1961 15079
rect 1995 15045 2007 15079
rect 1949 15039 2007 15045
rect 4157 15079 4215 15085
rect 4157 15045 4169 15079
rect 4203 15076 4215 15079
rect 6564 15076 6592 15116
rect 7190 15104 7196 15116
rect 7248 15104 7254 15156
rect 14734 15144 14740 15156
rect 7668 15116 14740 15144
rect 4203 15048 6592 15076
rect 4203 15045 4215 15048
rect 4157 15039 4215 15045
rect 6638 15036 6644 15088
rect 6696 15076 6702 15088
rect 6733 15079 6791 15085
rect 6733 15076 6745 15079
rect 6696 15048 6745 15076
rect 6696 15036 6702 15048
rect 6733 15045 6745 15048
rect 6779 15045 6791 15079
rect 6733 15039 6791 15045
rect 6822 15036 6828 15088
rect 6880 15076 6886 15088
rect 7668 15085 7696 15116
rect 14734 15104 14740 15116
rect 14792 15104 14798 15156
rect 15378 15104 15384 15156
rect 15436 15144 15442 15156
rect 16114 15144 16120 15156
rect 15436 15116 16120 15144
rect 15436 15104 15442 15116
rect 16114 15104 16120 15116
rect 16172 15104 16178 15156
rect 16482 15104 16488 15156
rect 16540 15144 16546 15156
rect 17129 15147 17187 15153
rect 17129 15144 17141 15147
rect 16540 15116 17141 15144
rect 16540 15104 16546 15116
rect 17129 15113 17141 15116
rect 17175 15113 17187 15147
rect 17129 15107 17187 15113
rect 18690 15104 18696 15156
rect 18748 15144 18754 15156
rect 19334 15144 19340 15156
rect 18748 15116 19340 15144
rect 18748 15104 18754 15116
rect 19334 15104 19340 15116
rect 19392 15104 19398 15156
rect 20714 15144 20720 15156
rect 20456 15116 20720 15144
rect 7653 15079 7711 15085
rect 6880 15048 7512 15076
rect 6880 15036 6886 15048
rect 4062 15008 4068 15020
rect 3975 14980 4068 15008
rect 4062 14968 4068 14980
rect 4120 15008 4126 15020
rect 4709 15011 4767 15017
rect 4120 14980 4476 15008
rect 4120 14968 4126 14980
rect 1857 14943 1915 14949
rect 1857 14909 1869 14943
rect 1903 14940 1915 14943
rect 2958 14940 2964 14952
rect 1903 14912 2774 14940
rect 2919 14912 2964 14940
rect 1903 14909 1915 14912
rect 1857 14903 1915 14909
rect 2409 14875 2467 14881
rect 2409 14841 2421 14875
rect 2455 14872 2467 14875
rect 2498 14872 2504 14884
rect 2455 14844 2504 14872
rect 2455 14841 2467 14844
rect 2409 14835 2467 14841
rect 2498 14832 2504 14844
rect 2556 14832 2562 14884
rect 2746 14872 2774 14912
rect 2958 14900 2964 14912
rect 3016 14900 3022 14952
rect 3142 14940 3148 14952
rect 3103 14912 3148 14940
rect 3142 14900 3148 14912
rect 3200 14900 3206 14952
rect 4448 14940 4476 14980
rect 4709 14977 4721 15011
rect 4755 15008 4767 15011
rect 5166 15008 5172 15020
rect 4755 14980 5172 15008
rect 4755 14977 4767 14980
rect 4709 14971 4767 14977
rect 5166 14968 5172 14980
rect 5224 14968 5230 15020
rect 5353 15011 5411 15017
rect 5353 14977 5365 15011
rect 5399 15006 5411 15011
rect 5442 15006 5448 15020
rect 5399 14978 5448 15006
rect 5399 14977 5411 14978
rect 5353 14971 5411 14977
rect 5442 14968 5448 14978
rect 5500 14968 5506 15020
rect 7484 15008 7512 15048
rect 7653 15045 7665 15079
rect 7699 15045 7711 15079
rect 7653 15039 7711 15045
rect 8018 15036 8024 15088
rect 8076 15076 8082 15088
rect 8205 15079 8263 15085
rect 8205 15076 8217 15079
rect 8076 15048 8217 15076
rect 8076 15036 8082 15048
rect 8205 15045 8217 15048
rect 8251 15045 8263 15079
rect 8205 15039 8263 15045
rect 8849 15079 8907 15085
rect 8849 15045 8861 15079
rect 8895 15076 8907 15079
rect 9674 15076 9680 15088
rect 8895 15048 9680 15076
rect 8895 15045 8907 15048
rect 8849 15039 8907 15045
rect 9674 15036 9680 15048
rect 9732 15036 9738 15088
rect 11977 15079 12035 15085
rect 11977 15045 11989 15079
rect 12023 15076 12035 15079
rect 13449 15079 13507 15085
rect 13449 15076 13461 15079
rect 12023 15048 13461 15076
rect 12023 15045 12035 15048
rect 11977 15039 12035 15045
rect 13449 15045 13461 15048
rect 13495 15045 13507 15079
rect 13449 15039 13507 15045
rect 15105 15079 15163 15085
rect 15105 15045 15117 15079
rect 15151 15076 15163 15079
rect 20456 15076 20484 15116
rect 20714 15104 20720 15116
rect 20772 15144 20778 15156
rect 24854 15144 24860 15156
rect 20772 15116 21496 15144
rect 24815 15116 24860 15144
rect 20772 15104 20778 15116
rect 20898 15076 20904 15088
rect 15151 15048 20484 15076
rect 20859 15048 20904 15076
rect 15151 15045 15163 15048
rect 15105 15039 15163 15045
rect 20898 15036 20904 15048
rect 20956 15036 20962 15088
rect 8113 15011 8171 15017
rect 8113 15008 8125 15011
rect 7484 14980 8125 15008
rect 8113 14977 8125 14980
rect 8159 15008 8171 15011
rect 8386 15008 8392 15020
rect 8159 14980 8392 15008
rect 8159 14977 8171 14980
rect 8113 14971 8171 14977
rect 8386 14968 8392 14980
rect 8444 14968 8450 15020
rect 8754 15008 8760 15020
rect 8715 14980 8760 15008
rect 8754 14968 8760 14980
rect 8812 14968 8818 15020
rect 9766 15008 9772 15020
rect 9727 14980 9772 15008
rect 9766 14968 9772 14980
rect 9824 14968 9830 15020
rect 13357 15011 13415 15017
rect 13357 15008 13369 15011
rect 12820 14980 13369 15008
rect 5902 14940 5908 14952
rect 4448 14912 5908 14940
rect 5902 14900 5908 14912
rect 5960 14900 5966 14952
rect 6270 14900 6276 14952
rect 6328 14940 6334 14952
rect 6641 14943 6699 14949
rect 6641 14940 6653 14943
rect 6328 14912 6653 14940
rect 6328 14900 6334 14912
rect 6641 14909 6653 14912
rect 6687 14909 6699 14943
rect 6641 14903 6699 14909
rect 6730 14900 6736 14952
rect 6788 14940 6794 14952
rect 11698 14940 11704 14952
rect 6788 14912 11704 14940
rect 6788 14900 6794 14912
rect 11698 14900 11704 14912
rect 11756 14900 11762 14952
rect 11882 14940 11888 14952
rect 11843 14912 11888 14940
rect 11882 14900 11888 14912
rect 11940 14900 11946 14952
rect 12066 14900 12072 14952
rect 12124 14940 12130 14952
rect 12820 14940 12848 14980
rect 13357 14977 13369 14980
rect 13403 14977 13415 15011
rect 16022 15008 16028 15020
rect 13357 14971 13415 14977
rect 13556 14980 16028 15008
rect 12124 14912 12848 14940
rect 12124 14900 12130 14912
rect 12894 14900 12900 14952
rect 12952 14940 12958 14952
rect 13556 14940 13584 14980
rect 16022 14968 16028 14980
rect 16080 14968 16086 15020
rect 17034 15008 17040 15020
rect 16995 14980 17040 15008
rect 17034 14968 17040 14980
rect 17092 14968 17098 15020
rect 18782 15008 18788 15020
rect 18743 14980 18788 15008
rect 18782 14968 18788 14980
rect 18840 14968 18846 15020
rect 18877 15011 18935 15017
rect 18877 14977 18889 15011
rect 18923 15008 18935 15011
rect 21468 15008 21496 15116
rect 24854 15104 24860 15116
rect 24912 15104 24918 15156
rect 24946 15104 24952 15156
rect 25004 15144 25010 15156
rect 26050 15144 26056 15156
rect 25004 15116 26056 15144
rect 25004 15104 25010 15116
rect 26050 15104 26056 15116
rect 26108 15104 26114 15156
rect 26510 15144 26516 15156
rect 26471 15116 26516 15144
rect 26510 15104 26516 15116
rect 26568 15104 26574 15156
rect 27706 15144 27712 15156
rect 27667 15116 27712 15144
rect 27706 15104 27712 15116
rect 27764 15104 27770 15156
rect 35161 15147 35219 15153
rect 35161 15113 35173 15147
rect 35207 15144 35219 15147
rect 36906 15144 36912 15156
rect 35207 15116 36912 15144
rect 35207 15113 35219 15116
rect 35161 15107 35219 15113
rect 36906 15104 36912 15116
rect 36964 15104 36970 15156
rect 23385 15079 23443 15085
rect 23385 15076 23397 15079
rect 22066 15048 23397 15076
rect 22066 15008 22094 15048
rect 23385 15045 23397 15048
rect 23431 15045 23443 15079
rect 23385 15039 23443 15045
rect 23474 15036 23480 15088
rect 23532 15076 23538 15088
rect 24029 15079 24087 15085
rect 23532 15048 23577 15076
rect 23532 15036 23538 15048
rect 24029 15045 24041 15079
rect 24075 15076 24087 15079
rect 27890 15076 27896 15088
rect 24075 15048 27896 15076
rect 24075 15045 24087 15048
rect 24029 15039 24087 15045
rect 27890 15036 27896 15048
rect 27948 15036 27954 15088
rect 18923 14980 19196 15008
rect 21468 14980 22094 15008
rect 24765 15011 24823 15017
rect 18923 14977 18935 14980
rect 18877 14971 18935 14977
rect 12952 14912 13584 14940
rect 12952 14900 12958 14912
rect 13630 14900 13636 14952
rect 13688 14940 13694 14952
rect 14461 14943 14519 14949
rect 14461 14940 14473 14943
rect 13688 14912 14473 14940
rect 13688 14900 13694 14912
rect 14461 14909 14473 14912
rect 14507 14909 14519 14943
rect 14642 14940 14648 14952
rect 14603 14912 14648 14940
rect 14461 14903 14519 14909
rect 14642 14900 14648 14912
rect 14700 14900 14706 14952
rect 16114 14900 16120 14952
rect 16172 14940 16178 14952
rect 19058 14940 19064 14952
rect 16172 14912 19064 14940
rect 16172 14900 16178 14912
rect 19058 14900 19064 14912
rect 19116 14900 19122 14952
rect 9398 14872 9404 14884
rect 2746 14844 9404 14872
rect 9398 14832 9404 14844
rect 9456 14832 9462 14884
rect 9950 14872 9956 14884
rect 9508 14844 9956 14872
rect 3602 14804 3608 14816
rect 3563 14776 3608 14804
rect 3602 14764 3608 14776
rect 3660 14764 3666 14816
rect 5445 14807 5503 14813
rect 5445 14773 5457 14807
rect 5491 14804 5503 14807
rect 9508 14804 9536 14844
rect 9950 14832 9956 14844
rect 10008 14832 10014 14884
rect 10226 14832 10232 14884
rect 10284 14872 10290 14884
rect 15838 14872 15844 14884
rect 10284 14844 15844 14872
rect 10284 14832 10290 14844
rect 15838 14832 15844 14844
rect 15896 14832 15902 14884
rect 19168 14872 19196 14980
rect 24765 14977 24777 15011
rect 24811 15008 24823 15011
rect 26421 15011 26479 15017
rect 26421 15008 26433 15011
rect 24811 14980 26433 15008
rect 24811 14977 24823 14980
rect 24765 14971 24823 14977
rect 26421 14977 26433 14980
rect 26467 14977 26479 15011
rect 27430 15008 27436 15020
rect 27391 14980 27436 15008
rect 26421 14971 26479 14977
rect 19334 14900 19340 14952
rect 19392 14940 19398 14952
rect 20809 14943 20867 14949
rect 19392 14912 20760 14940
rect 19392 14900 19398 14912
rect 19610 14872 19616 14884
rect 15948 14844 19012 14872
rect 19168 14844 19616 14872
rect 5491 14776 9536 14804
rect 9861 14807 9919 14813
rect 5491 14773 5503 14776
rect 5445 14767 5503 14773
rect 9861 14773 9873 14807
rect 9907 14804 9919 14807
rect 10042 14804 10048 14816
rect 9907 14776 10048 14804
rect 9907 14773 9919 14776
rect 9861 14767 9919 14773
rect 10042 14764 10048 14776
rect 10100 14764 10106 14816
rect 11514 14764 11520 14816
rect 11572 14804 11578 14816
rect 15948 14804 15976 14844
rect 11572 14776 15976 14804
rect 11572 14764 11578 14776
rect 16022 14764 16028 14816
rect 16080 14804 16086 14816
rect 18690 14804 18696 14816
rect 16080 14776 18696 14804
rect 16080 14764 16086 14776
rect 18690 14764 18696 14776
rect 18748 14764 18754 14816
rect 18984 14804 19012 14844
rect 19610 14832 19616 14844
rect 19668 14832 19674 14884
rect 20732 14872 20760 14912
rect 20809 14909 20821 14943
rect 20855 14940 20867 14943
rect 21082 14940 21088 14952
rect 20855 14912 21088 14940
rect 20855 14909 20867 14912
rect 20809 14903 20867 14909
rect 21082 14900 21088 14912
rect 21140 14900 21146 14952
rect 21376 14912 22876 14940
rect 21376 14881 21404 14912
rect 21361 14875 21419 14881
rect 21361 14872 21373 14875
rect 20732 14844 21373 14872
rect 21361 14841 21373 14844
rect 21407 14841 21419 14875
rect 21361 14835 21419 14841
rect 22738 14804 22744 14816
rect 18984 14776 22744 14804
rect 22738 14764 22744 14776
rect 22796 14764 22802 14816
rect 22848 14804 22876 14912
rect 22922 14900 22928 14952
rect 22980 14940 22986 14952
rect 25314 14940 25320 14952
rect 22980 14912 25320 14940
rect 22980 14900 22986 14912
rect 25314 14900 25320 14912
rect 25372 14900 25378 14952
rect 26436 14940 26464 14971
rect 27430 14968 27436 14980
rect 27488 14968 27494 15020
rect 29362 15008 29368 15020
rect 29323 14980 29368 15008
rect 29362 14968 29368 14980
rect 29420 14968 29426 15020
rect 29825 15011 29883 15017
rect 29825 14977 29837 15011
rect 29871 15008 29883 15011
rect 29871 14980 31754 15008
rect 29871 14977 29883 14980
rect 29825 14971 29883 14977
rect 26436 14912 27476 14940
rect 27448 14872 27476 14912
rect 27522 14900 27528 14952
rect 27580 14940 27586 14952
rect 29917 14943 29975 14949
rect 29917 14940 29929 14943
rect 27580 14912 29929 14940
rect 27580 14900 27586 14912
rect 29917 14909 29929 14912
rect 29963 14909 29975 14943
rect 31726 14940 31754 14980
rect 34514 14968 34520 15020
rect 34572 15008 34578 15020
rect 35345 15011 35403 15017
rect 35345 15008 35357 15011
rect 34572 14980 35357 15008
rect 34572 14968 34578 14980
rect 35345 14977 35357 14980
rect 35391 14977 35403 15011
rect 35345 14971 35403 14977
rect 37734 14968 37740 15020
rect 37792 15008 37798 15020
rect 38013 15011 38071 15017
rect 38013 15008 38025 15011
rect 37792 14980 38025 15008
rect 37792 14968 37798 14980
rect 38013 14977 38025 14980
rect 38059 14977 38071 15011
rect 38013 14971 38071 14977
rect 37090 14940 37096 14952
rect 31726 14912 37096 14940
rect 29917 14903 29975 14909
rect 37090 14900 37096 14912
rect 37148 14900 37154 14952
rect 35434 14872 35440 14884
rect 27448 14844 35440 14872
rect 35434 14832 35440 14844
rect 35492 14832 35498 14884
rect 23566 14804 23572 14816
rect 22848 14776 23572 14804
rect 23566 14764 23572 14776
rect 23624 14764 23630 14816
rect 28994 14764 29000 14816
rect 29052 14804 29058 14816
rect 29181 14807 29239 14813
rect 29181 14804 29193 14807
rect 29052 14776 29193 14804
rect 29052 14764 29058 14776
rect 29181 14773 29193 14776
rect 29227 14773 29239 14807
rect 29181 14767 29239 14773
rect 37829 14807 37887 14813
rect 37829 14773 37841 14807
rect 37875 14804 37887 14807
rect 37918 14804 37924 14816
rect 37875 14776 37924 14804
rect 37875 14773 37887 14776
rect 37829 14767 37887 14773
rect 37918 14764 37924 14776
rect 37976 14764 37982 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 3602 14560 3608 14612
rect 3660 14600 3666 14612
rect 5537 14603 5595 14609
rect 5537 14600 5549 14603
rect 3660 14572 5549 14600
rect 3660 14560 3666 14572
rect 5537 14569 5549 14572
rect 5583 14600 5595 14603
rect 11882 14600 11888 14612
rect 5583 14572 11888 14600
rect 5583 14569 5595 14572
rect 5537 14563 5595 14569
rect 11882 14560 11888 14572
rect 11940 14560 11946 14612
rect 12066 14560 12072 14612
rect 12124 14600 12130 14612
rect 20162 14600 20168 14612
rect 12124 14572 13584 14600
rect 12124 14560 12130 14572
rect 3329 14535 3387 14541
rect 3329 14501 3341 14535
rect 3375 14532 3387 14535
rect 5718 14532 5724 14544
rect 3375 14504 5724 14532
rect 3375 14501 3387 14504
rect 3329 14495 3387 14501
rect 5718 14492 5724 14504
rect 5776 14492 5782 14544
rect 9309 14535 9367 14541
rect 9309 14501 9321 14535
rect 9355 14532 9367 14535
rect 12434 14532 12440 14544
rect 9355 14504 12440 14532
rect 9355 14501 9367 14504
rect 9309 14495 9367 14501
rect 12434 14492 12440 14504
rect 12492 14492 12498 14544
rect 13556 14532 13584 14572
rect 14476 14572 20168 14600
rect 14366 14532 14372 14544
rect 13556 14504 14372 14532
rect 14366 14492 14372 14504
rect 14424 14492 14430 14544
rect 2498 14464 2504 14476
rect 2459 14436 2504 14464
rect 2498 14424 2504 14436
rect 2556 14424 2562 14476
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14464 4123 14467
rect 7006 14464 7012 14476
rect 4111 14436 7012 14464
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 7006 14424 7012 14436
rect 7064 14424 7070 14476
rect 7101 14467 7159 14473
rect 7101 14433 7113 14467
rect 7147 14464 7159 14467
rect 8570 14464 8576 14476
rect 7147 14436 8576 14464
rect 7147 14433 7159 14436
rect 7101 14427 7159 14433
rect 8570 14424 8576 14436
rect 8628 14424 8634 14476
rect 9953 14467 10011 14473
rect 9953 14464 9965 14467
rect 8680 14436 9965 14464
rect 2866 14356 2872 14408
rect 2924 14396 2930 14408
rect 3237 14399 3295 14405
rect 3237 14396 3249 14399
rect 2924 14368 3249 14396
rect 2924 14356 2930 14368
rect 3237 14365 3249 14368
rect 3283 14396 3295 14399
rect 3973 14399 4031 14405
rect 3973 14396 3985 14399
rect 3283 14368 3985 14396
rect 3283 14365 3295 14368
rect 3237 14359 3295 14365
rect 3973 14365 3985 14368
rect 4019 14396 4031 14399
rect 4893 14399 4951 14405
rect 4019 14368 4108 14396
rect 4019 14365 4031 14368
rect 3973 14359 4031 14365
rect 4080 14340 4108 14368
rect 4893 14365 4905 14399
rect 4939 14365 4951 14399
rect 4893 14359 4951 14365
rect 5077 14399 5135 14405
rect 5077 14365 5089 14399
rect 5123 14396 5135 14399
rect 5626 14396 5632 14408
rect 5123 14368 5632 14396
rect 5123 14365 5135 14368
rect 5077 14359 5135 14365
rect 2130 14328 2136 14340
rect 2091 14300 2136 14328
rect 2130 14288 2136 14300
rect 2188 14288 2194 14340
rect 2222 14288 2228 14340
rect 2280 14328 2286 14340
rect 2280 14300 2325 14328
rect 2280 14288 2286 14300
rect 4062 14288 4068 14340
rect 4120 14288 4126 14340
rect 4908 14328 4936 14359
rect 5626 14356 5632 14368
rect 5684 14356 5690 14408
rect 7558 14356 7564 14408
rect 7616 14396 7622 14408
rect 7653 14399 7711 14405
rect 7653 14396 7665 14399
rect 7616 14368 7665 14396
rect 7616 14356 7622 14368
rect 7653 14365 7665 14368
rect 7699 14365 7711 14399
rect 7653 14359 7711 14365
rect 5902 14328 5908 14340
rect 4908 14300 5908 14328
rect 5902 14288 5908 14300
rect 5960 14328 5966 14340
rect 6089 14331 6147 14337
rect 6089 14328 6101 14331
rect 5960 14300 6101 14328
rect 5960 14288 5966 14300
rect 6089 14297 6101 14300
rect 6135 14297 6147 14331
rect 6089 14291 6147 14297
rect 6178 14288 6184 14340
rect 6236 14328 6242 14340
rect 8680 14328 8708 14436
rect 9953 14433 9965 14436
rect 9999 14464 10011 14467
rect 10226 14464 10232 14476
rect 9999 14436 10232 14464
rect 9999 14433 10011 14436
rect 9953 14427 10011 14433
rect 10226 14424 10232 14436
rect 10284 14424 10290 14476
rect 10597 14467 10655 14473
rect 10597 14433 10609 14467
rect 10643 14464 10655 14467
rect 11146 14464 11152 14476
rect 10643 14436 11152 14464
rect 10643 14433 10655 14436
rect 10597 14427 10655 14433
rect 11146 14424 11152 14436
rect 11204 14464 11210 14476
rect 12066 14464 12072 14476
rect 11204 14436 12072 14464
rect 11204 14424 11210 14436
rect 12066 14424 12072 14436
rect 12124 14424 12130 14476
rect 14476 14464 14504 14572
rect 20162 14560 20168 14572
rect 20220 14600 20226 14612
rect 21174 14600 21180 14612
rect 20220 14572 21180 14600
rect 20220 14560 20226 14572
rect 21174 14560 21180 14572
rect 21232 14560 21238 14612
rect 21358 14560 21364 14612
rect 21416 14600 21422 14612
rect 21910 14600 21916 14612
rect 21416 14572 21916 14600
rect 21416 14560 21422 14572
rect 21910 14560 21916 14572
rect 21968 14600 21974 14612
rect 26050 14600 26056 14612
rect 21968 14572 26056 14600
rect 21968 14560 21974 14572
rect 26050 14560 26056 14572
rect 26108 14560 26114 14612
rect 15838 14492 15844 14544
rect 15896 14532 15902 14544
rect 15896 14504 21220 14532
rect 15896 14492 15902 14504
rect 13004 14436 14504 14464
rect 14553 14467 14611 14473
rect 8938 14356 8944 14408
rect 8996 14396 9002 14408
rect 9217 14399 9275 14405
rect 9217 14396 9229 14399
rect 8996 14368 9229 14396
rect 8996 14356 9002 14368
rect 9217 14365 9229 14368
rect 9263 14365 9275 14399
rect 13004 14396 13032 14436
rect 14553 14433 14565 14467
rect 14599 14464 14611 14467
rect 15010 14464 15016 14476
rect 14599 14436 15016 14464
rect 14599 14433 14611 14436
rect 14553 14427 14611 14433
rect 15010 14424 15016 14436
rect 15068 14424 15074 14476
rect 16022 14464 16028 14476
rect 15856 14436 16028 14464
rect 9217 14359 9275 14365
rect 12728 14368 13032 14396
rect 6236 14300 6281 14328
rect 6380 14300 8708 14328
rect 6236 14288 6242 14300
rect 5166 14220 5172 14272
rect 5224 14260 5230 14272
rect 5442 14260 5448 14272
rect 5224 14232 5448 14260
rect 5224 14220 5230 14232
rect 5442 14220 5448 14232
rect 5500 14260 5506 14272
rect 6380 14260 6408 14300
rect 10042 14288 10048 14340
rect 10100 14328 10106 14340
rect 10100 14300 10145 14328
rect 10100 14288 10106 14300
rect 11054 14288 11060 14340
rect 11112 14328 11118 14340
rect 11885 14331 11943 14337
rect 11885 14328 11897 14331
rect 11112 14300 11897 14328
rect 11112 14288 11118 14300
rect 11885 14297 11897 14300
rect 11931 14297 11943 14331
rect 11885 14291 11943 14297
rect 11974 14288 11980 14340
rect 12032 14328 12038 14340
rect 12728 14328 12756 14368
rect 13078 14356 13084 14408
rect 13136 14396 13142 14408
rect 13541 14399 13599 14405
rect 13541 14396 13553 14399
rect 13136 14368 13553 14396
rect 13136 14356 13142 14368
rect 13541 14365 13553 14368
rect 13587 14365 13599 14399
rect 13541 14359 13599 14365
rect 12894 14328 12900 14340
rect 12032 14300 12077 14328
rect 12360 14300 12756 14328
rect 12855 14300 12900 14328
rect 12032 14288 12038 14300
rect 5500 14232 6408 14260
rect 5500 14220 5506 14232
rect 7650 14220 7656 14272
rect 7708 14260 7714 14272
rect 7745 14263 7803 14269
rect 7745 14260 7757 14263
rect 7708 14232 7757 14260
rect 7708 14220 7714 14232
rect 7745 14229 7757 14232
rect 7791 14229 7803 14263
rect 7745 14223 7803 14229
rect 7834 14220 7840 14272
rect 7892 14260 7898 14272
rect 12360 14260 12388 14300
rect 12894 14288 12900 14300
rect 12952 14288 12958 14340
rect 14645 14331 14703 14337
rect 14645 14328 14657 14331
rect 13004 14300 14657 14328
rect 7892 14232 12388 14260
rect 7892 14220 7898 14232
rect 12434 14220 12440 14272
rect 12492 14260 12498 14272
rect 13004 14260 13032 14300
rect 14645 14297 14657 14300
rect 14691 14297 14703 14331
rect 15194 14328 15200 14340
rect 15155 14300 15200 14328
rect 14645 14291 14703 14297
rect 15194 14288 15200 14300
rect 15252 14288 15258 14340
rect 12492 14232 13032 14260
rect 12492 14220 12498 14232
rect 13262 14220 13268 14272
rect 13320 14260 13326 14272
rect 13633 14263 13691 14269
rect 13633 14260 13645 14263
rect 13320 14232 13645 14260
rect 13320 14220 13326 14232
rect 13633 14229 13645 14232
rect 13679 14229 13691 14263
rect 13633 14223 13691 14229
rect 14366 14220 14372 14272
rect 14424 14260 14430 14272
rect 15856 14260 15884 14436
rect 16022 14424 16028 14436
rect 16080 14424 16086 14476
rect 16298 14464 16304 14476
rect 16259 14436 16304 14464
rect 16298 14424 16304 14436
rect 16356 14424 16362 14476
rect 16666 14424 16672 14476
rect 16724 14464 16730 14476
rect 19242 14464 19248 14476
rect 16724 14436 19248 14464
rect 16724 14424 16730 14436
rect 19242 14424 19248 14436
rect 19300 14424 19306 14476
rect 19521 14467 19579 14473
rect 19521 14433 19533 14467
rect 19567 14464 19579 14467
rect 21082 14464 21088 14476
rect 19567 14436 21088 14464
rect 19567 14433 19579 14436
rect 19521 14427 19579 14433
rect 21082 14424 21088 14436
rect 21140 14424 21146 14476
rect 20162 14356 20168 14408
rect 20220 14396 20226 14408
rect 20220 14368 20265 14396
rect 20220 14356 20226 14368
rect 16025 14331 16083 14337
rect 16025 14297 16037 14331
rect 16071 14297 16083 14331
rect 16025 14291 16083 14297
rect 16117 14331 16175 14337
rect 16117 14297 16129 14331
rect 16163 14328 16175 14331
rect 16390 14328 16396 14340
rect 16163 14300 16396 14328
rect 16163 14297 16175 14300
rect 16117 14291 16175 14297
rect 14424 14232 15884 14260
rect 16040 14260 16068 14291
rect 16390 14288 16396 14300
rect 16448 14288 16454 14340
rect 19610 14288 19616 14340
rect 19668 14328 19674 14340
rect 21192 14328 21220 14504
rect 23400 14504 24716 14532
rect 23400 14473 23428 14504
rect 23385 14467 23443 14473
rect 23385 14433 23397 14467
rect 23431 14433 23443 14467
rect 23385 14427 23443 14433
rect 23566 14424 23572 14476
rect 23624 14464 23630 14476
rect 24688 14473 24716 14504
rect 26142 14492 26148 14544
rect 26200 14532 26206 14544
rect 26200 14504 30604 14532
rect 26200 14492 26206 14504
rect 23661 14467 23719 14473
rect 23661 14464 23673 14467
rect 23624 14436 23673 14464
rect 23624 14424 23630 14436
rect 23661 14433 23673 14436
rect 23707 14433 23719 14467
rect 23661 14427 23719 14433
rect 24673 14467 24731 14473
rect 24673 14433 24685 14467
rect 24719 14464 24731 14467
rect 29178 14464 29184 14476
rect 24719 14436 29184 14464
rect 24719 14433 24731 14436
rect 24673 14427 24731 14433
rect 29178 14424 29184 14436
rect 29236 14424 29242 14476
rect 30576 14473 30604 14504
rect 30561 14467 30619 14473
rect 30561 14433 30573 14467
rect 30607 14433 30619 14467
rect 30561 14427 30619 14433
rect 28994 14396 29000 14408
rect 28955 14368 29000 14396
rect 28994 14356 29000 14368
rect 29052 14356 29058 14408
rect 31938 14396 31944 14408
rect 31899 14368 31944 14396
rect 31938 14356 31944 14368
rect 31996 14356 32002 14408
rect 38013 14399 38071 14405
rect 38013 14396 38025 14399
rect 35866 14368 38025 14396
rect 22922 14328 22928 14340
rect 19668 14300 19713 14328
rect 21192 14300 22928 14328
rect 19668 14288 19674 14300
rect 22922 14288 22928 14300
rect 22980 14288 22986 14340
rect 23477 14331 23535 14337
rect 23477 14297 23489 14331
rect 23523 14328 23535 14331
rect 23658 14328 23664 14340
rect 23523 14300 23664 14328
rect 23523 14297 23535 14300
rect 23477 14291 23535 14297
rect 23658 14288 23664 14300
rect 23716 14288 23722 14340
rect 24765 14331 24823 14337
rect 24765 14297 24777 14331
rect 24811 14297 24823 14331
rect 24765 14291 24823 14297
rect 21266 14260 21272 14272
rect 16040 14232 21272 14260
rect 14424 14220 14430 14232
rect 21266 14220 21272 14232
rect 21324 14220 21330 14272
rect 23290 14220 23296 14272
rect 23348 14260 23354 14272
rect 24780 14260 24808 14291
rect 25590 14288 25596 14340
rect 25648 14328 25654 14340
rect 25685 14331 25743 14337
rect 25685 14328 25697 14331
rect 25648 14300 25697 14328
rect 25648 14288 25654 14300
rect 25685 14297 25697 14300
rect 25731 14297 25743 14331
rect 30282 14328 30288 14340
rect 30243 14300 30288 14328
rect 25685 14291 25743 14297
rect 30282 14288 30288 14300
rect 30340 14288 30346 14340
rect 30374 14288 30380 14340
rect 30432 14328 30438 14340
rect 30432 14300 30477 14328
rect 30432 14288 30438 14300
rect 23348 14232 24808 14260
rect 23348 14220 23354 14232
rect 28442 14220 28448 14272
rect 28500 14260 28506 14272
rect 28813 14263 28871 14269
rect 28813 14260 28825 14263
rect 28500 14232 28825 14260
rect 28500 14220 28506 14232
rect 28813 14229 28825 14232
rect 28859 14229 28871 14263
rect 28813 14223 28871 14229
rect 31757 14263 31815 14269
rect 31757 14229 31769 14263
rect 31803 14260 31815 14263
rect 35866 14260 35894 14368
rect 38013 14365 38025 14368
rect 38059 14365 38071 14399
rect 38013 14359 38071 14365
rect 38194 14260 38200 14272
rect 31803 14232 35894 14260
rect 38155 14232 38200 14260
rect 31803 14229 31815 14232
rect 31757 14223 31815 14229
rect 38194 14220 38200 14232
rect 38252 14220 38258 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 2041 14059 2099 14065
rect 2041 14025 2053 14059
rect 2087 14056 2099 14059
rect 2130 14056 2136 14068
rect 2087 14028 2136 14056
rect 2087 14025 2099 14028
rect 2041 14019 2099 14025
rect 2130 14016 2136 14028
rect 2188 14016 2194 14068
rect 2961 14059 3019 14065
rect 2961 14025 2973 14059
rect 3007 14056 3019 14059
rect 3418 14056 3424 14068
rect 3007 14028 3424 14056
rect 3007 14025 3019 14028
rect 2961 14019 3019 14025
rect 3418 14016 3424 14028
rect 3476 14016 3482 14068
rect 4982 14016 4988 14068
rect 5040 14056 5046 14068
rect 5169 14059 5227 14065
rect 5169 14056 5181 14059
rect 5040 14028 5181 14056
rect 5040 14016 5046 14028
rect 5169 14025 5181 14028
rect 5215 14025 5227 14059
rect 5169 14019 5227 14025
rect 6641 14059 6699 14065
rect 6641 14025 6653 14059
rect 6687 14056 6699 14059
rect 9490 14056 9496 14068
rect 6687 14028 9496 14056
rect 6687 14025 6699 14028
rect 6641 14019 6699 14025
rect 9490 14016 9496 14028
rect 9548 14016 9554 14068
rect 16298 14056 16304 14068
rect 13372 14028 16304 14056
rect 3694 13988 3700 14000
rect 3655 13960 3700 13988
rect 3694 13948 3700 13960
rect 3752 13948 3758 14000
rect 4617 13991 4675 13997
rect 4617 13957 4629 13991
rect 4663 13988 4675 13991
rect 5442 13988 5448 14000
rect 4663 13960 5448 13988
rect 4663 13957 4675 13960
rect 4617 13951 4675 13957
rect 5442 13948 5448 13960
rect 5500 13948 5506 14000
rect 7650 13988 7656 14000
rect 7611 13960 7656 13988
rect 7650 13948 7656 13960
rect 7708 13948 7714 14000
rect 9214 13948 9220 14000
rect 9272 13988 9278 14000
rect 9272 13960 9317 13988
rect 9272 13948 9278 13960
rect 9398 13948 9404 14000
rect 9456 13988 9462 14000
rect 9766 13988 9772 14000
rect 9456 13960 9772 13988
rect 9456 13948 9462 13960
rect 9766 13948 9772 13960
rect 9824 13948 9830 14000
rect 10594 13988 10600 14000
rect 10555 13960 10600 13988
rect 10594 13948 10600 13960
rect 10652 13948 10658 14000
rect 11882 13988 11888 14000
rect 11843 13960 11888 13988
rect 11882 13948 11888 13960
rect 11940 13948 11946 14000
rect 1394 13880 1400 13932
rect 1452 13920 1458 13932
rect 1857 13923 1915 13929
rect 1857 13920 1869 13923
rect 1452 13892 1869 13920
rect 1452 13880 1458 13892
rect 1857 13889 1869 13892
rect 1903 13889 1915 13923
rect 2866 13920 2872 13932
rect 2827 13892 2872 13920
rect 1857 13883 1915 13889
rect 2866 13880 2872 13892
rect 2924 13880 2930 13932
rect 5077 13923 5135 13929
rect 5077 13889 5089 13923
rect 5123 13918 5135 13923
rect 5123 13890 5212 13918
rect 5123 13889 5135 13890
rect 5077 13883 5135 13889
rect 2958 13812 2964 13864
rect 3016 13852 3022 13864
rect 3326 13852 3332 13864
rect 3016 13824 3332 13852
rect 3016 13812 3022 13824
rect 3326 13812 3332 13824
rect 3384 13852 3390 13864
rect 3605 13855 3663 13861
rect 3605 13852 3617 13855
rect 3384 13824 3617 13852
rect 3384 13812 3390 13824
rect 3605 13821 3617 13824
rect 3651 13821 3663 13855
rect 3605 13815 3663 13821
rect 5184 13852 5212 13890
rect 6362 13880 6368 13932
rect 6420 13920 6426 13932
rect 6549 13923 6607 13929
rect 6549 13920 6561 13923
rect 6420 13892 6561 13920
rect 6420 13880 6426 13892
rect 6549 13889 6561 13892
rect 6595 13889 6607 13923
rect 6549 13883 6607 13889
rect 6730 13852 6736 13864
rect 5184 13824 6736 13852
rect 3418 13744 3424 13796
rect 3476 13784 3482 13796
rect 5184 13784 5212 13824
rect 6730 13812 6736 13824
rect 6788 13812 6794 13864
rect 7561 13855 7619 13861
rect 7561 13821 7573 13855
rect 7607 13852 7619 13855
rect 7834 13852 7840 13864
rect 7607 13824 7840 13852
rect 7607 13821 7619 13824
rect 7561 13815 7619 13821
rect 7834 13812 7840 13824
rect 7892 13812 7898 13864
rect 7929 13855 7987 13861
rect 7929 13821 7941 13855
rect 7975 13821 7987 13855
rect 9122 13852 9128 13864
rect 9083 13824 9128 13852
rect 7929 13815 7987 13821
rect 3476 13756 5212 13784
rect 7944 13784 7972 13815
rect 9122 13812 9128 13824
rect 9180 13812 9186 13864
rect 9398 13852 9404 13864
rect 9359 13824 9404 13852
rect 9398 13812 9404 13824
rect 9456 13812 9462 13864
rect 10502 13852 10508 13864
rect 10463 13824 10508 13852
rect 10502 13812 10508 13824
rect 10560 13812 10566 13864
rect 11149 13855 11207 13861
rect 11149 13821 11161 13855
rect 11195 13852 11207 13855
rect 11238 13852 11244 13864
rect 11195 13824 11244 13852
rect 11195 13821 11207 13824
rect 11149 13815 11207 13821
rect 11238 13812 11244 13824
rect 11296 13812 11302 13864
rect 11514 13812 11520 13864
rect 11572 13852 11578 13864
rect 11793 13855 11851 13861
rect 11793 13852 11805 13855
rect 11572 13824 11805 13852
rect 11572 13812 11578 13824
rect 11793 13821 11805 13824
rect 11839 13821 11851 13855
rect 12066 13852 12072 13864
rect 12027 13824 12072 13852
rect 11793 13815 11851 13821
rect 12066 13812 12072 13824
rect 12124 13812 12130 13864
rect 13372 13784 13400 14028
rect 16298 14016 16304 14028
rect 16356 14016 16362 14068
rect 20990 14056 20996 14068
rect 16408 14028 19288 14056
rect 13909 13991 13967 13997
rect 13909 13957 13921 13991
rect 13955 13988 13967 13991
rect 14090 13988 14096 14000
rect 13955 13960 14096 13988
rect 13955 13957 13967 13960
rect 13909 13951 13967 13957
rect 14090 13948 14096 13960
rect 14148 13948 14154 14000
rect 15746 13948 15752 14000
rect 15804 13988 15810 14000
rect 16408 13988 16436 14028
rect 15804 13960 16436 13988
rect 17589 13991 17647 13997
rect 15804 13948 15810 13960
rect 17589 13957 17601 13991
rect 17635 13988 17647 13991
rect 18325 13991 18383 13997
rect 18325 13988 18337 13991
rect 17635 13960 18337 13988
rect 17635 13957 17647 13960
rect 17589 13951 17647 13957
rect 18325 13957 18337 13960
rect 18371 13957 18383 13991
rect 18325 13951 18383 13957
rect 19058 13948 19064 14000
rect 19116 13948 19122 14000
rect 19260 13997 19288 14028
rect 19628 14028 20576 14056
rect 20951 14028 20996 14056
rect 19245 13991 19303 13997
rect 19245 13957 19257 13991
rect 19291 13957 19303 13991
rect 19245 13951 19303 13957
rect 14461 13923 14519 13929
rect 14461 13889 14473 13923
rect 14507 13920 14519 13923
rect 16666 13920 16672 13932
rect 14507 13892 16672 13920
rect 14507 13889 14519 13892
rect 14461 13883 14519 13889
rect 16666 13880 16672 13892
rect 16724 13880 16730 13932
rect 16853 13923 16911 13929
rect 16853 13889 16865 13923
rect 16899 13920 16911 13923
rect 17310 13920 17316 13932
rect 16899 13892 17316 13920
rect 16899 13889 16911 13892
rect 16853 13883 16911 13889
rect 17310 13880 17316 13892
rect 17368 13880 17374 13932
rect 17494 13920 17500 13932
rect 17455 13892 17500 13920
rect 17494 13880 17500 13892
rect 17552 13880 17558 13932
rect 19076 13920 19104 13948
rect 19628 13920 19656 14028
rect 19886 13988 19892 14000
rect 19847 13960 19892 13988
rect 19886 13948 19892 13960
rect 19944 13948 19950 14000
rect 20548 13988 20576 14028
rect 20990 14016 20996 14028
rect 21048 14016 21054 14068
rect 21082 14016 21088 14068
rect 21140 14056 21146 14068
rect 24029 14059 24087 14065
rect 24029 14056 24041 14059
rect 21140 14028 24041 14056
rect 21140 14016 21146 14028
rect 24029 14025 24041 14028
rect 24075 14025 24087 14059
rect 24029 14019 24087 14025
rect 30282 14016 30288 14068
rect 30340 14056 30346 14068
rect 30837 14059 30895 14065
rect 30837 14056 30849 14059
rect 30340 14028 30849 14056
rect 30340 14016 30346 14028
rect 30837 14025 30849 14028
rect 30883 14025 30895 14059
rect 30837 14019 30895 14025
rect 25958 13988 25964 14000
rect 20548 13960 20944 13988
rect 25919 13960 25964 13988
rect 20916 13929 20944 13960
rect 25958 13948 25964 13960
rect 26016 13948 26022 14000
rect 26050 13948 26056 14000
rect 26108 13988 26114 14000
rect 26513 13991 26571 13997
rect 26513 13988 26525 13991
rect 26108 13960 26525 13988
rect 26108 13948 26114 13960
rect 26513 13957 26525 13960
rect 26559 13957 26571 13991
rect 26513 13951 26571 13957
rect 28905 13991 28963 13997
rect 28905 13957 28917 13991
rect 28951 13988 28963 13991
rect 30466 13988 30472 14000
rect 28951 13960 30472 13988
rect 28951 13957 28963 13960
rect 28905 13951 28963 13957
rect 30466 13948 30472 13960
rect 30524 13948 30530 14000
rect 19076 13892 19656 13920
rect 20901 13923 20959 13929
rect 20901 13889 20913 13923
rect 20947 13920 20959 13923
rect 21542 13920 21548 13932
rect 20947 13892 21548 13920
rect 20947 13889 20959 13892
rect 20901 13883 20959 13889
rect 21542 13880 21548 13892
rect 21600 13880 21606 13932
rect 21818 13880 21824 13932
rect 21876 13920 21882 13932
rect 22002 13920 22008 13932
rect 21876 13892 22008 13920
rect 21876 13880 21882 13892
rect 22002 13880 22008 13892
rect 22060 13880 22066 13932
rect 23937 13923 23995 13929
rect 23937 13889 23949 13923
rect 23983 13920 23995 13923
rect 25222 13920 25228 13932
rect 23983 13892 25228 13920
rect 23983 13889 23995 13892
rect 23937 13883 23995 13889
rect 25222 13880 25228 13892
rect 25280 13880 25286 13932
rect 28442 13920 28448 13932
rect 28403 13892 28448 13920
rect 28442 13880 28448 13892
rect 28500 13880 28506 13932
rect 30745 13923 30803 13929
rect 30745 13889 30757 13923
rect 30791 13920 30803 13923
rect 36906 13920 36912 13932
rect 30791 13892 36912 13920
rect 30791 13889 30803 13892
rect 30745 13883 30803 13889
rect 36906 13880 36912 13892
rect 36964 13880 36970 13932
rect 13630 13812 13636 13864
rect 13688 13852 13694 13864
rect 13817 13855 13875 13861
rect 13817 13852 13829 13855
rect 13688 13824 13829 13852
rect 13688 13812 13694 13824
rect 13817 13821 13829 13824
rect 13863 13821 13875 13855
rect 13817 13815 13875 13821
rect 13906 13812 13912 13864
rect 13964 13852 13970 13864
rect 14090 13852 14096 13864
rect 13964 13824 14096 13852
rect 13964 13812 13970 13824
rect 14090 13812 14096 13824
rect 14148 13812 14154 13864
rect 16945 13855 17003 13861
rect 16945 13821 16957 13855
rect 16991 13852 17003 13855
rect 17126 13852 17132 13864
rect 16991 13824 17132 13852
rect 16991 13821 17003 13824
rect 16945 13815 17003 13821
rect 17126 13812 17132 13824
rect 17184 13812 17190 13864
rect 18233 13855 18291 13861
rect 18233 13821 18245 13855
rect 18279 13852 18291 13855
rect 19334 13852 19340 13864
rect 18279 13824 19340 13852
rect 18279 13821 18291 13824
rect 18233 13815 18291 13821
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 19797 13855 19855 13861
rect 19797 13821 19809 13855
rect 19843 13821 19855 13855
rect 19797 13815 19855 13821
rect 20441 13855 20499 13861
rect 20441 13821 20453 13855
rect 20487 13852 20499 13855
rect 22186 13852 22192 13864
rect 20487 13824 22192 13852
rect 20487 13821 20499 13824
rect 20441 13815 20499 13821
rect 7944 13756 13400 13784
rect 3476 13744 3482 13756
rect 3970 13676 3976 13728
rect 4028 13716 4034 13728
rect 7944 13716 7972 13756
rect 17494 13744 17500 13796
rect 17552 13784 17558 13796
rect 19812 13784 19840 13815
rect 22186 13812 22192 13824
rect 22244 13812 22250 13864
rect 25869 13855 25927 13861
rect 25869 13821 25881 13855
rect 25915 13852 25927 13855
rect 26510 13852 26516 13864
rect 25915 13824 26516 13852
rect 25915 13821 25927 13824
rect 25869 13815 25927 13821
rect 26510 13812 26516 13824
rect 26568 13812 26574 13864
rect 27522 13812 27528 13864
rect 27580 13852 27586 13864
rect 28261 13855 28319 13861
rect 28261 13852 28273 13855
rect 27580 13824 28273 13852
rect 27580 13812 27586 13824
rect 28261 13821 28273 13824
rect 28307 13821 28319 13855
rect 28261 13815 28319 13821
rect 17552 13756 19840 13784
rect 17552 13744 17558 13756
rect 19886 13744 19892 13796
rect 19944 13784 19950 13796
rect 22097 13787 22155 13793
rect 22097 13784 22109 13787
rect 19944 13756 22109 13784
rect 19944 13744 19950 13756
rect 22097 13753 22109 13756
rect 22143 13753 22155 13787
rect 22097 13747 22155 13753
rect 4028 13688 7972 13716
rect 4028 13676 4034 13688
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 2590 13512 2596 13524
rect 2551 13484 2596 13512
rect 2590 13472 2596 13484
rect 2648 13472 2654 13524
rect 3326 13512 3332 13524
rect 3287 13484 3332 13512
rect 3326 13472 3332 13484
rect 3384 13472 3390 13524
rect 3694 13472 3700 13524
rect 3752 13512 3758 13524
rect 4065 13515 4123 13521
rect 4065 13512 4077 13515
rect 3752 13484 4077 13512
rect 3752 13472 3758 13484
rect 4065 13481 4077 13484
rect 4111 13481 4123 13515
rect 4706 13512 4712 13524
rect 4667 13484 4712 13512
rect 4065 13475 4123 13481
rect 4706 13472 4712 13484
rect 4764 13472 4770 13524
rect 5721 13515 5779 13521
rect 5721 13481 5733 13515
rect 5767 13512 5779 13515
rect 6178 13512 6184 13524
rect 5767 13484 6184 13512
rect 5767 13481 5779 13484
rect 5721 13475 5779 13481
rect 6178 13472 6184 13484
rect 6236 13472 6242 13524
rect 8205 13515 8263 13521
rect 8205 13481 8217 13515
rect 8251 13512 8263 13515
rect 9214 13512 9220 13524
rect 8251 13484 9220 13512
rect 8251 13481 8263 13484
rect 8205 13475 8263 13481
rect 9214 13472 9220 13484
rect 9272 13472 9278 13524
rect 10781 13515 10839 13521
rect 10781 13481 10793 13515
rect 10827 13512 10839 13515
rect 11882 13512 11888 13524
rect 10827 13484 11888 13512
rect 10827 13481 10839 13484
rect 10781 13475 10839 13481
rect 11882 13472 11888 13484
rect 11940 13472 11946 13524
rect 11992 13484 16528 13512
rect 7561 13447 7619 13453
rect 7561 13413 7573 13447
rect 7607 13444 7619 13447
rect 8294 13444 8300 13456
rect 7607 13416 8300 13444
rect 7607 13413 7619 13416
rect 7561 13407 7619 13413
rect 8294 13404 8300 13416
rect 8352 13444 8358 13456
rect 9122 13444 9128 13456
rect 8352 13416 9128 13444
rect 8352 13404 8358 13416
rect 9122 13404 9128 13416
rect 9180 13404 9186 13456
rect 1857 13379 1915 13385
rect 1857 13345 1869 13379
rect 1903 13376 1915 13379
rect 11992 13376 12020 13484
rect 12342 13404 12348 13456
rect 12400 13444 12406 13456
rect 16390 13444 16396 13456
rect 12400 13416 16396 13444
rect 12400 13404 12406 13416
rect 16390 13404 16396 13416
rect 16448 13404 16454 13456
rect 16500 13444 16528 13484
rect 16666 13472 16672 13524
rect 16724 13512 16730 13524
rect 21450 13512 21456 13524
rect 16724 13484 21456 13512
rect 16724 13472 16730 13484
rect 21450 13472 21456 13484
rect 21508 13472 21514 13524
rect 22097 13515 22155 13521
rect 22097 13481 22109 13515
rect 22143 13512 22155 13515
rect 22370 13512 22376 13524
rect 22143 13484 22376 13512
rect 22143 13481 22155 13484
rect 22097 13475 22155 13481
rect 22370 13472 22376 13484
rect 22428 13472 22434 13524
rect 25958 13512 25964 13524
rect 25919 13484 25964 13512
rect 25958 13472 25964 13484
rect 26016 13472 26022 13524
rect 31938 13444 31944 13456
rect 16500 13416 31944 13444
rect 31938 13404 31944 13416
rect 31996 13404 32002 13456
rect 21453 13379 21511 13385
rect 1903 13348 12020 13376
rect 12406 13348 21404 13376
rect 1903 13345 1915 13348
rect 1857 13339 1915 13345
rect 1670 13308 1676 13320
rect 1631 13280 1676 13308
rect 1670 13268 1676 13280
rect 1728 13268 1734 13320
rect 2501 13311 2559 13317
rect 2501 13277 2513 13311
rect 2547 13277 2559 13311
rect 2501 13271 2559 13277
rect 2516 13240 2544 13271
rect 2958 13268 2964 13320
rect 3016 13308 3022 13320
rect 3234 13308 3240 13320
rect 3016 13280 3240 13308
rect 3016 13268 3022 13280
rect 3234 13268 3240 13280
rect 3292 13268 3298 13320
rect 3973 13311 4031 13317
rect 3973 13277 3985 13311
rect 4019 13308 4031 13311
rect 4154 13308 4160 13320
rect 4019 13280 4160 13308
rect 4019 13277 4031 13280
rect 3973 13271 4031 13277
rect 4154 13268 4160 13280
rect 4212 13268 4218 13320
rect 4617 13311 4675 13317
rect 4617 13277 4629 13311
rect 4663 13308 4675 13311
rect 5350 13308 5356 13320
rect 4663 13280 5356 13308
rect 4663 13277 4675 13280
rect 4617 13271 4675 13277
rect 5350 13268 5356 13280
rect 5408 13268 5414 13320
rect 5442 13268 5448 13320
rect 5500 13308 5506 13320
rect 7484 13317 7512 13348
rect 5629 13311 5687 13317
rect 5629 13308 5641 13311
rect 5500 13280 5641 13308
rect 5500 13268 5506 13280
rect 5629 13277 5641 13280
rect 5675 13277 5687 13311
rect 5629 13271 5687 13277
rect 7469 13311 7527 13317
rect 7469 13277 7481 13311
rect 7515 13277 7527 13311
rect 8110 13308 8116 13320
rect 8071 13280 8116 13308
rect 7469 13271 7527 13277
rect 8110 13268 8116 13280
rect 8168 13268 8174 13320
rect 9490 13308 9496 13320
rect 9451 13280 9496 13308
rect 9490 13268 9496 13280
rect 9548 13268 9554 13320
rect 10134 13268 10140 13320
rect 10192 13308 10198 13320
rect 10689 13311 10747 13317
rect 10689 13308 10701 13311
rect 10192 13280 10701 13308
rect 10192 13268 10198 13280
rect 10689 13277 10701 13280
rect 10735 13277 10747 13311
rect 10689 13271 10747 13277
rect 5074 13240 5080 13252
rect 2516 13212 5080 13240
rect 5074 13200 5080 13212
rect 5132 13200 5138 13252
rect 5534 13240 5540 13252
rect 5184 13212 5540 13240
rect 4154 13132 4160 13184
rect 4212 13172 4218 13184
rect 5184 13172 5212 13212
rect 5534 13200 5540 13212
rect 5592 13240 5598 13252
rect 12406 13240 12434 13348
rect 12710 13268 12716 13320
rect 12768 13308 12774 13320
rect 14274 13308 14280 13320
rect 12768 13280 14280 13308
rect 12768 13268 12774 13280
rect 14274 13268 14280 13280
rect 14332 13268 14338 13320
rect 17678 13308 17684 13320
rect 17328 13280 17684 13308
rect 5592 13212 12434 13240
rect 14737 13243 14795 13249
rect 5592 13200 5598 13212
rect 14737 13209 14749 13243
rect 14783 13209 14795 13243
rect 14737 13203 14795 13209
rect 14829 13243 14887 13249
rect 14829 13209 14841 13243
rect 14875 13240 14887 13243
rect 15562 13240 15568 13252
rect 14875 13212 15568 13240
rect 14875 13209 14887 13212
rect 14829 13203 14887 13209
rect 9306 13172 9312 13184
rect 4212 13144 5212 13172
rect 9267 13144 9312 13172
rect 4212 13132 4218 13144
rect 9306 13132 9312 13144
rect 9364 13132 9370 13184
rect 13722 13132 13728 13184
rect 13780 13172 13786 13184
rect 14752 13172 14780 13203
rect 15562 13200 15568 13212
rect 15620 13200 15626 13252
rect 15746 13240 15752 13252
rect 15707 13212 15752 13240
rect 15746 13200 15752 13212
rect 15804 13200 15810 13252
rect 16298 13240 16304 13252
rect 16259 13212 16304 13240
rect 16298 13200 16304 13212
rect 16356 13200 16362 13252
rect 16393 13243 16451 13249
rect 16393 13209 16405 13243
rect 16439 13240 16451 13243
rect 17218 13240 17224 13252
rect 16439 13212 17224 13240
rect 16439 13209 16451 13212
rect 16393 13203 16451 13209
rect 17218 13200 17224 13212
rect 17276 13200 17282 13252
rect 17328 13249 17356 13280
rect 17678 13268 17684 13280
rect 17736 13268 17742 13320
rect 21376 13317 21404 13348
rect 21453 13345 21465 13379
rect 21499 13376 21511 13379
rect 23290 13376 23296 13388
rect 21499 13348 23296 13376
rect 21499 13345 21511 13348
rect 21453 13339 21511 13345
rect 23290 13336 23296 13348
rect 23348 13336 23354 13388
rect 21361 13311 21419 13317
rect 21361 13277 21373 13311
rect 21407 13277 21419 13311
rect 21361 13271 21419 13277
rect 21910 13268 21916 13320
rect 21968 13308 21974 13320
rect 22005 13311 22063 13317
rect 22005 13308 22017 13311
rect 21968 13280 22017 13308
rect 21968 13268 21974 13280
rect 22005 13277 22017 13280
rect 22051 13308 22063 13311
rect 23382 13308 23388 13320
rect 22051 13280 22876 13308
rect 23343 13280 23388 13308
rect 22051 13277 22063 13280
rect 22005 13271 22063 13277
rect 17313 13243 17371 13249
rect 17313 13209 17325 13243
rect 17359 13209 17371 13243
rect 17313 13203 17371 13209
rect 17494 13200 17500 13252
rect 17552 13240 17558 13252
rect 18233 13243 18291 13249
rect 18233 13240 18245 13243
rect 17552 13212 18245 13240
rect 17552 13200 17558 13212
rect 18233 13209 18245 13212
rect 18279 13209 18291 13243
rect 18233 13203 18291 13209
rect 18325 13243 18383 13249
rect 18325 13209 18337 13243
rect 18371 13209 18383 13243
rect 18325 13203 18383 13209
rect 18877 13243 18935 13249
rect 18877 13209 18889 13243
rect 18923 13240 18935 13243
rect 22646 13240 22652 13252
rect 18923 13212 22652 13240
rect 18923 13209 18935 13212
rect 18877 13203 18935 13209
rect 16666 13172 16672 13184
rect 13780 13144 16672 13172
rect 13780 13132 13786 13144
rect 16666 13132 16672 13144
rect 16724 13132 16730 13184
rect 16850 13132 16856 13184
rect 16908 13172 16914 13184
rect 18340 13172 18368 13203
rect 22646 13200 22652 13212
rect 22704 13200 22710 13252
rect 22848 13240 22876 13280
rect 23382 13268 23388 13280
rect 23440 13268 23446 13320
rect 25682 13268 25688 13320
rect 25740 13308 25746 13320
rect 25869 13311 25927 13317
rect 25869 13308 25881 13311
rect 25740 13280 25881 13308
rect 25740 13268 25746 13280
rect 25869 13277 25881 13280
rect 25915 13277 25927 13311
rect 25869 13271 25927 13277
rect 25958 13268 25964 13320
rect 26016 13308 26022 13320
rect 26513 13311 26571 13317
rect 26513 13308 26525 13311
rect 26016 13280 26525 13308
rect 26016 13268 26022 13280
rect 26513 13277 26525 13280
rect 26559 13277 26571 13311
rect 26513 13271 26571 13277
rect 27890 13268 27896 13320
rect 27948 13308 27954 13320
rect 31389 13311 31447 13317
rect 31389 13308 31401 13311
rect 27948 13280 31401 13308
rect 27948 13268 27954 13280
rect 31389 13277 31401 13280
rect 31435 13277 31447 13311
rect 31389 13271 31447 13277
rect 32306 13268 32312 13320
rect 32364 13308 32370 13320
rect 38013 13311 38071 13317
rect 38013 13308 38025 13311
rect 32364 13280 38025 13308
rect 32364 13268 32370 13280
rect 38013 13277 38025 13280
rect 38059 13277 38071 13311
rect 38013 13271 38071 13277
rect 23934 13240 23940 13252
rect 22848 13212 23940 13240
rect 23934 13200 23940 13212
rect 23992 13200 23998 13252
rect 25222 13240 25228 13252
rect 25135 13212 25228 13240
rect 25222 13200 25228 13212
rect 25280 13240 25286 13252
rect 37734 13240 37740 13252
rect 25280 13212 37740 13240
rect 25280 13200 25286 13212
rect 37734 13200 37740 13212
rect 37792 13200 37798 13252
rect 16908 13144 18368 13172
rect 23477 13175 23535 13181
rect 16908 13132 16914 13144
rect 23477 13141 23489 13175
rect 23523 13172 23535 13175
rect 23750 13172 23756 13184
rect 23523 13144 23756 13172
rect 23523 13141 23535 13144
rect 23477 13135 23535 13141
rect 23750 13132 23756 13144
rect 23808 13132 23814 13184
rect 25314 13172 25320 13184
rect 25275 13144 25320 13172
rect 25314 13132 25320 13144
rect 25372 13132 25378 13184
rect 26050 13132 26056 13184
rect 26108 13172 26114 13184
rect 26605 13175 26663 13181
rect 26605 13172 26617 13175
rect 26108 13144 26617 13172
rect 26108 13132 26114 13144
rect 26605 13141 26617 13144
rect 26651 13141 26663 13175
rect 26605 13135 26663 13141
rect 31481 13175 31539 13181
rect 31481 13141 31493 13175
rect 31527 13172 31539 13175
rect 32490 13172 32496 13184
rect 31527 13144 32496 13172
rect 31527 13141 31539 13144
rect 31481 13135 31539 13141
rect 32490 13132 32496 13144
rect 32548 13132 32554 13184
rect 38194 13172 38200 13184
rect 38155 13144 38200 13172
rect 38194 13132 38200 13144
rect 38252 13132 38258 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 2869 12971 2927 12977
rect 2869 12937 2881 12971
rect 2915 12968 2927 12971
rect 3050 12968 3056 12980
rect 2915 12940 3056 12968
rect 2915 12937 2927 12940
rect 2869 12931 2927 12937
rect 3050 12928 3056 12940
rect 3108 12928 3114 12980
rect 3513 12971 3571 12977
rect 3513 12937 3525 12971
rect 3559 12968 3571 12971
rect 3786 12968 3792 12980
rect 3559 12940 3792 12968
rect 3559 12937 3571 12940
rect 3513 12931 3571 12937
rect 3786 12928 3792 12940
rect 3844 12928 3850 12980
rect 4157 12971 4215 12977
rect 4157 12937 4169 12971
rect 4203 12968 4215 12971
rect 4614 12968 4620 12980
rect 4203 12940 4620 12968
rect 4203 12937 4215 12940
rect 4157 12931 4215 12937
rect 4614 12928 4620 12940
rect 4672 12928 4678 12980
rect 5077 12971 5135 12977
rect 5077 12937 5089 12971
rect 5123 12968 5135 12971
rect 5123 12940 12434 12968
rect 5123 12937 5135 12940
rect 5077 12931 5135 12937
rect 1765 12903 1823 12909
rect 1765 12869 1777 12903
rect 1811 12900 1823 12903
rect 2130 12900 2136 12912
rect 1811 12872 2136 12900
rect 1811 12869 1823 12872
rect 1765 12863 1823 12869
rect 2130 12860 2136 12872
rect 2188 12860 2194 12912
rect 7190 12900 7196 12912
rect 7151 12872 7196 12900
rect 7190 12860 7196 12872
rect 7248 12860 7254 12912
rect 7745 12903 7803 12909
rect 7745 12869 7757 12903
rect 7791 12900 7803 12903
rect 11054 12900 11060 12912
rect 7791 12872 11060 12900
rect 7791 12869 7803 12872
rect 7745 12863 7803 12869
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12832 2835 12835
rect 2866 12832 2872 12844
rect 2823 12804 2872 12832
rect 2823 12801 2835 12804
rect 2777 12795 2835 12801
rect 2866 12792 2872 12804
rect 2924 12792 2930 12844
rect 3418 12832 3424 12844
rect 3379 12804 3424 12832
rect 3418 12792 3424 12804
rect 3476 12792 3482 12844
rect 3878 12792 3884 12844
rect 3936 12832 3942 12844
rect 4065 12835 4123 12841
rect 4065 12832 4077 12835
rect 3936 12804 4077 12832
rect 3936 12792 3942 12804
rect 4065 12801 4077 12804
rect 4111 12801 4123 12835
rect 4982 12832 4988 12844
rect 4943 12804 4988 12832
rect 4065 12795 4123 12801
rect 4982 12792 4988 12804
rect 5040 12792 5046 12844
rect 1670 12764 1676 12776
rect 1631 12736 1676 12764
rect 1670 12724 1676 12736
rect 1728 12724 1734 12776
rect 7101 12767 7159 12773
rect 7101 12733 7113 12767
rect 7147 12764 7159 12767
rect 8294 12764 8300 12776
rect 7147 12736 8300 12764
rect 7147 12733 7159 12736
rect 7101 12727 7159 12733
rect 8294 12724 8300 12736
rect 8352 12724 8358 12776
rect 2225 12699 2283 12705
rect 2225 12665 2237 12699
rect 2271 12696 2283 12699
rect 2314 12696 2320 12708
rect 2271 12668 2320 12696
rect 2271 12665 2283 12668
rect 2225 12659 2283 12665
rect 2314 12656 2320 12668
rect 2372 12696 2378 12708
rect 8404 12696 8432 12872
rect 11054 12860 11060 12872
rect 11112 12860 11118 12912
rect 12406 12900 12434 12940
rect 14642 12928 14648 12980
rect 14700 12968 14706 12980
rect 14829 12971 14887 12977
rect 14829 12968 14841 12971
rect 14700 12940 14841 12968
rect 14700 12928 14706 12940
rect 14829 12937 14841 12940
rect 14875 12937 14887 12971
rect 15562 12968 15568 12980
rect 15523 12940 15568 12968
rect 14829 12931 14887 12937
rect 15562 12928 15568 12940
rect 15620 12928 15626 12980
rect 16850 12968 16856 12980
rect 16811 12940 16856 12968
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 17218 12928 17224 12980
rect 17276 12968 17282 12980
rect 18877 12971 18935 12977
rect 18877 12968 18889 12971
rect 17276 12940 18889 12968
rect 17276 12928 17282 12940
rect 18877 12937 18889 12940
rect 18923 12937 18935 12971
rect 18877 12931 18935 12937
rect 18966 12928 18972 12980
rect 19024 12968 19030 12980
rect 25314 12968 25320 12980
rect 19024 12940 25320 12968
rect 19024 12928 19030 12940
rect 25314 12928 25320 12940
rect 25372 12928 25378 12980
rect 29178 12968 29184 12980
rect 29139 12940 29184 12968
rect 29178 12928 29184 12940
rect 29236 12928 29242 12980
rect 32306 12968 32312 12980
rect 32267 12940 32312 12968
rect 32306 12928 32312 12940
rect 32364 12928 32370 12980
rect 17773 12903 17831 12909
rect 12406 12872 17172 12900
rect 15013 12835 15071 12841
rect 15013 12801 15025 12835
rect 15059 12832 15071 12835
rect 15378 12832 15384 12844
rect 15059 12804 15384 12832
rect 15059 12801 15071 12804
rect 15013 12795 15071 12801
rect 15378 12792 15384 12804
rect 15436 12792 15442 12844
rect 15473 12835 15531 12841
rect 15473 12801 15485 12835
rect 15519 12801 15531 12835
rect 17034 12832 17040 12844
rect 16995 12804 17040 12832
rect 15473 12795 15531 12801
rect 13814 12724 13820 12776
rect 13872 12764 13878 12776
rect 15488 12764 15516 12795
rect 17034 12792 17040 12804
rect 17092 12792 17098 12844
rect 17144 12832 17172 12872
rect 17773 12869 17785 12903
rect 17819 12900 17831 12903
rect 17862 12900 17868 12912
rect 17819 12872 17868 12900
rect 17819 12869 17831 12872
rect 17773 12863 17831 12869
rect 17862 12860 17868 12872
rect 17920 12860 17926 12912
rect 22830 12900 22836 12912
rect 22112 12872 22836 12900
rect 17494 12832 17500 12844
rect 17144 12804 17500 12832
rect 17494 12792 17500 12804
rect 17552 12792 17558 12844
rect 22112 12841 22140 12872
rect 22830 12860 22836 12872
rect 22888 12860 22894 12912
rect 23750 12900 23756 12912
rect 23711 12872 23756 12900
rect 23750 12860 23756 12872
rect 23808 12860 23814 12912
rect 18785 12835 18843 12841
rect 18785 12801 18797 12835
rect 18831 12832 18843 12835
rect 20349 12835 20407 12841
rect 20349 12832 20361 12835
rect 18831 12804 20361 12832
rect 18831 12801 18843 12804
rect 18785 12795 18843 12801
rect 20349 12801 20361 12804
rect 20395 12801 20407 12835
rect 20349 12795 20407 12801
rect 22097 12835 22155 12841
rect 22097 12801 22109 12835
rect 22143 12801 22155 12835
rect 22097 12795 22155 12801
rect 13872 12736 15516 12764
rect 17681 12767 17739 12773
rect 13872 12724 13878 12736
rect 17681 12733 17693 12767
rect 17727 12764 17739 12767
rect 17862 12764 17868 12776
rect 17727 12736 17868 12764
rect 17727 12733 17739 12736
rect 17681 12727 17739 12733
rect 17862 12724 17868 12736
rect 17920 12724 17926 12776
rect 18800 12764 18828 12795
rect 22462 12792 22468 12844
rect 22520 12832 22526 12844
rect 22741 12835 22799 12841
rect 22741 12832 22753 12835
rect 22520 12804 22753 12832
rect 22520 12792 22526 12804
rect 22741 12801 22753 12804
rect 22787 12801 22799 12835
rect 22741 12795 22799 12801
rect 29089 12835 29147 12841
rect 29089 12801 29101 12835
rect 29135 12832 29147 12835
rect 32490 12832 32496 12844
rect 29135 12804 31754 12832
rect 32451 12804 32496 12832
rect 29135 12801 29147 12804
rect 29089 12795 29147 12801
rect 18156 12736 18828 12764
rect 2372 12668 8432 12696
rect 2372 12656 2378 12668
rect 16390 12656 16396 12708
rect 16448 12696 16454 12708
rect 18156 12696 18184 12736
rect 23474 12724 23480 12776
rect 23532 12764 23538 12776
rect 23661 12767 23719 12773
rect 23661 12764 23673 12767
rect 23532 12736 23673 12764
rect 23532 12724 23538 12736
rect 23661 12733 23673 12736
rect 23707 12733 23719 12767
rect 23661 12727 23719 12733
rect 23937 12767 23995 12773
rect 23937 12733 23949 12767
rect 23983 12733 23995 12767
rect 23937 12727 23995 12733
rect 16448 12668 18184 12696
rect 18233 12699 18291 12705
rect 16448 12656 16454 12668
rect 18233 12665 18245 12699
rect 18279 12665 18291 12699
rect 18233 12659 18291 12665
rect 15194 12588 15200 12640
rect 15252 12628 15258 12640
rect 18248 12628 18276 12659
rect 21634 12656 21640 12708
rect 21692 12696 21698 12708
rect 22833 12699 22891 12705
rect 22833 12696 22845 12699
rect 21692 12668 22845 12696
rect 21692 12656 21698 12668
rect 22833 12665 22845 12668
rect 22879 12665 22891 12699
rect 22833 12659 22891 12665
rect 23566 12656 23572 12708
rect 23624 12696 23630 12708
rect 23952 12696 23980 12727
rect 23624 12668 23980 12696
rect 31726 12696 31754 12804
rect 32490 12792 32496 12804
rect 32548 12792 32554 12844
rect 38286 12832 38292 12844
rect 38247 12804 38292 12832
rect 38286 12792 38292 12804
rect 38344 12792 38350 12844
rect 38105 12699 38163 12705
rect 38105 12696 38117 12699
rect 31726 12668 38117 12696
rect 23624 12656 23630 12668
rect 38105 12665 38117 12668
rect 38151 12665 38163 12699
rect 38105 12659 38163 12665
rect 15252 12600 18276 12628
rect 15252 12588 15258 12600
rect 20070 12588 20076 12640
rect 20128 12628 20134 12640
rect 20441 12631 20499 12637
rect 20441 12628 20453 12631
rect 20128 12600 20453 12628
rect 20128 12588 20134 12600
rect 20441 12597 20453 12600
rect 20487 12597 20499 12631
rect 20441 12591 20499 12597
rect 20806 12588 20812 12640
rect 20864 12628 20870 12640
rect 22189 12631 22247 12637
rect 22189 12628 22201 12631
rect 20864 12600 22201 12628
rect 20864 12588 20870 12600
rect 22189 12597 22201 12600
rect 22235 12597 22247 12631
rect 22189 12591 22247 12597
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 2406 12424 2412 12436
rect 2367 12396 2412 12424
rect 2406 12384 2412 12396
rect 2464 12384 2470 12436
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 3053 12427 3111 12433
rect 3053 12424 3065 12427
rect 2832 12396 3065 12424
rect 2832 12384 2838 12396
rect 3053 12393 3065 12396
rect 3099 12393 3111 12427
rect 3053 12387 3111 12393
rect 7009 12427 7067 12433
rect 7009 12393 7021 12427
rect 7055 12424 7067 12427
rect 7190 12424 7196 12436
rect 7055 12396 7196 12424
rect 7055 12393 7067 12396
rect 7009 12387 7067 12393
rect 7190 12384 7196 12396
rect 7248 12384 7254 12436
rect 8570 12384 8576 12436
rect 8628 12424 8634 12436
rect 8628 12396 14964 12424
rect 8628 12384 8634 12396
rect 1762 12356 1768 12368
rect 1723 12328 1768 12356
rect 1762 12316 1768 12328
rect 1820 12316 1826 12368
rect 5629 12359 5687 12365
rect 5629 12325 5641 12359
rect 5675 12356 5687 12359
rect 10594 12356 10600 12368
rect 5675 12328 10600 12356
rect 5675 12325 5687 12328
rect 5629 12319 5687 12325
rect 10594 12316 10600 12328
rect 10652 12316 10658 12368
rect 13446 12356 13452 12368
rect 11624 12328 13452 12356
rect 2406 12288 2412 12300
rect 2319 12260 2412 12288
rect 2332 12229 2360 12260
rect 2406 12248 2412 12260
rect 2464 12288 2470 12300
rect 3418 12288 3424 12300
rect 2464 12260 3424 12288
rect 2464 12248 2470 12260
rect 3418 12248 3424 12260
rect 3476 12248 3482 12300
rect 5077 12291 5135 12297
rect 5077 12257 5089 12291
rect 5123 12288 5135 12291
rect 11514 12288 11520 12300
rect 5123 12260 11520 12288
rect 5123 12257 5135 12260
rect 5077 12251 5135 12257
rect 11514 12248 11520 12260
rect 11572 12248 11578 12300
rect 1581 12223 1639 12229
rect 1581 12189 1593 12223
rect 1627 12189 1639 12223
rect 1581 12183 1639 12189
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12189 2375 12223
rect 2958 12220 2964 12232
rect 2919 12192 2964 12220
rect 2317 12183 2375 12189
rect 1596 12152 1624 12183
rect 2958 12180 2964 12192
rect 3016 12180 3022 12232
rect 5534 12220 5540 12232
rect 5495 12192 5540 12220
rect 5534 12180 5540 12192
rect 5592 12180 5598 12232
rect 6454 12180 6460 12232
rect 6512 12220 6518 12232
rect 11624 12229 11652 12328
rect 13446 12316 13452 12328
rect 13504 12316 13510 12368
rect 14936 12365 14964 12396
rect 15378 12384 15384 12436
rect 15436 12424 15442 12436
rect 15933 12427 15991 12433
rect 15933 12424 15945 12427
rect 15436 12396 15945 12424
rect 15436 12384 15442 12396
rect 15933 12393 15945 12396
rect 15979 12393 15991 12427
rect 15933 12387 15991 12393
rect 18598 12384 18604 12436
rect 18656 12424 18662 12436
rect 23750 12424 23756 12436
rect 18656 12396 23756 12424
rect 18656 12384 18662 12396
rect 23750 12384 23756 12396
rect 23808 12384 23814 12436
rect 14921 12359 14979 12365
rect 14921 12325 14933 12359
rect 14967 12356 14979 12359
rect 18414 12356 18420 12368
rect 14967 12328 18420 12356
rect 14967 12325 14979 12328
rect 14921 12319 14979 12325
rect 18414 12316 18420 12328
rect 18472 12356 18478 12368
rect 19242 12356 19248 12368
rect 18472 12328 19248 12356
rect 18472 12316 18478 12328
rect 19242 12316 19248 12328
rect 19300 12316 19306 12368
rect 24854 12356 24860 12368
rect 21008 12328 24860 12356
rect 12529 12291 12587 12297
rect 12529 12257 12541 12291
rect 12575 12288 12587 12291
rect 13814 12288 13820 12300
rect 12575 12260 13820 12288
rect 12575 12257 12587 12260
rect 12529 12251 12587 12257
rect 13814 12248 13820 12260
rect 13872 12248 13878 12300
rect 14366 12288 14372 12300
rect 14279 12260 14372 12288
rect 14366 12248 14372 12260
rect 14424 12288 14430 12300
rect 16298 12288 16304 12300
rect 14424 12260 16304 12288
rect 14424 12248 14430 12260
rect 16298 12248 16304 12260
rect 16356 12248 16362 12300
rect 19981 12291 20039 12297
rect 19981 12257 19993 12291
rect 20027 12288 20039 12291
rect 20530 12288 20536 12300
rect 20027 12260 20536 12288
rect 20027 12257 20039 12260
rect 19981 12251 20039 12257
rect 20530 12248 20536 12260
rect 20588 12248 20594 12300
rect 21008 12297 21036 12328
rect 24854 12316 24860 12328
rect 24912 12316 24918 12368
rect 20993 12291 21051 12297
rect 20993 12257 21005 12291
rect 21039 12257 21051 12291
rect 22646 12288 22652 12300
rect 22607 12260 22652 12288
rect 20993 12251 21051 12257
rect 22646 12248 22652 12260
rect 22704 12248 22710 12300
rect 23566 12248 23572 12300
rect 23624 12288 23630 12300
rect 24673 12291 24731 12297
rect 24673 12288 24685 12291
rect 23624 12260 24685 12288
rect 23624 12248 23630 12260
rect 24673 12257 24685 12260
rect 24719 12257 24731 12291
rect 24673 12251 24731 12257
rect 25317 12291 25375 12297
rect 25317 12257 25329 12291
rect 25363 12288 25375 12291
rect 27157 12291 27215 12297
rect 27157 12288 27169 12291
rect 25363 12260 27169 12288
rect 25363 12257 25375 12260
rect 25317 12251 25375 12257
rect 27157 12257 27169 12260
rect 27203 12288 27215 12291
rect 30834 12288 30840 12300
rect 27203 12260 30840 12288
rect 27203 12257 27215 12260
rect 27157 12251 27215 12257
rect 30834 12248 30840 12260
rect 30892 12248 30898 12300
rect 6917 12223 6975 12229
rect 6917 12220 6929 12223
rect 6512 12192 6929 12220
rect 6512 12180 6518 12192
rect 6917 12189 6929 12192
rect 6963 12189 6975 12223
rect 6917 12183 6975 12189
rect 11609 12223 11667 12229
rect 11609 12189 11621 12223
rect 11655 12189 11667 12223
rect 11609 12183 11667 12189
rect 11698 12180 11704 12232
rect 11756 12220 11762 12232
rect 12437 12223 12495 12229
rect 12437 12220 12449 12223
rect 11756 12192 12449 12220
rect 11756 12180 11762 12192
rect 12437 12189 12449 12192
rect 12483 12189 12495 12223
rect 12437 12183 12495 12189
rect 13081 12223 13139 12229
rect 13081 12189 13093 12223
rect 13127 12189 13139 12223
rect 16114 12220 16120 12232
rect 16075 12192 16120 12220
rect 13081 12183 13139 12189
rect 1596 12124 2774 12152
rect 2746 12084 2774 12124
rect 3786 12112 3792 12164
rect 3844 12152 3850 12164
rect 4065 12155 4123 12161
rect 4065 12152 4077 12155
rect 3844 12124 4077 12152
rect 3844 12112 3850 12124
rect 4065 12121 4077 12124
rect 4111 12121 4123 12155
rect 4065 12115 4123 12121
rect 4157 12155 4215 12161
rect 4157 12121 4169 12155
rect 4203 12152 4215 12155
rect 4614 12152 4620 12164
rect 4203 12124 4620 12152
rect 4203 12121 4215 12124
rect 4157 12115 4215 12121
rect 4614 12112 4620 12124
rect 4672 12112 4678 12164
rect 10318 12112 10324 12164
rect 10376 12152 10382 12164
rect 10376 12124 12434 12152
rect 10376 12112 10382 12124
rect 7926 12084 7932 12096
rect 2746 12056 7932 12084
rect 7926 12044 7932 12056
rect 7984 12044 7990 12096
rect 11330 12044 11336 12096
rect 11388 12084 11394 12096
rect 11701 12087 11759 12093
rect 11701 12084 11713 12087
rect 11388 12056 11713 12084
rect 11388 12044 11394 12056
rect 11701 12053 11713 12056
rect 11747 12053 11759 12087
rect 12406 12084 12434 12124
rect 13096 12084 13124 12183
rect 16114 12180 16120 12192
rect 16172 12180 16178 12232
rect 23750 12220 23756 12232
rect 23711 12192 23756 12220
rect 23750 12180 23756 12192
rect 23808 12180 23814 12232
rect 14461 12155 14519 12161
rect 14461 12121 14473 12155
rect 14507 12152 14519 12155
rect 14734 12152 14740 12164
rect 14507 12124 14740 12152
rect 14507 12121 14519 12124
rect 14461 12115 14519 12121
rect 14734 12112 14740 12124
rect 14792 12112 14798 12164
rect 15856 12124 16574 12152
rect 12406 12056 13124 12084
rect 13173 12087 13231 12093
rect 11701 12047 11759 12053
rect 13173 12053 13185 12087
rect 13219 12084 13231 12087
rect 15856 12084 15884 12124
rect 13219 12056 15884 12084
rect 16546 12084 16574 12124
rect 20070 12112 20076 12164
rect 20128 12152 20134 12164
rect 22741 12155 22799 12161
rect 20128 12124 20173 12152
rect 20128 12112 20134 12124
rect 22741 12121 22753 12155
rect 22787 12121 22799 12155
rect 22741 12115 22799 12121
rect 23293 12155 23351 12161
rect 23293 12121 23305 12155
rect 23339 12152 23351 12155
rect 24302 12152 24308 12164
rect 23339 12124 24308 12152
rect 23339 12121 23351 12124
rect 23293 12115 23351 12121
rect 17310 12084 17316 12096
rect 16546 12056 17316 12084
rect 13219 12053 13231 12056
rect 13173 12047 13231 12053
rect 17310 12044 17316 12056
rect 17368 12044 17374 12096
rect 22756 12084 22784 12115
rect 24302 12112 24308 12124
rect 24360 12112 24366 12164
rect 24762 12112 24768 12164
rect 24820 12152 24826 12164
rect 26510 12152 26516 12164
rect 24820 12124 24865 12152
rect 26471 12124 26516 12152
rect 24820 12112 24826 12124
rect 26510 12112 26516 12124
rect 26568 12112 26574 12164
rect 26605 12155 26663 12161
rect 26605 12121 26617 12155
rect 26651 12152 26663 12155
rect 26970 12152 26976 12164
rect 26651 12124 26976 12152
rect 26651 12121 26663 12124
rect 26605 12115 26663 12121
rect 26970 12112 26976 12124
rect 27028 12112 27034 12164
rect 23845 12087 23903 12093
rect 23845 12084 23857 12087
rect 22756 12056 23857 12084
rect 23845 12053 23857 12056
rect 23891 12053 23903 12087
rect 23845 12047 23903 12053
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 4341 11883 4399 11889
rect 4341 11880 4353 11883
rect 3016 11852 4353 11880
rect 3016 11840 3022 11852
rect 4341 11849 4353 11852
rect 4387 11849 4399 11883
rect 5626 11880 5632 11892
rect 5587 11852 5632 11880
rect 4341 11843 4399 11849
rect 5626 11840 5632 11852
rect 5684 11840 5690 11892
rect 7926 11880 7932 11892
rect 7887 11852 7932 11880
rect 7926 11840 7932 11852
rect 7984 11840 7990 11892
rect 14093 11883 14151 11889
rect 8128 11852 12434 11880
rect 1949 11815 2007 11821
rect 1949 11781 1961 11815
rect 1995 11812 2007 11815
rect 2314 11812 2320 11824
rect 1995 11784 2320 11812
rect 1995 11781 2007 11784
rect 1949 11775 2007 11781
rect 2314 11772 2320 11784
rect 2372 11772 2378 11824
rect 2685 11815 2743 11821
rect 2685 11781 2697 11815
rect 2731 11812 2743 11815
rect 2866 11812 2872 11824
rect 2731 11784 2872 11812
rect 2731 11781 2743 11784
rect 2685 11775 2743 11781
rect 2866 11772 2872 11784
rect 2924 11772 2930 11824
rect 6730 11812 6736 11824
rect 6691 11784 6736 11812
rect 6730 11772 6736 11784
rect 6788 11772 6794 11824
rect 7285 11815 7343 11821
rect 7285 11781 7297 11815
rect 7331 11812 7343 11815
rect 7834 11812 7840 11824
rect 7331 11784 7840 11812
rect 7331 11781 7343 11784
rect 7285 11775 7343 11781
rect 7834 11772 7840 11784
rect 7892 11772 7898 11824
rect 1857 11747 1915 11753
rect 1857 11713 1869 11747
rect 1903 11744 1915 11747
rect 2406 11744 2412 11756
rect 1903 11716 2412 11744
rect 1903 11713 1915 11716
rect 1857 11707 1915 11713
rect 2406 11704 2412 11716
rect 2464 11704 2470 11756
rect 3602 11704 3608 11756
rect 3660 11744 3666 11756
rect 4525 11747 4583 11753
rect 4525 11744 4537 11747
rect 3660 11716 4537 11744
rect 3660 11704 3666 11716
rect 4525 11713 4537 11716
rect 4571 11713 4583 11747
rect 4525 11707 4583 11713
rect 5537 11747 5595 11753
rect 5537 11713 5549 11747
rect 5583 11744 5595 11747
rect 6454 11744 6460 11756
rect 5583 11716 6460 11744
rect 5583 11713 5595 11716
rect 5537 11707 5595 11713
rect 6454 11704 6460 11716
rect 6512 11704 6518 11756
rect 8128 11753 8156 11852
rect 8757 11815 8815 11821
rect 8757 11781 8769 11815
rect 8803 11812 8815 11815
rect 9677 11815 9735 11821
rect 8803 11784 9628 11812
rect 8803 11781 8815 11784
rect 8757 11775 8815 11781
rect 8113 11747 8171 11753
rect 8113 11713 8125 11747
rect 8159 11713 8171 11747
rect 8113 11707 8171 11713
rect 2593 11679 2651 11685
rect 2593 11645 2605 11679
rect 2639 11676 2651 11679
rect 3697 11679 3755 11685
rect 3697 11676 3709 11679
rect 2639 11648 3709 11676
rect 2639 11645 2651 11648
rect 2593 11639 2651 11645
rect 3697 11645 3709 11648
rect 3743 11645 3755 11679
rect 3697 11639 3755 11645
rect 6641 11679 6699 11685
rect 6641 11645 6653 11679
rect 6687 11645 6699 11679
rect 6641 11639 6699 11645
rect 2498 11568 2504 11620
rect 2556 11608 2562 11620
rect 3145 11611 3203 11617
rect 3145 11608 3157 11611
rect 2556 11580 3157 11608
rect 2556 11568 2562 11580
rect 3145 11577 3157 11580
rect 3191 11577 3203 11611
rect 6656 11608 6684 11639
rect 6822 11636 6828 11688
rect 6880 11676 6886 11688
rect 8665 11679 8723 11685
rect 8665 11676 8677 11679
rect 6880 11648 8677 11676
rect 6880 11636 6886 11648
rect 8665 11645 8677 11648
rect 8711 11645 8723 11679
rect 9600 11676 9628 11784
rect 9677 11781 9689 11815
rect 9723 11781 9735 11815
rect 9677 11775 9735 11781
rect 9692 11744 9720 11775
rect 9766 11772 9772 11824
rect 9824 11812 9830 11824
rect 11974 11812 11980 11824
rect 9824 11784 11980 11812
rect 9824 11772 9830 11784
rect 11974 11772 11980 11784
rect 12032 11772 12038 11824
rect 12406 11812 12434 11852
rect 14093 11849 14105 11883
rect 14139 11880 14151 11883
rect 14366 11880 14372 11892
rect 14139 11852 14372 11880
rect 14139 11849 14151 11852
rect 14093 11843 14151 11849
rect 14366 11840 14372 11852
rect 14424 11840 14430 11892
rect 14734 11880 14740 11892
rect 14695 11852 14740 11880
rect 14734 11840 14740 11852
rect 14792 11840 14798 11892
rect 16853 11883 16911 11889
rect 16853 11849 16865 11883
rect 16899 11880 16911 11883
rect 17034 11880 17040 11892
rect 16899 11852 17040 11880
rect 16899 11849 16911 11852
rect 16853 11843 16911 11849
rect 17034 11840 17040 11852
rect 17092 11840 17098 11892
rect 19334 11840 19340 11892
rect 19392 11880 19398 11892
rect 19518 11880 19524 11892
rect 19392 11852 19524 11880
rect 19392 11840 19398 11852
rect 19518 11840 19524 11852
rect 19576 11840 19582 11892
rect 23290 11840 23296 11892
rect 23348 11880 23354 11892
rect 27525 11883 27583 11889
rect 27525 11880 27537 11883
rect 23348 11852 27537 11880
rect 23348 11840 23354 11852
rect 27525 11849 27537 11852
rect 27571 11849 27583 11883
rect 27525 11843 27583 11849
rect 21910 11812 21916 11824
rect 12406 11784 21916 11812
rect 21910 11772 21916 11784
rect 21968 11772 21974 11824
rect 13722 11744 13728 11756
rect 9692 11716 13728 11744
rect 13722 11704 13728 11716
rect 13780 11704 13786 11756
rect 14001 11747 14059 11753
rect 14001 11713 14013 11747
rect 14047 11713 14059 11747
rect 14001 11707 14059 11713
rect 10502 11676 10508 11688
rect 9600 11648 10508 11676
rect 8665 11639 8723 11645
rect 10502 11636 10508 11648
rect 10560 11636 10566 11688
rect 10686 11676 10692 11688
rect 10647 11648 10692 11676
rect 10686 11636 10692 11648
rect 10744 11636 10750 11688
rect 14016 11676 14044 11707
rect 14182 11704 14188 11756
rect 14240 11744 14246 11756
rect 14550 11744 14556 11756
rect 14240 11716 14556 11744
rect 14240 11704 14246 11716
rect 14550 11704 14556 11716
rect 14608 11744 14614 11756
rect 14645 11747 14703 11753
rect 14645 11744 14657 11747
rect 14608 11716 14657 11744
rect 14608 11704 14614 11716
rect 14645 11713 14657 11716
rect 14691 11713 14703 11747
rect 14645 11707 14703 11713
rect 17037 11747 17095 11753
rect 17037 11713 17049 11747
rect 17083 11744 17095 11747
rect 17218 11744 17224 11756
rect 17083 11716 17224 11744
rect 17083 11713 17095 11716
rect 17037 11707 17095 11713
rect 17218 11704 17224 11716
rect 17276 11704 17282 11756
rect 20714 11704 20720 11756
rect 20772 11744 20778 11756
rect 22005 11747 22063 11753
rect 22005 11744 22017 11747
rect 20772 11716 22017 11744
rect 20772 11704 20778 11716
rect 22005 11713 22017 11716
rect 22051 11713 22063 11747
rect 22005 11707 22063 11713
rect 27433 11747 27491 11753
rect 27433 11713 27445 11747
rect 27479 11744 27491 11747
rect 34514 11744 34520 11756
rect 27479 11716 34520 11744
rect 27479 11713 27491 11716
rect 27433 11707 27491 11713
rect 34514 11704 34520 11716
rect 34572 11704 34578 11756
rect 15654 11676 15660 11688
rect 10796 11648 15660 11676
rect 7926 11608 7932 11620
rect 6656 11580 7932 11608
rect 3145 11571 3203 11577
rect 7926 11568 7932 11580
rect 7984 11568 7990 11620
rect 5718 11500 5724 11552
rect 5776 11540 5782 11552
rect 9766 11540 9772 11552
rect 5776 11512 9772 11540
rect 5776 11500 5782 11512
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 10410 11500 10416 11552
rect 10468 11540 10474 11552
rect 10796 11540 10824 11648
rect 15654 11636 15660 11648
rect 15712 11636 15718 11688
rect 25593 11679 25651 11685
rect 25593 11645 25605 11679
rect 25639 11676 25651 11679
rect 25774 11676 25780 11688
rect 25639 11648 25780 11676
rect 25639 11645 25651 11648
rect 25593 11639 25651 11645
rect 25774 11636 25780 11648
rect 25832 11636 25838 11688
rect 28166 11676 28172 11688
rect 28127 11648 28172 11676
rect 28166 11636 28172 11648
rect 28224 11636 28230 11688
rect 28350 11676 28356 11688
rect 28311 11648 28356 11676
rect 28350 11636 28356 11648
rect 28408 11636 28414 11688
rect 11146 11568 11152 11620
rect 11204 11608 11210 11620
rect 11606 11608 11612 11620
rect 11204 11580 11612 11608
rect 11204 11568 11210 11580
rect 11606 11568 11612 11580
rect 11664 11568 11670 11620
rect 16022 11608 16028 11620
rect 12406 11580 16028 11608
rect 10468 11512 10824 11540
rect 10468 11500 10474 11512
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 12406 11540 12434 11580
rect 16022 11568 16028 11580
rect 16080 11568 16086 11620
rect 28534 11608 28540 11620
rect 28495 11580 28540 11608
rect 28534 11568 28540 11580
rect 28592 11568 28598 11620
rect 10928 11512 12434 11540
rect 10928 11500 10934 11512
rect 14182 11500 14188 11552
rect 14240 11540 14246 11552
rect 18230 11540 18236 11552
rect 14240 11512 18236 11540
rect 14240 11500 14246 11512
rect 18230 11500 18236 11512
rect 18288 11500 18294 11552
rect 22097 11543 22155 11549
rect 22097 11509 22109 11543
rect 22143 11540 22155 11543
rect 22186 11540 22192 11552
rect 22143 11512 22192 11540
rect 22143 11509 22155 11512
rect 22097 11503 22155 11509
rect 22186 11500 22192 11512
rect 22244 11500 22250 11552
rect 24210 11500 24216 11552
rect 24268 11540 24274 11552
rect 27338 11540 27344 11552
rect 24268 11512 27344 11540
rect 24268 11500 24274 11512
rect 27338 11500 27344 11512
rect 27396 11500 27402 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 1673 11339 1731 11345
rect 1673 11305 1685 11339
rect 1719 11336 1731 11339
rect 1854 11336 1860 11348
rect 1719 11308 1860 11336
rect 1719 11305 1731 11308
rect 1673 11299 1731 11305
rect 1854 11296 1860 11308
rect 1912 11296 1918 11348
rect 6822 11336 6828 11348
rect 4816 11308 6828 11336
rect 3329 11203 3387 11209
rect 3329 11169 3341 11203
rect 3375 11200 3387 11203
rect 3970 11200 3976 11212
rect 3375 11172 3976 11200
rect 3375 11169 3387 11172
rect 3329 11163 3387 11169
rect 3970 11160 3976 11172
rect 4028 11160 4034 11212
rect 4816 11209 4844 11308
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 10502 11296 10508 11348
rect 10560 11336 10566 11348
rect 11885 11339 11943 11345
rect 11885 11336 11897 11339
rect 10560 11308 11897 11336
rect 10560 11296 10566 11308
rect 11885 11305 11897 11308
rect 11931 11305 11943 11339
rect 11885 11299 11943 11305
rect 11974 11296 11980 11348
rect 12032 11336 12038 11348
rect 14182 11336 14188 11348
rect 12032 11308 14188 11336
rect 12032 11296 12038 11308
rect 14182 11296 14188 11308
rect 14240 11296 14246 11348
rect 17034 11296 17040 11348
rect 17092 11336 17098 11348
rect 22094 11336 22100 11348
rect 17092 11308 22100 11336
rect 17092 11296 17098 11308
rect 22094 11296 22100 11308
rect 22152 11296 22158 11348
rect 22649 11339 22707 11345
rect 22649 11305 22661 11339
rect 22695 11336 22707 11339
rect 26421 11339 26479 11345
rect 26421 11336 26433 11339
rect 22695 11308 26433 11336
rect 22695 11305 22707 11308
rect 22649 11299 22707 11305
rect 26421 11305 26433 11308
rect 26467 11336 26479 11339
rect 26510 11336 26516 11348
rect 26467 11308 26516 11336
rect 26467 11305 26479 11308
rect 26421 11299 26479 11305
rect 26510 11296 26516 11308
rect 26568 11296 26574 11348
rect 27338 11296 27344 11348
rect 27396 11336 27402 11348
rect 27433 11339 27491 11345
rect 27433 11336 27445 11339
rect 27396 11308 27445 11336
rect 27396 11296 27402 11308
rect 27433 11305 27445 11308
rect 27479 11305 27491 11339
rect 27433 11299 27491 11305
rect 37090 11296 37096 11348
rect 37148 11336 37154 11348
rect 38105 11339 38163 11345
rect 38105 11336 38117 11339
rect 37148 11308 38117 11336
rect 37148 11296 37154 11308
rect 38105 11305 38117 11308
rect 38151 11305 38163 11339
rect 38105 11299 38163 11305
rect 6641 11271 6699 11277
rect 6641 11237 6653 11271
rect 6687 11268 6699 11271
rect 14642 11268 14648 11280
rect 6687 11240 11468 11268
rect 6687 11237 6699 11240
rect 6641 11231 6699 11237
rect 4801 11203 4859 11209
rect 4801 11169 4813 11203
rect 4847 11169 4859 11203
rect 5166 11200 5172 11212
rect 5127 11172 5172 11200
rect 4801 11163 4859 11169
rect 5166 11160 5172 11172
rect 5224 11160 5230 11212
rect 8202 11160 8208 11212
rect 8260 11200 8266 11212
rect 10686 11200 10692 11212
rect 8260 11172 9352 11200
rect 10647 11172 10692 11200
rect 8260 11160 8266 11172
rect 1302 11092 1308 11144
rect 1360 11132 1366 11144
rect 1581 11135 1639 11141
rect 1581 11132 1593 11135
rect 1360 11104 1593 11132
rect 1360 11092 1366 11104
rect 1581 11101 1593 11104
rect 1627 11101 1639 11135
rect 1581 11095 1639 11101
rect 6086 11092 6092 11144
rect 6144 11132 6150 11144
rect 6549 11135 6607 11141
rect 6549 11132 6561 11135
rect 6144 11104 6561 11132
rect 6144 11092 6150 11104
rect 6549 11101 6561 11104
rect 6595 11101 6607 11135
rect 6549 11095 6607 11101
rect 7098 11092 7104 11144
rect 7156 11132 7162 11144
rect 7193 11135 7251 11141
rect 7193 11132 7205 11135
rect 7156 11104 7205 11132
rect 7156 11092 7162 11104
rect 7193 11101 7205 11104
rect 7239 11101 7251 11135
rect 7193 11095 7251 11101
rect 8570 11092 8576 11144
rect 8628 11132 8634 11144
rect 9324 11141 9352 11172
rect 10686 11160 10692 11172
rect 10744 11160 10750 11212
rect 11146 11200 11152 11212
rect 11107 11172 11152 11200
rect 11146 11160 11152 11172
rect 11204 11160 11210 11212
rect 9309 11135 9367 11141
rect 8628 11104 8673 11132
rect 8628 11092 8634 11104
rect 9309 11101 9321 11135
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 9858 11092 9864 11144
rect 9916 11132 9922 11144
rect 9953 11135 10011 11141
rect 9953 11132 9965 11135
rect 9916 11104 9965 11132
rect 9916 11092 9922 11104
rect 9953 11101 9965 11104
rect 9999 11101 10011 11135
rect 9953 11095 10011 11101
rect 10045 11135 10103 11141
rect 10045 11101 10057 11135
rect 10091 11132 10103 11135
rect 10502 11132 10508 11144
rect 10091 11104 10508 11132
rect 10091 11101 10103 11104
rect 10045 11095 10103 11101
rect 10502 11092 10508 11104
rect 10560 11092 10566 11144
rect 2314 11064 2320 11076
rect 2275 11036 2320 11064
rect 2314 11024 2320 11036
rect 2372 11024 2378 11076
rect 2406 11024 2412 11076
rect 2464 11064 2470 11076
rect 2464 11036 2509 11064
rect 2464 11024 2470 11036
rect 4890 11024 4896 11076
rect 4948 11064 4954 11076
rect 7285 11067 7343 11073
rect 4948 11036 4993 11064
rect 4948 11024 4954 11036
rect 7285 11033 7297 11067
rect 7331 11064 7343 11067
rect 7926 11064 7932 11076
rect 7331 11036 7788 11064
rect 7887 11036 7932 11064
rect 7331 11033 7343 11036
rect 7285 11027 7343 11033
rect 7760 10996 7788 11036
rect 7926 11024 7932 11036
rect 7984 11024 7990 11076
rect 8021 11067 8079 11073
rect 8021 11033 8033 11067
rect 8067 11033 8079 11067
rect 8021 11027 8079 11033
rect 9401 11067 9459 11073
rect 9401 11033 9413 11067
rect 9447 11064 9459 11067
rect 10781 11067 10839 11073
rect 10781 11064 10793 11067
rect 9447 11036 10793 11064
rect 9447 11033 9459 11036
rect 9401 11027 9459 11033
rect 10781 11033 10793 11036
rect 10827 11033 10839 11067
rect 11440 11064 11468 11240
rect 12820 11240 14648 11268
rect 11606 11160 11612 11212
rect 11664 11200 11670 11212
rect 12820 11200 12848 11240
rect 14642 11228 14648 11240
rect 14700 11268 14706 11280
rect 14921 11271 14979 11277
rect 14921 11268 14933 11271
rect 14700 11240 14933 11268
rect 14700 11228 14706 11240
rect 14921 11237 14933 11240
rect 14967 11237 14979 11271
rect 14921 11231 14979 11237
rect 15933 11271 15991 11277
rect 15933 11237 15945 11271
rect 15979 11268 15991 11271
rect 37826 11268 37832 11280
rect 15979 11240 37832 11268
rect 15979 11237 15991 11240
rect 15933 11231 15991 11237
rect 37826 11228 37832 11240
rect 37884 11228 37890 11280
rect 11664 11172 12848 11200
rect 14369 11203 14427 11209
rect 11664 11160 11670 11172
rect 14369 11169 14381 11203
rect 14415 11200 14427 11203
rect 17678 11200 17684 11212
rect 14415 11172 17684 11200
rect 14415 11169 14427 11172
rect 14369 11163 14427 11169
rect 17678 11160 17684 11172
rect 17736 11200 17742 11212
rect 22005 11203 22063 11209
rect 22005 11200 22017 11203
rect 17736 11172 22017 11200
rect 17736 11160 17742 11172
rect 22005 11169 22017 11172
rect 22051 11169 22063 11203
rect 22186 11200 22192 11212
rect 22147 11172 22192 11200
rect 22005 11163 22063 11169
rect 22186 11160 22192 11172
rect 22244 11160 22250 11212
rect 24673 11203 24731 11209
rect 24673 11169 24685 11203
rect 24719 11200 24731 11203
rect 25774 11200 25780 11212
rect 24719 11172 25452 11200
rect 25735 11172 25780 11200
rect 24719 11169 24731 11172
rect 24673 11163 24731 11169
rect 11793 11135 11851 11141
rect 11793 11101 11805 11135
rect 11839 11132 11851 11135
rect 12986 11132 12992 11144
rect 11839 11104 12992 11132
rect 11839 11101 11851 11104
rect 11793 11095 11851 11101
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 15654 11092 15660 11144
rect 15712 11132 15718 11144
rect 15749 11135 15807 11141
rect 15749 11132 15761 11135
rect 15712 11104 15761 11132
rect 15712 11092 15718 11104
rect 15749 11101 15761 11104
rect 15795 11101 15807 11135
rect 23198 11132 23204 11144
rect 15749 11095 15807 11101
rect 21376 11104 23204 11132
rect 14461 11067 14519 11073
rect 14461 11064 14473 11067
rect 11440 11036 14473 11064
rect 10781 11027 10839 11033
rect 14461 11033 14473 11036
rect 14507 11033 14519 11067
rect 14461 11027 14519 11033
rect 8036 10996 8064 11027
rect 17034 11024 17040 11076
rect 17092 11064 17098 11076
rect 17221 11067 17279 11073
rect 17221 11064 17233 11067
rect 17092 11036 17233 11064
rect 17092 11024 17098 11036
rect 17221 11033 17233 11036
rect 17267 11033 17279 11067
rect 17221 11027 17279 11033
rect 17310 11024 17316 11076
rect 17368 11064 17374 11076
rect 18230 11064 18236 11076
rect 17368 11036 17413 11064
rect 18143 11036 18236 11064
rect 17368 11024 17374 11036
rect 18230 11024 18236 11036
rect 18288 11064 18294 11076
rect 20530 11064 20536 11076
rect 18288 11036 20392 11064
rect 20491 11036 20536 11064
rect 18288 11024 18294 11036
rect 7760 10968 8064 10996
rect 20364 10996 20392 11036
rect 20530 11024 20536 11036
rect 20588 11024 20594 11076
rect 20625 11067 20683 11073
rect 20625 11033 20637 11067
rect 20671 11064 20683 11067
rect 20806 11064 20812 11076
rect 20671 11036 20812 11064
rect 20671 11033 20683 11036
rect 20625 11027 20683 11033
rect 20806 11024 20812 11036
rect 20864 11024 20870 11076
rect 21376 11064 21404 11104
rect 23198 11092 23204 11104
rect 23256 11092 23262 11144
rect 20916 11036 21404 11064
rect 21545 11067 21603 11073
rect 20916 10996 20944 11036
rect 21545 11033 21557 11067
rect 21591 11064 21603 11067
rect 22094 11064 22100 11076
rect 21591 11036 22100 11064
rect 21591 11033 21603 11036
rect 21545 11027 21603 11033
rect 22094 11024 22100 11036
rect 22152 11064 22158 11076
rect 23106 11064 23112 11076
rect 22152 11036 23112 11064
rect 22152 11024 22158 11036
rect 23106 11024 23112 11036
rect 23164 11024 23170 11076
rect 24762 11064 24768 11076
rect 24723 11036 24768 11064
rect 24762 11024 24768 11036
rect 24820 11024 24826 11076
rect 25314 11064 25320 11076
rect 25275 11036 25320 11064
rect 25314 11024 25320 11036
rect 25372 11024 25378 11076
rect 25424 11064 25452 11172
rect 25774 11160 25780 11172
rect 25832 11160 25838 11212
rect 28166 11200 28172 11212
rect 28127 11172 28172 11200
rect 28166 11160 28172 11172
rect 28224 11160 28230 11212
rect 25498 11092 25504 11144
rect 25556 11132 25562 11144
rect 25961 11135 26019 11141
rect 25961 11132 25973 11135
rect 25556 11104 25973 11132
rect 25556 11092 25562 11104
rect 25961 11101 25973 11104
rect 26007 11101 26019 11135
rect 25961 11095 26019 11101
rect 27246 11092 27252 11144
rect 27304 11132 27310 11144
rect 27341 11135 27399 11141
rect 27341 11132 27353 11135
rect 27304 11104 27353 11132
rect 27304 11092 27310 11104
rect 27341 11101 27353 11104
rect 27387 11101 27399 11135
rect 38286 11132 38292 11144
rect 38247 11104 38292 11132
rect 27341 11095 27399 11101
rect 38286 11092 38292 11104
rect 38344 11092 38350 11144
rect 28534 11064 28540 11076
rect 25424 11036 28540 11064
rect 28534 11024 28540 11036
rect 28592 11024 28598 11076
rect 20364 10968 20944 10996
rect 23750 10956 23756 11008
rect 23808 10996 23814 11008
rect 25406 10996 25412 11008
rect 23808 10968 25412 10996
rect 23808 10956 23814 10968
rect 25406 10956 25412 10968
rect 25464 10956 25470 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 2314 10752 2320 10804
rect 2372 10792 2378 10804
rect 2869 10795 2927 10801
rect 2869 10792 2881 10795
rect 2372 10764 2881 10792
rect 2372 10752 2378 10764
rect 2869 10761 2881 10764
rect 2915 10761 2927 10795
rect 2869 10755 2927 10761
rect 4433 10795 4491 10801
rect 4433 10761 4445 10795
rect 4479 10792 4491 10795
rect 4890 10792 4896 10804
rect 4479 10764 4896 10792
rect 4479 10761 4491 10764
rect 4433 10755 4491 10761
rect 4890 10752 4896 10764
rect 4948 10752 4954 10804
rect 5077 10795 5135 10801
rect 5077 10761 5089 10795
rect 5123 10792 5135 10795
rect 6730 10792 6736 10804
rect 5123 10764 6736 10792
rect 5123 10761 5135 10764
rect 5077 10755 5135 10761
rect 6730 10752 6736 10764
rect 6788 10752 6794 10804
rect 13906 10752 13912 10804
rect 13964 10792 13970 10804
rect 14645 10795 14703 10801
rect 14645 10792 14657 10795
rect 13964 10764 14657 10792
rect 13964 10752 13970 10764
rect 14645 10761 14657 10764
rect 14691 10761 14703 10795
rect 17678 10792 17684 10804
rect 17639 10764 17684 10792
rect 14645 10755 14703 10761
rect 17678 10752 17684 10764
rect 17736 10752 17742 10804
rect 23293 10795 23351 10801
rect 23293 10761 23305 10795
rect 23339 10761 23351 10795
rect 23293 10755 23351 10761
rect 23937 10795 23995 10801
rect 23937 10761 23949 10795
rect 23983 10792 23995 10795
rect 24762 10792 24768 10804
rect 23983 10764 24768 10792
rect 23983 10761 23995 10764
rect 23937 10755 23995 10761
rect 1854 10724 1860 10736
rect 1815 10696 1860 10724
rect 1854 10684 1860 10696
rect 1912 10684 1918 10736
rect 2406 10684 2412 10736
rect 2464 10724 2470 10736
rect 3605 10727 3663 10733
rect 3605 10724 3617 10727
rect 2464 10696 3617 10724
rect 2464 10684 2470 10696
rect 3605 10693 3617 10696
rect 3651 10693 3663 10727
rect 4798 10724 4804 10736
rect 3605 10687 3663 10693
rect 4356 10696 4804 10724
rect 3510 10656 3516 10668
rect 3471 10628 3516 10656
rect 3510 10616 3516 10628
rect 3568 10616 3574 10668
rect 4356 10665 4384 10696
rect 4798 10684 4804 10696
rect 4856 10684 4862 10736
rect 6641 10727 6699 10733
rect 6641 10693 6653 10727
rect 6687 10724 6699 10727
rect 6822 10724 6828 10736
rect 6687 10696 6828 10724
rect 6687 10693 6699 10696
rect 6641 10687 6699 10693
rect 6822 10684 6828 10696
rect 6880 10684 6886 10736
rect 12986 10684 12992 10736
rect 13044 10724 13050 10736
rect 15289 10727 15347 10733
rect 13044 10696 15240 10724
rect 13044 10684 13050 10696
rect 4341 10659 4399 10665
rect 4341 10625 4353 10659
rect 4387 10625 4399 10659
rect 4341 10619 4399 10625
rect 4706 10616 4712 10668
rect 4764 10656 4770 10668
rect 4985 10659 5043 10665
rect 4985 10656 4997 10659
rect 4764 10628 4997 10656
rect 4764 10616 4770 10628
rect 4985 10625 4997 10628
rect 5031 10625 5043 10659
rect 5626 10656 5632 10668
rect 5587 10628 5632 10656
rect 4985 10619 5043 10625
rect 5626 10616 5632 10628
rect 5684 10616 5690 10668
rect 6546 10656 6552 10668
rect 6507 10628 6552 10656
rect 6546 10616 6552 10628
rect 6604 10616 6610 10668
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10656 11759 10659
rect 13538 10656 13544 10668
rect 11747 10628 13544 10656
rect 11747 10625 11759 10628
rect 11701 10619 11759 10625
rect 13538 10616 13544 10628
rect 13596 10616 13602 10668
rect 14550 10656 14556 10668
rect 14511 10628 14556 10656
rect 14550 10616 14556 10628
rect 14608 10616 14614 10668
rect 15212 10665 15240 10696
rect 15289 10693 15301 10727
rect 15335 10724 15347 10727
rect 19153 10727 19211 10733
rect 19153 10724 19165 10727
rect 15335 10696 19165 10724
rect 15335 10693 15347 10696
rect 15289 10687 15347 10693
rect 19153 10693 19165 10696
rect 19199 10693 19211 10727
rect 23308 10724 23336 10755
rect 24762 10752 24768 10764
rect 24820 10752 24826 10804
rect 25866 10792 25872 10804
rect 25148 10764 25872 10792
rect 25148 10724 25176 10764
rect 25866 10752 25872 10764
rect 25924 10752 25930 10804
rect 27341 10795 27399 10801
rect 27341 10761 27353 10795
rect 27387 10761 27399 10795
rect 27341 10755 27399 10761
rect 28169 10795 28227 10801
rect 28169 10761 28181 10795
rect 28215 10792 28227 10795
rect 28350 10792 28356 10804
rect 28215 10764 28356 10792
rect 28215 10761 28227 10764
rect 28169 10755 28227 10761
rect 23308 10696 24164 10724
rect 19153 10687 19211 10693
rect 15197 10659 15255 10665
rect 15197 10625 15209 10659
rect 15243 10625 15255 10659
rect 17589 10659 17647 10665
rect 17589 10656 17601 10659
rect 15197 10619 15255 10625
rect 16546 10628 17601 10656
rect 1765 10591 1823 10597
rect 1765 10557 1777 10591
rect 1811 10557 1823 10591
rect 1765 10551 1823 10557
rect 2409 10591 2467 10597
rect 2409 10557 2421 10591
rect 2455 10588 2467 10591
rect 2498 10588 2504 10600
rect 2455 10560 2504 10588
rect 2455 10557 2467 10560
rect 2409 10551 2467 10557
rect 1780 10520 1808 10551
rect 2498 10548 2504 10560
rect 2556 10548 2562 10600
rect 5350 10548 5356 10600
rect 5408 10588 5414 10600
rect 16546 10588 16574 10628
rect 17589 10625 17601 10628
rect 17635 10656 17647 10659
rect 18417 10659 18475 10665
rect 17635 10628 18368 10656
rect 17635 10625 17647 10628
rect 17589 10619 17647 10625
rect 5408 10560 16574 10588
rect 5408 10548 5414 10560
rect 3602 10520 3608 10532
rect 1780 10492 3608 10520
rect 3602 10480 3608 10492
rect 3660 10480 3666 10532
rect 3234 10412 3240 10464
rect 3292 10452 3298 10464
rect 5721 10455 5779 10461
rect 5721 10452 5733 10455
rect 3292 10424 5733 10452
rect 3292 10412 3298 10424
rect 5721 10421 5733 10424
rect 5767 10421 5779 10455
rect 5721 10415 5779 10421
rect 11793 10455 11851 10461
rect 11793 10421 11805 10455
rect 11839 10452 11851 10455
rect 11882 10452 11888 10464
rect 11839 10424 11888 10452
rect 11839 10421 11851 10424
rect 11793 10415 11851 10421
rect 11882 10412 11888 10424
rect 11940 10412 11946 10464
rect 17770 10412 17776 10464
rect 17828 10452 17834 10464
rect 18233 10455 18291 10461
rect 18233 10452 18245 10455
rect 17828 10424 18245 10452
rect 17828 10412 17834 10424
rect 18233 10421 18245 10424
rect 18279 10421 18291 10455
rect 18340 10452 18368 10628
rect 18417 10625 18429 10659
rect 18463 10656 18475 10659
rect 18690 10656 18696 10668
rect 18463 10628 18696 10656
rect 18463 10625 18475 10628
rect 18417 10619 18475 10625
rect 18690 10616 18696 10628
rect 18748 10616 18754 10668
rect 20714 10656 20720 10668
rect 20675 10628 20720 10656
rect 20714 10616 20720 10628
rect 20772 10616 20778 10668
rect 22002 10656 22008 10668
rect 21963 10628 22008 10656
rect 22002 10616 22008 10628
rect 22060 10616 22066 10668
rect 22649 10659 22707 10665
rect 22649 10625 22661 10659
rect 22695 10625 22707 10659
rect 23474 10656 23480 10668
rect 23435 10628 23480 10656
rect 22649 10619 22707 10625
rect 19058 10588 19064 10600
rect 19019 10560 19064 10588
rect 19058 10548 19064 10560
rect 19116 10548 19122 10600
rect 19426 10588 19432 10600
rect 19387 10560 19432 10588
rect 19426 10548 19432 10560
rect 19484 10548 19490 10600
rect 22664 10588 22692 10619
rect 23474 10616 23480 10628
rect 23532 10616 23538 10668
rect 24136 10665 24164 10696
rect 24228 10696 25176 10724
rect 24121 10659 24179 10665
rect 24121 10625 24133 10659
rect 24167 10625 24179 10659
rect 24121 10619 24179 10625
rect 24228 10588 24256 10696
rect 25222 10684 25228 10736
rect 25280 10724 25286 10736
rect 26053 10727 26111 10733
rect 26053 10724 26065 10727
rect 25280 10696 26065 10724
rect 25280 10684 25286 10696
rect 26053 10693 26065 10696
rect 26099 10693 26111 10727
rect 27356 10724 27384 10755
rect 28350 10752 28356 10764
rect 28408 10752 28414 10804
rect 27356 10696 28396 10724
rect 26053 10687 26111 10693
rect 24762 10656 24768 10668
rect 24723 10628 24768 10656
rect 24762 10616 24768 10628
rect 24820 10616 24826 10668
rect 25406 10656 25412 10668
rect 25367 10628 25412 10656
rect 25406 10616 25412 10628
rect 25464 10616 25470 10668
rect 27338 10616 27344 10668
rect 27396 10656 27402 10668
rect 28368 10665 28396 10696
rect 27525 10659 27583 10665
rect 27525 10656 27537 10659
rect 27396 10628 27537 10656
rect 27396 10616 27402 10628
rect 27525 10625 27537 10628
rect 27571 10625 27583 10659
rect 27525 10619 27583 10625
rect 28353 10659 28411 10665
rect 28353 10625 28365 10659
rect 28399 10625 28411 10659
rect 28353 10619 28411 10625
rect 22664 10560 24256 10588
rect 24302 10548 24308 10600
rect 24360 10588 24366 10600
rect 25961 10591 26019 10597
rect 24360 10560 25636 10588
rect 24360 10548 24366 10560
rect 20714 10480 20720 10532
rect 20772 10520 20778 10532
rect 23842 10520 23848 10532
rect 20772 10492 23848 10520
rect 20772 10480 20778 10492
rect 23842 10480 23848 10492
rect 23900 10480 23906 10532
rect 24581 10523 24639 10529
rect 24581 10489 24593 10523
rect 24627 10520 24639 10523
rect 25498 10520 25504 10532
rect 24627 10492 25504 10520
rect 24627 10489 24639 10492
rect 24581 10483 24639 10489
rect 25498 10480 25504 10492
rect 25556 10480 25562 10532
rect 25608 10520 25636 10560
rect 25961 10557 25973 10591
rect 26007 10588 26019 10591
rect 26326 10588 26332 10600
rect 26007 10560 26332 10588
rect 26007 10557 26019 10560
rect 25961 10551 26019 10557
rect 26326 10548 26332 10560
rect 26384 10548 26390 10600
rect 26605 10591 26663 10597
rect 26605 10557 26617 10591
rect 26651 10588 26663 10591
rect 29914 10588 29920 10600
rect 26651 10560 29920 10588
rect 26651 10557 26663 10560
rect 26605 10551 26663 10557
rect 26620 10520 26648 10551
rect 29914 10548 29920 10560
rect 29972 10548 29978 10600
rect 25608 10492 26648 10520
rect 20070 10452 20076 10464
rect 18340 10424 20076 10452
rect 18233 10415 18291 10421
rect 20070 10412 20076 10424
rect 20128 10412 20134 10464
rect 20806 10452 20812 10464
rect 20767 10424 20812 10452
rect 20806 10412 20812 10424
rect 20864 10412 20870 10464
rect 20898 10412 20904 10464
rect 20956 10452 20962 10464
rect 22097 10455 22155 10461
rect 22097 10452 22109 10455
rect 20956 10424 22109 10452
rect 20956 10412 20962 10424
rect 22097 10421 22109 10424
rect 22143 10421 22155 10455
rect 22097 10415 22155 10421
rect 22554 10412 22560 10464
rect 22612 10452 22618 10464
rect 22741 10455 22799 10461
rect 22741 10452 22753 10455
rect 22612 10424 22753 10452
rect 22612 10412 22618 10424
rect 22741 10421 22753 10424
rect 22787 10421 22799 10455
rect 22741 10415 22799 10421
rect 25225 10455 25283 10461
rect 25225 10421 25237 10455
rect 25271 10452 25283 10455
rect 25406 10452 25412 10464
rect 25271 10424 25412 10452
rect 25271 10421 25283 10424
rect 25225 10415 25283 10421
rect 25406 10412 25412 10424
rect 25464 10412 25470 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 2133 10251 2191 10257
rect 2133 10217 2145 10251
rect 2179 10248 2191 10251
rect 2222 10248 2228 10260
rect 2179 10220 2228 10248
rect 2179 10217 2191 10220
rect 2133 10211 2191 10217
rect 2222 10208 2228 10220
rect 2280 10208 2286 10260
rect 2777 10251 2835 10257
rect 2777 10217 2789 10251
rect 2823 10248 2835 10251
rect 3142 10248 3148 10260
rect 2823 10220 3148 10248
rect 2823 10217 2835 10220
rect 2777 10211 2835 10217
rect 3142 10208 3148 10220
rect 3200 10208 3206 10260
rect 18233 10251 18291 10257
rect 18233 10217 18245 10251
rect 18279 10248 18291 10251
rect 20073 10251 20131 10257
rect 20073 10248 20085 10251
rect 18279 10220 20085 10248
rect 18279 10217 18291 10220
rect 18233 10211 18291 10217
rect 20073 10217 20085 10220
rect 20119 10248 20131 10251
rect 23566 10248 23572 10260
rect 20119 10220 23572 10248
rect 20119 10217 20131 10220
rect 20073 10211 20131 10217
rect 23566 10208 23572 10220
rect 23624 10208 23630 10260
rect 23661 10251 23719 10257
rect 23661 10217 23673 10251
rect 23707 10248 23719 10251
rect 24762 10248 24768 10260
rect 23707 10220 24768 10248
rect 23707 10217 23719 10220
rect 23661 10211 23719 10217
rect 24762 10208 24768 10220
rect 24820 10208 24826 10260
rect 25222 10248 25228 10260
rect 25183 10220 25228 10248
rect 25222 10208 25228 10220
rect 25280 10208 25286 10260
rect 13170 10140 13176 10192
rect 13228 10180 13234 10192
rect 23474 10180 23480 10192
rect 13228 10152 23480 10180
rect 13228 10140 13234 10152
rect 3694 10112 3700 10124
rect 2700 10084 3700 10112
rect 2038 10044 2044 10056
rect 1999 10016 2044 10044
rect 2038 10004 2044 10016
rect 2096 10004 2102 10056
rect 2314 10004 2320 10056
rect 2372 10044 2378 10056
rect 2700 10053 2728 10084
rect 3694 10072 3700 10084
rect 3752 10072 3758 10124
rect 14737 10115 14795 10121
rect 14737 10081 14749 10115
rect 14783 10112 14795 10115
rect 16209 10115 16267 10121
rect 16209 10112 16221 10115
rect 14783 10084 16221 10112
rect 14783 10081 14795 10084
rect 14737 10075 14795 10081
rect 16209 10081 16221 10084
rect 16255 10081 16267 10115
rect 17770 10112 17776 10124
rect 17731 10084 17776 10112
rect 16209 10075 16267 10081
rect 17770 10072 17776 10084
rect 17828 10072 17834 10124
rect 17862 10072 17868 10124
rect 17920 10112 17926 10124
rect 19429 10115 19487 10121
rect 19429 10112 19441 10115
rect 17920 10084 19441 10112
rect 17920 10072 17926 10084
rect 19429 10081 19441 10084
rect 19475 10081 19487 10115
rect 19429 10075 19487 10081
rect 19613 10115 19671 10121
rect 19613 10081 19625 10115
rect 19659 10112 19671 10115
rect 20806 10112 20812 10124
rect 19659 10084 20812 10112
rect 19659 10081 19671 10084
rect 19613 10075 19671 10081
rect 20806 10072 20812 10084
rect 20864 10072 20870 10124
rect 2685 10047 2743 10053
rect 2685 10044 2697 10047
rect 2372 10016 2697 10044
rect 2372 10004 2378 10016
rect 2685 10013 2697 10016
rect 2731 10013 2743 10047
rect 2685 10007 2743 10013
rect 3418 10004 3424 10056
rect 3476 10044 3482 10056
rect 4157 10047 4215 10053
rect 4157 10044 4169 10047
rect 3476 10016 4169 10044
rect 3476 10004 3482 10016
rect 4157 10013 4169 10016
rect 4203 10013 4215 10047
rect 4157 10007 4215 10013
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10044 5871 10047
rect 7282 10044 7288 10056
rect 5859 10016 7288 10044
rect 5859 10013 5871 10016
rect 5813 10007 5871 10013
rect 7282 10004 7288 10016
rect 7340 10004 7346 10056
rect 17589 10047 17647 10053
rect 17589 10044 17601 10047
rect 16546 10016 17601 10044
rect 13814 9936 13820 9988
rect 13872 9976 13878 9988
rect 14829 9979 14887 9985
rect 14829 9976 14841 9979
rect 13872 9948 14841 9976
rect 13872 9936 13878 9948
rect 14829 9945 14841 9948
rect 14875 9945 14887 9979
rect 15746 9976 15752 9988
rect 15707 9948 15752 9976
rect 14829 9939 14887 9945
rect 15746 9936 15752 9948
rect 15804 9936 15810 9988
rect 3694 9868 3700 9920
rect 3752 9908 3758 9920
rect 3973 9911 4031 9917
rect 3973 9908 3985 9911
rect 3752 9880 3985 9908
rect 3752 9868 3758 9880
rect 3973 9877 3985 9880
rect 4019 9877 4031 9911
rect 5902 9908 5908 9920
rect 5815 9880 5908 9908
rect 3973 9871 4031 9877
rect 5902 9868 5908 9880
rect 5960 9908 5966 9920
rect 16546 9908 16574 10016
rect 17589 10013 17601 10016
rect 17635 10013 17647 10047
rect 17589 10007 17647 10013
rect 18877 10047 18935 10053
rect 18877 10013 18889 10047
rect 18923 10044 18935 10047
rect 20714 10044 20720 10056
rect 18923 10016 20720 10044
rect 18923 10013 18935 10016
rect 18877 10007 18935 10013
rect 17402 9936 17408 9988
rect 17460 9976 17466 9988
rect 18892 9976 18920 10007
rect 20714 10004 20720 10016
rect 20772 10004 20778 10056
rect 21376 10053 21404 10152
rect 23474 10140 23480 10152
rect 23532 10140 23538 10192
rect 22465 10115 22523 10121
rect 22465 10081 22477 10115
rect 22511 10112 22523 10115
rect 24302 10112 24308 10124
rect 22511 10084 24308 10112
rect 22511 10081 22523 10084
rect 22465 10075 22523 10081
rect 24302 10072 24308 10084
rect 24360 10072 24366 10124
rect 28626 10072 28632 10124
rect 28684 10112 28690 10124
rect 37737 10115 37795 10121
rect 37737 10112 37749 10115
rect 28684 10084 37749 10112
rect 28684 10072 28690 10084
rect 37737 10081 37749 10084
rect 37783 10081 37795 10115
rect 37737 10075 37795 10081
rect 21361 10047 21419 10053
rect 21361 10013 21373 10047
rect 21407 10013 21419 10047
rect 23842 10044 23848 10056
rect 23803 10016 23848 10044
rect 21361 10007 21419 10013
rect 23842 10004 23848 10016
rect 23900 10004 23906 10056
rect 25406 10044 25412 10056
rect 25367 10016 25412 10044
rect 25406 10004 25412 10016
rect 25464 10004 25470 10056
rect 37182 10004 37188 10056
rect 37240 10044 37246 10056
rect 37461 10047 37519 10053
rect 37461 10044 37473 10047
rect 37240 10016 37473 10044
rect 37240 10004 37246 10016
rect 37461 10013 37473 10016
rect 37507 10013 37519 10047
rect 37461 10007 37519 10013
rect 17460 9948 18920 9976
rect 17460 9936 17466 9948
rect 19242 9936 19248 9988
rect 19300 9976 19306 9988
rect 19300 9948 21588 9976
rect 19300 9936 19306 9948
rect 18690 9908 18696 9920
rect 5960 9880 16574 9908
rect 18651 9880 18696 9908
rect 5960 9868 5966 9880
rect 18690 9868 18696 9880
rect 18748 9868 18754 9920
rect 20714 9868 20720 9920
rect 20772 9908 20778 9920
rect 21453 9911 21511 9917
rect 21453 9908 21465 9911
rect 20772 9880 21465 9908
rect 20772 9868 20778 9880
rect 21453 9877 21465 9880
rect 21499 9877 21511 9911
rect 21560 9908 21588 9948
rect 22554 9936 22560 9988
rect 22612 9976 22618 9988
rect 23109 9979 23167 9985
rect 22612 9948 22657 9976
rect 22612 9936 22618 9948
rect 23109 9945 23121 9979
rect 23155 9945 23167 9979
rect 23109 9939 23167 9945
rect 23124 9908 23152 9939
rect 21560 9880 23152 9908
rect 21453 9871 21511 9877
rect 25682 9868 25688 9920
rect 25740 9908 25746 9920
rect 25869 9911 25927 9917
rect 25869 9908 25881 9911
rect 25740 9880 25881 9908
rect 25740 9868 25746 9880
rect 25869 9877 25881 9880
rect 25915 9877 25927 9911
rect 25869 9871 25927 9877
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 1765 9707 1823 9713
rect 1765 9673 1777 9707
rect 1811 9704 1823 9707
rect 1854 9704 1860 9716
rect 1811 9676 1860 9704
rect 1811 9673 1823 9676
rect 1765 9667 1823 9673
rect 1854 9664 1860 9676
rect 1912 9664 1918 9716
rect 18693 9707 18751 9713
rect 18693 9673 18705 9707
rect 18739 9704 18751 9707
rect 19058 9704 19064 9716
rect 18739 9676 19064 9704
rect 18739 9673 18751 9676
rect 18693 9667 18751 9673
rect 19058 9664 19064 9676
rect 19116 9664 19122 9716
rect 20898 9704 20904 9716
rect 20548 9676 20904 9704
rect 2130 9596 2136 9648
rect 2188 9636 2194 9648
rect 2409 9639 2467 9645
rect 2409 9636 2421 9639
rect 2188 9608 2421 9636
rect 2188 9596 2194 9608
rect 2409 9605 2421 9608
rect 2455 9605 2467 9639
rect 2409 9599 2467 9605
rect 2866 9596 2872 9648
rect 2924 9636 2930 9648
rect 3145 9639 3203 9645
rect 3145 9636 3157 9639
rect 2924 9608 3157 9636
rect 2924 9596 2930 9608
rect 3145 9605 3157 9608
rect 3191 9605 3203 9639
rect 3786 9636 3792 9648
rect 3747 9608 3792 9636
rect 3145 9599 3203 9605
rect 3786 9596 3792 9608
rect 3844 9596 3850 9648
rect 14734 9596 14740 9648
rect 14792 9636 14798 9648
rect 17037 9639 17095 9645
rect 17037 9636 17049 9639
rect 14792 9608 17049 9636
rect 14792 9596 14798 9608
rect 17037 9605 17049 9608
rect 17083 9605 17095 9639
rect 17037 9599 17095 9605
rect 17126 9596 17132 9648
rect 17184 9636 17190 9648
rect 17681 9639 17739 9645
rect 17184 9608 17229 9636
rect 17184 9596 17190 9608
rect 17681 9605 17693 9639
rect 17727 9636 17739 9639
rect 19426 9636 19432 9648
rect 17727 9608 19432 9636
rect 17727 9605 17739 9608
rect 17681 9599 17739 9605
rect 19426 9596 19432 9608
rect 19484 9596 19490 9648
rect 19521 9639 19579 9645
rect 19521 9605 19533 9639
rect 19567 9636 19579 9639
rect 20548 9636 20576 9676
rect 20898 9664 20904 9676
rect 20956 9664 20962 9716
rect 20714 9636 20720 9648
rect 19567 9608 20576 9636
rect 20675 9608 20720 9636
rect 19567 9605 19579 9608
rect 19521 9599 19579 9605
rect 20714 9596 20720 9608
rect 20772 9596 20778 9648
rect 24302 9596 24308 9648
rect 24360 9636 24366 9648
rect 30285 9639 30343 9645
rect 30285 9636 30297 9639
rect 24360 9608 30297 9636
rect 24360 9596 24366 9608
rect 30285 9605 30297 9608
rect 30331 9605 30343 9639
rect 30285 9599 30343 9605
rect 1118 9528 1124 9580
rect 1176 9568 1182 9580
rect 1673 9571 1731 9577
rect 1673 9568 1685 9571
rect 1176 9540 1685 9568
rect 1176 9528 1182 9540
rect 1673 9537 1685 9540
rect 1719 9537 1731 9571
rect 2314 9568 2320 9580
rect 2275 9540 2320 9568
rect 1673 9531 1731 9537
rect 2314 9528 2320 9540
rect 2372 9528 2378 9580
rect 3050 9568 3056 9580
rect 3011 9540 3056 9568
rect 3050 9528 3056 9540
rect 3108 9528 3114 9580
rect 3694 9568 3700 9580
rect 3655 9540 3700 9568
rect 3694 9528 3700 9540
rect 3752 9528 3758 9580
rect 5626 9528 5632 9580
rect 5684 9568 5690 9580
rect 7101 9571 7159 9577
rect 7101 9568 7113 9571
rect 5684 9540 7113 9568
rect 5684 9528 5690 9540
rect 7101 9537 7113 9540
rect 7147 9537 7159 9571
rect 7101 9531 7159 9537
rect 13998 9528 14004 9580
rect 14056 9568 14062 9580
rect 14185 9571 14243 9577
rect 14185 9568 14197 9571
rect 14056 9540 14197 9568
rect 14056 9528 14062 9540
rect 14185 9537 14197 9540
rect 14231 9568 14243 9571
rect 14458 9568 14464 9580
rect 14231 9540 14464 9568
rect 14231 9537 14243 9540
rect 14185 9531 14243 9537
rect 14458 9528 14464 9540
rect 14516 9568 14522 9580
rect 18598 9568 18604 9580
rect 14516 9540 15608 9568
rect 18511 9540 18604 9568
rect 14516 9528 14522 9540
rect 7193 9503 7251 9509
rect 7193 9469 7205 9503
rect 7239 9500 7251 9503
rect 7926 9500 7932 9512
rect 7239 9472 7932 9500
rect 7239 9469 7251 9472
rect 7193 9463 7251 9469
rect 7926 9460 7932 9472
rect 7984 9500 7990 9512
rect 15289 9503 15347 9509
rect 15289 9500 15301 9503
rect 7984 9472 15301 9500
rect 7984 9460 7990 9472
rect 15289 9469 15301 9472
rect 15335 9469 15347 9503
rect 15289 9463 15347 9469
rect 15378 9460 15384 9512
rect 15436 9500 15442 9512
rect 15473 9503 15531 9509
rect 15473 9500 15485 9503
rect 15436 9472 15485 9500
rect 15436 9460 15442 9472
rect 15473 9469 15485 9472
rect 15519 9469 15531 9503
rect 15580 9500 15608 9540
rect 18598 9528 18604 9540
rect 18656 9568 18662 9580
rect 20073 9571 20131 9577
rect 18656 9540 19012 9568
rect 18656 9528 18662 9540
rect 17678 9500 17684 9512
rect 15580 9472 17684 9500
rect 15473 9463 15531 9469
rect 17678 9460 17684 9472
rect 17736 9460 17742 9512
rect 18984 9432 19012 9540
rect 20073 9537 20085 9571
rect 20119 9568 20131 9571
rect 20162 9568 20168 9580
rect 20119 9540 20168 9568
rect 20119 9537 20131 9540
rect 20073 9531 20131 9537
rect 20162 9528 20168 9540
rect 20220 9528 20226 9580
rect 25222 9568 25228 9580
rect 25183 9540 25228 9568
rect 25222 9528 25228 9540
rect 25280 9528 25286 9580
rect 25682 9568 25688 9580
rect 25643 9540 25688 9568
rect 25682 9528 25688 9540
rect 25740 9528 25746 9580
rect 26326 9568 26332 9580
rect 26287 9540 26332 9568
rect 26326 9528 26332 9540
rect 26384 9528 26390 9580
rect 27157 9571 27215 9577
rect 27157 9537 27169 9571
rect 27203 9568 27215 9571
rect 27706 9568 27712 9580
rect 27203 9540 27712 9568
rect 27203 9537 27215 9540
rect 27157 9531 27215 9537
rect 27706 9528 27712 9540
rect 27764 9528 27770 9580
rect 30193 9571 30251 9577
rect 30193 9537 30205 9571
rect 30239 9568 30251 9571
rect 30239 9540 35894 9568
rect 30239 9537 30251 9540
rect 30193 9531 30251 9537
rect 19426 9500 19432 9512
rect 19387 9472 19432 9500
rect 19426 9460 19432 9472
rect 19484 9460 19490 9512
rect 20625 9503 20683 9509
rect 20625 9500 20637 9503
rect 19812 9472 20637 9500
rect 19702 9432 19708 9444
rect 18984 9404 19708 9432
rect 19702 9392 19708 9404
rect 19760 9392 19766 9444
rect 19812 9376 19840 9472
rect 20625 9469 20637 9472
rect 20671 9469 20683 9503
rect 20625 9463 20683 9469
rect 21269 9503 21327 9509
rect 21269 9469 21281 9503
rect 21315 9500 21327 9503
rect 25314 9500 25320 9512
rect 21315 9472 25320 9500
rect 21315 9469 21327 9472
rect 21269 9463 21327 9469
rect 25314 9460 25320 9472
rect 25372 9460 25378 9512
rect 25869 9503 25927 9509
rect 25869 9469 25881 9503
rect 25915 9500 25927 9503
rect 26510 9500 26516 9512
rect 25915 9472 26516 9500
rect 25915 9469 25927 9472
rect 25869 9463 25927 9469
rect 26510 9460 26516 9472
rect 26568 9460 26574 9512
rect 27341 9503 27399 9509
rect 27341 9469 27353 9503
rect 27387 9469 27399 9503
rect 35866 9500 35894 9540
rect 37182 9500 37188 9512
rect 35866 9472 37188 9500
rect 27341 9463 27399 9469
rect 25958 9392 25964 9444
rect 26016 9432 26022 9444
rect 27356 9432 27384 9463
rect 37182 9460 37188 9472
rect 37240 9460 37246 9512
rect 26016 9404 27384 9432
rect 26016 9392 26022 9404
rect 14277 9367 14335 9373
rect 14277 9333 14289 9367
rect 14323 9364 14335 9367
rect 14458 9364 14464 9376
rect 14323 9336 14464 9364
rect 14323 9333 14335 9336
rect 14277 9327 14335 9333
rect 14458 9324 14464 9336
rect 14516 9324 14522 9376
rect 15933 9367 15991 9373
rect 15933 9333 15945 9367
rect 15979 9364 15991 9367
rect 19794 9364 19800 9376
rect 15979 9336 19800 9364
rect 15979 9333 15991 9336
rect 15933 9327 15991 9333
rect 19794 9324 19800 9336
rect 19852 9324 19858 9376
rect 25041 9367 25099 9373
rect 25041 9333 25053 9367
rect 25087 9364 25099 9367
rect 26234 9364 26240 9376
rect 25087 9336 26240 9364
rect 25087 9333 25099 9336
rect 25041 9327 25099 9333
rect 26234 9324 26240 9336
rect 26292 9324 26298 9376
rect 26326 9324 26332 9376
rect 26384 9364 26390 9376
rect 27525 9367 27583 9373
rect 27525 9364 27537 9367
rect 26384 9336 27537 9364
rect 26384 9324 26390 9336
rect 27525 9333 27537 9336
rect 27571 9333 27583 9367
rect 27525 9327 27583 9333
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 2593 9163 2651 9169
rect 2593 9129 2605 9163
rect 2639 9160 2651 9163
rect 4614 9160 4620 9172
rect 2639 9132 4620 9160
rect 2639 9129 2651 9132
rect 2593 9123 2651 9129
rect 4614 9120 4620 9132
rect 4672 9120 4678 9172
rect 17862 9160 17868 9172
rect 17823 9132 17868 9160
rect 17862 9120 17868 9132
rect 17920 9120 17926 9172
rect 19794 9160 19800 9172
rect 19755 9132 19800 9160
rect 19794 9120 19800 9132
rect 19852 9120 19858 9172
rect 25958 9160 25964 9172
rect 25919 9132 25964 9160
rect 25958 9120 25964 9132
rect 26016 9120 26022 9172
rect 26510 9160 26516 9172
rect 26471 9132 26516 9160
rect 26510 9120 26516 9132
rect 26568 9120 26574 9172
rect 2038 9092 2044 9104
rect 1999 9064 2044 9092
rect 2038 9052 2044 9064
rect 2096 9052 2102 9104
rect 3050 9052 3056 9104
rect 3108 9092 3114 9104
rect 3237 9095 3295 9101
rect 3237 9092 3249 9095
rect 3108 9064 3249 9092
rect 3108 9052 3114 9064
rect 3237 9061 3249 9064
rect 3283 9092 3295 9095
rect 9582 9092 9588 9104
rect 3283 9064 9588 9092
rect 3283 9061 3295 9064
rect 3237 9055 3295 9061
rect 9582 9052 9588 9064
rect 9640 9052 9646 9104
rect 13538 9052 13544 9104
rect 13596 9092 13602 9104
rect 14645 9095 14703 9101
rect 14645 9092 14657 9095
rect 13596 9064 14657 9092
rect 13596 9052 13602 9064
rect 14645 9061 14657 9064
rect 14691 9061 14703 9095
rect 14645 9055 14703 9061
rect 18708 9064 23796 9092
rect 4798 9024 4804 9036
rect 2516 8996 4804 9024
rect 2516 8965 2544 8996
rect 4798 8984 4804 8996
rect 4856 8984 4862 9036
rect 10962 8984 10968 9036
rect 11020 9024 11026 9036
rect 11517 9027 11575 9033
rect 11517 9024 11529 9027
rect 11020 8996 11529 9024
rect 11020 8984 11026 8996
rect 11517 8993 11529 8996
rect 11563 9024 11575 9027
rect 14277 9027 14335 9033
rect 11563 8996 14228 9024
rect 11563 8993 11575 8996
rect 11517 8987 11575 8993
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8925 2559 8959
rect 3142 8956 3148 8968
rect 3103 8928 3148 8956
rect 2501 8919 2559 8925
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 1578 8848 1584 8900
rect 1636 8888 1642 8900
rect 1857 8891 1915 8897
rect 1857 8888 1869 8891
rect 1636 8860 1869 8888
rect 1636 8848 1642 8860
rect 1857 8857 1869 8860
rect 1903 8888 1915 8891
rect 4982 8888 4988 8900
rect 1903 8860 4988 8888
rect 1903 8857 1915 8860
rect 1857 8851 1915 8857
rect 4982 8848 4988 8860
rect 5040 8848 5046 8900
rect 11238 8888 11244 8900
rect 11199 8860 11244 8888
rect 11238 8848 11244 8860
rect 11296 8848 11302 8900
rect 11330 8848 11336 8900
rect 11388 8888 11394 8900
rect 14200 8888 14228 8996
rect 14277 8993 14289 9027
rect 14323 9024 14335 9027
rect 15930 9024 15936 9036
rect 14323 8996 15424 9024
rect 15891 8996 15936 9024
rect 14323 8993 14335 8996
rect 14277 8987 14335 8993
rect 14458 8956 14464 8968
rect 14419 8928 14464 8956
rect 14458 8916 14464 8928
rect 14516 8916 14522 8968
rect 15396 8956 15424 8996
rect 15930 8984 15936 8996
rect 15988 8984 15994 9036
rect 16206 8984 16212 9036
rect 16264 9024 16270 9036
rect 18708 9024 18736 9064
rect 16264 8996 18736 9024
rect 16264 8984 16270 8996
rect 17770 8956 17776 8968
rect 15396 8928 17632 8956
rect 17731 8928 17776 8956
rect 15470 8888 15476 8900
rect 11388 8860 11433 8888
rect 14200 8860 15476 8888
rect 11388 8848 11394 8860
rect 15470 8848 15476 8860
rect 15528 8848 15534 8900
rect 15749 8891 15807 8897
rect 15749 8857 15761 8891
rect 15795 8888 15807 8891
rect 15795 8860 16574 8888
rect 15795 8857 15807 8860
rect 15749 8851 15807 8857
rect 16546 8820 16574 8860
rect 16850 8820 16856 8832
rect 16546 8792 16856 8820
rect 16850 8780 16856 8792
rect 16908 8780 16914 8832
rect 17604 8820 17632 8928
rect 17770 8916 17776 8928
rect 17828 8916 17834 8968
rect 18708 8965 18736 8996
rect 18785 9027 18843 9033
rect 18785 8993 18797 9027
rect 18831 9024 18843 9027
rect 19613 9027 19671 9033
rect 19613 9024 19625 9027
rect 18831 8996 19625 9024
rect 18831 8993 18843 8996
rect 18785 8987 18843 8993
rect 19613 8993 19625 8996
rect 19659 8993 19671 9027
rect 19613 8987 19671 8993
rect 23109 9027 23167 9033
rect 23109 8993 23121 9027
rect 23155 9024 23167 9027
rect 23290 9024 23296 9036
rect 23155 8996 23296 9024
rect 23155 8993 23167 8996
rect 23109 8987 23167 8993
rect 23290 8984 23296 8996
rect 23348 8984 23354 9036
rect 23474 9024 23480 9036
rect 23435 8996 23480 9024
rect 23474 8984 23480 8996
rect 23532 8984 23538 9036
rect 18693 8959 18751 8965
rect 18693 8925 18705 8959
rect 18739 8925 18751 8959
rect 18693 8919 18751 8925
rect 19058 8916 19064 8968
rect 19116 8956 19122 8968
rect 19429 8959 19487 8965
rect 19429 8956 19441 8959
rect 19116 8928 19441 8956
rect 19116 8916 19122 8928
rect 19429 8925 19441 8928
rect 19475 8925 19487 8959
rect 22370 8956 22376 8968
rect 19429 8919 19487 8925
rect 20456 8928 22376 8956
rect 17678 8848 17684 8900
rect 17736 8888 17742 8900
rect 20456 8888 20484 8928
rect 22370 8916 22376 8928
rect 22428 8916 22434 8968
rect 17736 8860 20484 8888
rect 23201 8891 23259 8897
rect 17736 8848 17742 8860
rect 23201 8857 23213 8891
rect 23247 8857 23259 8891
rect 23768 8888 23796 9064
rect 25222 8916 25228 8968
rect 25280 8956 25286 8968
rect 25869 8959 25927 8965
rect 25869 8956 25881 8959
rect 25280 8928 25881 8956
rect 25280 8916 25286 8928
rect 25869 8925 25881 8928
rect 25915 8925 25927 8959
rect 25869 8919 25927 8925
rect 26234 8916 26240 8968
rect 26292 8956 26298 8968
rect 26697 8959 26755 8965
rect 26697 8956 26709 8959
rect 26292 8928 26709 8956
rect 26292 8916 26298 8928
rect 26697 8925 26709 8928
rect 26743 8925 26755 8959
rect 35986 8956 35992 8968
rect 35947 8928 35992 8956
rect 26697 8919 26755 8925
rect 35986 8916 35992 8928
rect 36044 8916 36050 8968
rect 27338 8888 27344 8900
rect 23768 8860 27344 8888
rect 23201 8851 23259 8857
rect 20254 8820 20260 8832
rect 17604 8792 20260 8820
rect 20254 8780 20260 8792
rect 20312 8780 20318 8832
rect 22465 8823 22523 8829
rect 22465 8789 22477 8823
rect 22511 8820 22523 8823
rect 23216 8820 23244 8851
rect 27338 8848 27344 8860
rect 27396 8848 27402 8900
rect 22511 8792 23244 8820
rect 36081 8823 36139 8829
rect 22511 8789 22523 8792
rect 22465 8783 22523 8789
rect 36081 8789 36093 8823
rect 36127 8820 36139 8823
rect 36446 8820 36452 8832
rect 36127 8792 36452 8820
rect 36127 8789 36139 8792
rect 36081 8783 36139 8789
rect 36446 8780 36452 8792
rect 36504 8780 36510 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1762 8616 1768 8628
rect 1723 8588 1768 8616
rect 1762 8576 1768 8588
rect 1820 8576 1826 8628
rect 15378 8616 15384 8628
rect 15339 8588 15384 8616
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15470 8576 15476 8628
rect 15528 8616 15534 8628
rect 19150 8616 19156 8628
rect 15528 8588 19156 8616
rect 15528 8576 15534 8588
rect 19150 8576 19156 8588
rect 19208 8576 19214 8628
rect 27249 8619 27307 8625
rect 27249 8585 27261 8619
rect 27295 8616 27307 8619
rect 27522 8616 27528 8628
rect 27295 8588 27528 8616
rect 27295 8585 27307 8588
rect 27249 8579 27307 8585
rect 27522 8576 27528 8588
rect 27580 8576 27586 8628
rect 36906 8576 36912 8628
rect 36964 8616 36970 8628
rect 38105 8619 38163 8625
rect 38105 8616 38117 8619
rect 36964 8588 38117 8616
rect 36964 8576 36970 8588
rect 38105 8585 38117 8588
rect 38151 8585 38163 8619
rect 38105 8579 38163 8585
rect 1670 8508 1676 8560
rect 1728 8548 1734 8560
rect 2409 8551 2467 8557
rect 2409 8548 2421 8551
rect 1728 8520 2421 8548
rect 1728 8508 1734 8520
rect 2409 8517 2421 8520
rect 2455 8517 2467 8551
rect 2409 8511 2467 8517
rect 12084 8520 16574 8548
rect 1486 8440 1492 8492
rect 1544 8480 1550 8492
rect 12084 8489 12112 8520
rect 1581 8483 1639 8489
rect 1581 8480 1593 8483
rect 1544 8452 1593 8480
rect 1544 8440 1550 8452
rect 1581 8449 1593 8452
rect 1627 8449 1639 8483
rect 1581 8443 1639 8449
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8449 2375 8483
rect 2317 8443 2375 8449
rect 12069 8483 12127 8489
rect 12069 8449 12081 8483
rect 12115 8449 12127 8483
rect 12069 8443 12127 8449
rect 1210 8372 1216 8424
rect 1268 8412 1274 8424
rect 2332 8412 2360 8443
rect 12158 8440 12164 8492
rect 12216 8480 12222 8492
rect 13173 8483 13231 8489
rect 13173 8480 13185 8483
rect 12216 8452 13185 8480
rect 12216 8440 12222 8452
rect 13173 8449 13185 8452
rect 13219 8449 13231 8483
rect 14642 8480 14648 8492
rect 14603 8452 14648 8480
rect 13173 8443 13231 8449
rect 14642 8440 14648 8452
rect 14700 8440 14706 8492
rect 15565 8483 15623 8489
rect 15565 8449 15577 8483
rect 15611 8480 15623 8483
rect 16206 8480 16212 8492
rect 15611 8452 16068 8480
rect 16167 8452 16212 8480
rect 15611 8449 15623 8452
rect 15565 8443 15623 8449
rect 1268 8384 2360 8412
rect 1268 8372 1274 8384
rect 2958 8372 2964 8424
rect 3016 8412 3022 8424
rect 3053 8415 3111 8421
rect 3053 8412 3065 8415
rect 3016 8384 3065 8412
rect 3016 8372 3022 8384
rect 3053 8381 3065 8384
rect 3099 8381 3111 8415
rect 3053 8375 3111 8381
rect 11146 8372 11152 8424
rect 11204 8412 11210 8424
rect 12176 8412 12204 8440
rect 11204 8384 12204 8412
rect 12253 8415 12311 8421
rect 11204 8372 11210 8384
rect 12253 8381 12265 8415
rect 12299 8412 12311 8415
rect 13265 8415 13323 8421
rect 13265 8412 13277 8415
rect 12299 8384 13277 8412
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 13265 8381 13277 8384
rect 13311 8381 13323 8415
rect 13265 8375 13323 8381
rect 14737 8347 14795 8353
rect 14737 8313 14749 8347
rect 14783 8344 14795 8347
rect 15654 8344 15660 8356
rect 14783 8316 15660 8344
rect 14783 8313 14795 8316
rect 14737 8307 14795 8313
rect 15654 8304 15660 8316
rect 15712 8304 15718 8356
rect 16040 8353 16068 8452
rect 16206 8440 16212 8452
rect 16264 8440 16270 8492
rect 16546 8412 16574 8520
rect 17218 8508 17224 8560
rect 17276 8548 17282 8560
rect 25222 8548 25228 8560
rect 17276 8520 25228 8548
rect 17276 8508 17282 8520
rect 25222 8508 25228 8520
rect 25280 8508 25286 8560
rect 20070 8440 20076 8492
rect 20128 8480 20134 8492
rect 20533 8483 20591 8489
rect 20533 8480 20545 8483
rect 20128 8452 20545 8480
rect 20128 8440 20134 8452
rect 20533 8449 20545 8452
rect 20579 8449 20591 8483
rect 20533 8443 20591 8449
rect 26234 8440 26240 8492
rect 26292 8480 26298 8492
rect 27157 8483 27215 8489
rect 27157 8480 27169 8483
rect 26292 8452 27169 8480
rect 26292 8440 26298 8452
rect 27157 8449 27169 8452
rect 27203 8449 27215 8483
rect 36446 8480 36452 8492
rect 36407 8452 36452 8480
rect 27157 8443 27215 8449
rect 36446 8440 36452 8452
rect 36504 8440 36510 8492
rect 38286 8480 38292 8492
rect 38247 8452 38292 8480
rect 38286 8440 38292 8452
rect 38344 8440 38350 8492
rect 23474 8412 23480 8424
rect 16546 8384 23480 8412
rect 23474 8372 23480 8384
rect 23532 8372 23538 8424
rect 16025 8347 16083 8353
rect 16025 8313 16037 8347
rect 16071 8313 16083 8347
rect 16025 8307 16083 8313
rect 20349 8347 20407 8353
rect 20349 8313 20361 8347
rect 20395 8344 20407 8347
rect 23382 8344 23388 8356
rect 20395 8316 23388 8344
rect 20395 8313 20407 8316
rect 20349 8307 20407 8313
rect 23382 8304 23388 8316
rect 23440 8304 23446 8356
rect 36265 8347 36323 8353
rect 36265 8313 36277 8347
rect 36311 8344 36323 8347
rect 38010 8344 38016 8356
rect 36311 8316 38016 8344
rect 36311 8313 36323 8316
rect 36265 8307 36323 8313
rect 38010 8304 38016 8316
rect 38068 8304 38074 8356
rect 12434 8276 12440 8288
rect 12395 8248 12440 8276
rect 12434 8236 12440 8248
rect 12492 8236 12498 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 19521 8075 19579 8081
rect 19521 8041 19533 8075
rect 19567 8072 19579 8075
rect 20530 8072 20536 8084
rect 19567 8044 20536 8072
rect 19567 8041 19579 8044
rect 19521 8035 19579 8041
rect 20530 8032 20536 8044
rect 20588 8032 20594 8084
rect 11238 7964 11244 8016
rect 11296 8004 11302 8016
rect 12158 8004 12164 8016
rect 11296 7976 12164 8004
rect 11296 7964 11302 7976
rect 12158 7964 12164 7976
rect 12216 8004 12222 8016
rect 15289 8007 15347 8013
rect 15289 8004 15301 8007
rect 12216 7976 15301 8004
rect 12216 7964 12222 7976
rect 15289 7973 15301 7976
rect 15335 7973 15347 8007
rect 15289 7967 15347 7973
rect 2133 7939 2191 7945
rect 2133 7905 2145 7939
rect 2179 7936 2191 7939
rect 3050 7936 3056 7948
rect 2179 7908 3056 7936
rect 2179 7905 2191 7908
rect 2133 7899 2191 7905
rect 3050 7896 3056 7908
rect 3108 7896 3114 7948
rect 3145 7939 3203 7945
rect 3145 7905 3157 7939
rect 3191 7936 3203 7939
rect 3602 7936 3608 7948
rect 3191 7908 3608 7936
rect 3191 7905 3203 7908
rect 3145 7899 3203 7905
rect 3602 7896 3608 7908
rect 3660 7896 3666 7948
rect 12434 7936 12440 7948
rect 10244 7908 12440 7936
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7868 4031 7871
rect 5534 7868 5540 7880
rect 4019 7840 5540 7868
rect 4019 7837 4031 7840
rect 3973 7831 4031 7837
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 10244 7877 10272 7908
rect 12434 7896 12440 7908
rect 12492 7936 12498 7948
rect 12529 7939 12587 7945
rect 12529 7936 12541 7939
rect 12492 7908 12541 7936
rect 12492 7896 12498 7908
rect 12529 7905 12541 7908
rect 12575 7905 12587 7939
rect 14734 7936 14740 7948
rect 14695 7908 14740 7936
rect 12529 7899 12587 7905
rect 14734 7896 14740 7908
rect 14792 7896 14798 7948
rect 15304 7936 15332 7967
rect 25869 7939 25927 7945
rect 15304 7908 15424 7936
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 11885 7871 11943 7877
rect 11885 7837 11897 7871
rect 11931 7837 11943 7871
rect 12066 7868 12072 7880
rect 12027 7840 12072 7868
rect 11885 7831 11943 7837
rect 2225 7803 2283 7809
rect 2225 7769 2237 7803
rect 2271 7769 2283 7803
rect 11900 7800 11928 7831
rect 12066 7828 12072 7840
rect 12124 7828 12130 7880
rect 13538 7800 13544 7812
rect 11900 7772 13544 7800
rect 2225 7763 2283 7769
rect 2240 7732 2268 7763
rect 13538 7760 13544 7772
rect 13596 7760 13602 7812
rect 14826 7760 14832 7812
rect 14884 7800 14890 7812
rect 15396 7800 15424 7908
rect 25869 7905 25881 7939
rect 25915 7936 25927 7939
rect 27433 7939 27491 7945
rect 27433 7936 27445 7939
rect 25915 7908 27445 7936
rect 25915 7905 25927 7908
rect 25869 7899 25927 7905
rect 27433 7905 27445 7908
rect 27479 7905 27491 7939
rect 27433 7899 27491 7905
rect 15654 7828 15660 7880
rect 15712 7868 15718 7880
rect 16577 7871 16635 7877
rect 16577 7868 16589 7871
rect 15712 7840 16589 7868
rect 15712 7828 15718 7840
rect 16577 7837 16589 7840
rect 16623 7837 16635 7871
rect 16577 7831 16635 7837
rect 17494 7828 17500 7880
rect 17552 7868 17558 7880
rect 19429 7871 19487 7877
rect 19429 7868 19441 7871
rect 17552 7840 19441 7868
rect 17552 7828 17558 7840
rect 19429 7837 19441 7840
rect 19475 7837 19487 7871
rect 19429 7831 19487 7837
rect 23477 7871 23535 7877
rect 23477 7837 23489 7871
rect 23523 7868 23535 7871
rect 25590 7868 25596 7880
rect 23523 7840 25596 7868
rect 23523 7837 23535 7840
rect 23477 7831 23535 7837
rect 25590 7828 25596 7840
rect 25648 7828 25654 7880
rect 27338 7868 27344 7880
rect 27299 7840 27344 7868
rect 27338 7828 27344 7840
rect 27396 7828 27402 7880
rect 38286 7868 38292 7880
rect 38247 7840 38292 7868
rect 38286 7828 38292 7840
rect 38344 7828 38350 7880
rect 20070 7800 20076 7812
rect 14884 7772 14929 7800
rect 15396 7772 20076 7800
rect 14884 7760 14890 7772
rect 20070 7760 20076 7772
rect 20128 7760 20134 7812
rect 21542 7800 21548 7812
rect 21503 7772 21548 7800
rect 21542 7760 21548 7772
rect 21600 7760 21606 7812
rect 21634 7760 21640 7812
rect 21692 7800 21698 7812
rect 21692 7772 21737 7800
rect 21692 7760 21698 7772
rect 22094 7760 22100 7812
rect 22152 7800 22158 7812
rect 22557 7803 22615 7809
rect 22557 7800 22569 7803
rect 22152 7772 22569 7800
rect 22152 7760 22158 7772
rect 22557 7769 22569 7772
rect 22603 7800 22615 7803
rect 25961 7803 26019 7809
rect 22603 7772 23704 7800
rect 22603 7769 22615 7772
rect 22557 7763 22615 7769
rect 4065 7735 4123 7741
rect 4065 7732 4077 7735
rect 2240 7704 4077 7732
rect 4065 7701 4077 7704
rect 4111 7701 4123 7735
rect 10318 7732 10324 7744
rect 10279 7704 10324 7732
rect 4065 7695 4123 7701
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 12894 7692 12900 7744
rect 12952 7732 12958 7744
rect 12989 7735 13047 7741
rect 12989 7732 13001 7735
rect 12952 7704 13001 7732
rect 12952 7692 12958 7704
rect 12989 7701 13001 7704
rect 13035 7701 13047 7735
rect 12989 7695 13047 7701
rect 16393 7735 16451 7741
rect 16393 7701 16405 7735
rect 16439 7732 16451 7735
rect 17862 7732 17868 7744
rect 16439 7704 17868 7732
rect 16439 7701 16451 7704
rect 16393 7695 16451 7701
rect 17862 7692 17868 7704
rect 17920 7692 17926 7744
rect 19426 7692 19432 7744
rect 19484 7732 19490 7744
rect 19978 7732 19984 7744
rect 19484 7704 19984 7732
rect 19484 7692 19490 7704
rect 19978 7692 19984 7704
rect 20036 7732 20042 7744
rect 23569 7735 23627 7741
rect 23569 7732 23581 7735
rect 20036 7704 23581 7732
rect 20036 7692 20042 7704
rect 23569 7701 23581 7704
rect 23615 7701 23627 7735
rect 23676 7732 23704 7772
rect 25961 7769 25973 7803
rect 26007 7800 26019 7803
rect 26050 7800 26056 7812
rect 26007 7772 26056 7800
rect 26007 7769 26019 7772
rect 25961 7763 26019 7769
rect 26050 7760 26056 7772
rect 26108 7760 26114 7812
rect 26881 7803 26939 7809
rect 26881 7800 26893 7803
rect 26206 7772 26893 7800
rect 26206 7732 26234 7772
rect 26881 7769 26893 7772
rect 26927 7769 26939 7803
rect 26881 7763 26939 7769
rect 23676 7704 26234 7732
rect 23569 7695 23627 7701
rect 36354 7692 36360 7744
rect 36412 7732 36418 7744
rect 38105 7735 38163 7741
rect 38105 7732 38117 7735
rect 36412 7704 38117 7732
rect 36412 7692 36418 7704
rect 38105 7701 38117 7704
rect 38151 7701 38163 7735
rect 38105 7695 38163 7701
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 1578 7528 1584 7540
rect 1539 7500 1584 7528
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 13538 7528 13544 7540
rect 13499 7500 13544 7528
rect 13538 7488 13544 7500
rect 13596 7488 13602 7540
rect 14737 7531 14795 7537
rect 14737 7497 14749 7531
rect 14783 7528 14795 7531
rect 14826 7528 14832 7540
rect 14783 7500 14832 7528
rect 14783 7497 14795 7500
rect 14737 7491 14795 7497
rect 14826 7488 14832 7500
rect 14884 7488 14890 7540
rect 21542 7488 21548 7540
rect 21600 7528 21606 7540
rect 22097 7531 22155 7537
rect 22097 7528 22109 7531
rect 21600 7500 22109 7528
rect 21600 7488 21606 7500
rect 22097 7497 22109 7500
rect 22143 7497 22155 7531
rect 22097 7491 22155 7497
rect 2958 7460 2964 7472
rect 2919 7432 2964 7460
rect 2958 7420 2964 7432
rect 3016 7420 3022 7472
rect 3053 7463 3111 7469
rect 3053 7429 3065 7463
rect 3099 7460 3111 7463
rect 3234 7460 3240 7472
rect 3099 7432 3240 7460
rect 3099 7429 3111 7432
rect 3053 7423 3111 7429
rect 3234 7420 3240 7432
rect 3292 7420 3298 7472
rect 3973 7463 4031 7469
rect 3973 7429 3985 7463
rect 4019 7460 4031 7463
rect 5718 7460 5724 7472
rect 4019 7432 5724 7460
rect 4019 7429 4031 7432
rect 3973 7423 4031 7429
rect 5718 7420 5724 7432
rect 5776 7420 5782 7472
rect 11882 7460 11888 7472
rect 11843 7432 11888 7460
rect 11882 7420 11888 7432
rect 11940 7420 11946 7472
rect 18322 7460 18328 7472
rect 18283 7432 18328 7460
rect 18322 7420 18328 7432
rect 18380 7420 18386 7472
rect 19150 7420 19156 7472
rect 19208 7460 19214 7472
rect 19245 7463 19303 7469
rect 19245 7460 19257 7463
rect 19208 7432 19257 7460
rect 19208 7420 19214 7432
rect 19245 7429 19257 7432
rect 19291 7429 19303 7463
rect 19245 7423 19303 7429
rect 19426 7420 19432 7472
rect 19484 7460 19490 7472
rect 19889 7463 19947 7469
rect 19889 7460 19901 7463
rect 19484 7432 19901 7460
rect 19484 7420 19490 7432
rect 19889 7429 19901 7432
rect 19935 7429 19947 7463
rect 19889 7423 19947 7429
rect 23109 7463 23167 7469
rect 23109 7429 23121 7463
rect 23155 7460 23167 7463
rect 23474 7460 23480 7472
rect 23155 7432 23480 7460
rect 23155 7429 23167 7432
rect 23109 7423 23167 7429
rect 23474 7420 23480 7432
rect 23532 7420 23538 7472
rect 1762 7392 1768 7404
rect 1723 7364 1768 7392
rect 1762 7352 1768 7364
rect 1820 7352 1826 7404
rect 1946 7352 1952 7404
rect 2004 7392 2010 7404
rect 2225 7395 2283 7401
rect 2225 7392 2237 7395
rect 2004 7364 2237 7392
rect 2004 7352 2010 7364
rect 2225 7361 2237 7364
rect 2271 7361 2283 7395
rect 2225 7355 2283 7361
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7392 6607 7395
rect 10962 7392 10968 7404
rect 6595 7364 10968 7392
rect 6595 7361 6607 7364
rect 6549 7355 6607 7361
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 11146 7392 11152 7404
rect 11107 7364 11152 7392
rect 11146 7352 11152 7364
rect 11204 7352 11210 7404
rect 12894 7392 12900 7404
rect 12855 7364 12900 7392
rect 12894 7352 12900 7364
rect 12952 7352 12958 7404
rect 14274 7352 14280 7404
rect 14332 7392 14338 7404
rect 14645 7395 14703 7401
rect 14645 7392 14657 7395
rect 14332 7364 14657 7392
rect 14332 7352 14338 7364
rect 14645 7361 14657 7364
rect 14691 7392 14703 7395
rect 15562 7392 15568 7404
rect 14691 7364 15568 7392
rect 14691 7361 14703 7364
rect 14645 7355 14703 7361
rect 15562 7352 15568 7364
rect 15620 7352 15626 7404
rect 22002 7392 22008 7404
rect 21963 7364 22008 7392
rect 22002 7352 22008 7364
rect 22060 7352 22066 7404
rect 11790 7324 11796 7336
rect 11751 7296 11796 7324
rect 11790 7284 11796 7296
rect 11848 7284 11854 7336
rect 12158 7324 12164 7336
rect 12119 7296 12164 7324
rect 12158 7284 12164 7296
rect 12216 7284 12222 7336
rect 13078 7324 13084 7336
rect 13039 7296 13084 7324
rect 13078 7284 13084 7296
rect 13136 7284 13142 7336
rect 17402 7324 17408 7336
rect 17363 7296 17408 7324
rect 17402 7284 17408 7296
rect 17460 7284 17466 7336
rect 18230 7324 18236 7336
rect 18191 7296 18236 7324
rect 18230 7284 18236 7296
rect 18288 7284 18294 7336
rect 19797 7327 19855 7333
rect 19797 7293 19809 7327
rect 19843 7324 19855 7327
rect 19886 7324 19892 7336
rect 19843 7296 19892 7324
rect 19843 7293 19855 7296
rect 19797 7287 19855 7293
rect 19886 7284 19892 7296
rect 19944 7284 19950 7336
rect 20070 7324 20076 7336
rect 20031 7296 20076 7324
rect 20070 7284 20076 7296
rect 20128 7284 20134 7336
rect 23017 7327 23075 7333
rect 23017 7293 23029 7327
rect 23063 7324 23075 7327
rect 24578 7324 24584 7336
rect 23063 7296 24584 7324
rect 23063 7293 23075 7296
rect 23017 7287 23075 7293
rect 24578 7284 24584 7296
rect 24636 7284 24642 7336
rect 23566 7256 23572 7268
rect 23527 7228 23572 7256
rect 23566 7216 23572 7228
rect 23624 7216 23630 7268
rect 2317 7191 2375 7197
rect 2317 7157 2329 7191
rect 2363 7188 2375 7191
rect 3234 7188 3240 7200
rect 2363 7160 3240 7188
rect 2363 7157 2375 7160
rect 2317 7151 2375 7157
rect 3234 7148 3240 7160
rect 3292 7148 3298 7200
rect 6641 7191 6699 7197
rect 6641 7157 6653 7191
rect 6687 7188 6699 7191
rect 6730 7188 6736 7200
rect 6687 7160 6736 7188
rect 6687 7157 6699 7160
rect 6641 7151 6699 7157
rect 6730 7148 6736 7160
rect 6788 7148 6794 7200
rect 10965 7191 11023 7197
rect 10965 7157 10977 7191
rect 11011 7188 11023 7191
rect 11698 7188 11704 7200
rect 11011 7160 11704 7188
rect 11011 7157 11023 7160
rect 10965 7151 11023 7157
rect 11698 7148 11704 7160
rect 11756 7148 11762 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 11517 6987 11575 6993
rect 11517 6953 11529 6987
rect 11563 6984 11575 6987
rect 12066 6984 12072 6996
rect 11563 6956 12072 6984
rect 11563 6953 11575 6956
rect 11517 6947 11575 6953
rect 12066 6944 12072 6956
rect 12124 6944 12130 6996
rect 23474 6984 23480 6996
rect 23435 6956 23480 6984
rect 23474 6944 23480 6956
rect 23532 6944 23538 6996
rect 12437 6851 12495 6857
rect 12437 6817 12449 6851
rect 12483 6848 12495 6851
rect 14734 6848 14740 6860
rect 12483 6820 14740 6848
rect 12483 6817 12495 6820
rect 12437 6811 12495 6817
rect 14734 6808 14740 6820
rect 14792 6808 14798 6860
rect 17313 6851 17371 6857
rect 17313 6817 17325 6851
rect 17359 6848 17371 6851
rect 17402 6848 17408 6860
rect 17359 6820 17408 6848
rect 17359 6817 17371 6820
rect 17313 6811 17371 6817
rect 17402 6808 17408 6820
rect 17460 6808 17466 6860
rect 17957 6851 18015 6857
rect 17957 6817 17969 6851
rect 18003 6848 18015 6851
rect 18230 6848 18236 6860
rect 18003 6820 18236 6848
rect 18003 6817 18015 6820
rect 17957 6811 18015 6817
rect 1762 6780 1768 6792
rect 1723 6752 1768 6780
rect 1762 6740 1768 6752
rect 1820 6740 1826 6792
rect 3234 6780 3240 6792
rect 3195 6752 3240 6780
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 6825 6783 6883 6789
rect 6825 6749 6837 6783
rect 6871 6780 6883 6783
rect 10318 6780 10324 6792
rect 6871 6752 10324 6780
rect 6871 6749 6883 6752
rect 6825 6743 6883 6749
rect 10318 6740 10324 6752
rect 10376 6740 10382 6792
rect 11698 6780 11704 6792
rect 11659 6752 11704 6780
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 12342 6780 12348 6792
rect 12303 6752 12348 6780
rect 12342 6740 12348 6752
rect 12400 6740 12406 6792
rect 14366 6740 14372 6792
rect 14424 6780 14430 6792
rect 15381 6783 15439 6789
rect 15381 6780 15393 6783
rect 14424 6752 15393 6780
rect 14424 6740 14430 6752
rect 15381 6749 15393 6752
rect 15427 6749 15439 6783
rect 15381 6743 15439 6749
rect 15565 6783 15623 6789
rect 15565 6749 15577 6783
rect 15611 6780 15623 6783
rect 15654 6780 15660 6792
rect 15611 6752 15660 6780
rect 15611 6749 15623 6752
rect 15565 6743 15623 6749
rect 15654 6740 15660 6752
rect 15712 6740 15718 6792
rect 17497 6783 17555 6789
rect 17497 6749 17509 6783
rect 17543 6780 17555 6783
rect 17586 6780 17592 6792
rect 17543 6752 17592 6780
rect 17543 6749 17555 6752
rect 17497 6743 17555 6749
rect 17586 6740 17592 6752
rect 17644 6740 17650 6792
rect 16025 6715 16083 6721
rect 16025 6681 16037 6715
rect 16071 6712 16083 6715
rect 17972 6712 18000 6811
rect 18230 6808 18236 6820
rect 18288 6808 18294 6860
rect 19797 6783 19855 6789
rect 19797 6749 19809 6783
rect 19843 6780 19855 6783
rect 20714 6780 20720 6792
rect 19843 6752 20720 6780
rect 19843 6749 19855 6752
rect 19797 6743 19855 6749
rect 20714 6740 20720 6752
rect 20772 6740 20778 6792
rect 22370 6740 22376 6792
rect 22428 6780 22434 6792
rect 23017 6783 23075 6789
rect 23017 6780 23029 6783
rect 22428 6752 23029 6780
rect 22428 6740 22434 6752
rect 23017 6749 23029 6752
rect 23063 6749 23075 6783
rect 23017 6743 23075 6749
rect 23661 6783 23719 6789
rect 23661 6749 23673 6783
rect 23707 6749 23719 6783
rect 23661 6743 23719 6749
rect 16071 6684 18000 6712
rect 16071 6681 16083 6684
rect 16025 6675 16083 6681
rect 1394 6604 1400 6656
rect 1452 6644 1458 6656
rect 1581 6647 1639 6653
rect 1581 6644 1593 6647
rect 1452 6616 1593 6644
rect 1452 6604 1458 6616
rect 1581 6613 1593 6616
rect 1627 6613 1639 6647
rect 3050 6644 3056 6656
rect 3011 6616 3056 6644
rect 1581 6607 1639 6613
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 6638 6644 6644 6656
rect 6599 6616 6644 6644
rect 6638 6604 6644 6616
rect 6696 6604 6702 6656
rect 15010 6604 15016 6656
rect 15068 6644 15074 6656
rect 19334 6644 19340 6656
rect 15068 6616 19340 6644
rect 15068 6604 15074 6616
rect 19334 6604 19340 6616
rect 19392 6644 19398 6656
rect 19889 6647 19947 6653
rect 19889 6644 19901 6647
rect 19392 6616 19901 6644
rect 19392 6604 19398 6616
rect 19889 6613 19901 6616
rect 19935 6613 19947 6647
rect 19889 6607 19947 6613
rect 22833 6647 22891 6653
rect 22833 6613 22845 6647
rect 22879 6644 22891 6647
rect 23676 6644 23704 6743
rect 22879 6616 23704 6644
rect 22879 6613 22891 6616
rect 22833 6607 22891 6613
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 1946 6440 1952 6452
rect 1907 6412 1952 6440
rect 1946 6400 1952 6412
rect 2004 6400 2010 6452
rect 11790 6400 11796 6452
rect 11848 6440 11854 6452
rect 11885 6443 11943 6449
rect 11885 6440 11897 6443
rect 11848 6412 11897 6440
rect 11848 6400 11854 6412
rect 11885 6409 11897 6412
rect 11931 6409 11943 6443
rect 11885 6403 11943 6409
rect 13078 6400 13084 6452
rect 13136 6440 13142 6452
rect 13173 6443 13231 6449
rect 13173 6440 13185 6443
rect 13136 6412 13185 6440
rect 13136 6400 13142 6412
rect 13173 6409 13185 6412
rect 13219 6409 13231 6443
rect 13173 6403 13231 6409
rect 13817 6443 13875 6449
rect 13817 6409 13829 6443
rect 13863 6409 13875 6443
rect 15654 6440 15660 6452
rect 15615 6412 15660 6440
rect 13817 6403 13875 6409
rect 1857 6375 1915 6381
rect 1857 6341 1869 6375
rect 1903 6372 1915 6375
rect 2866 6372 2872 6384
rect 1903 6344 2872 6372
rect 1903 6341 1915 6344
rect 1857 6335 1915 6341
rect 2866 6332 2872 6344
rect 2924 6332 2930 6384
rect 6730 6304 6736 6316
rect 6691 6276 6736 6304
rect 6730 6264 6736 6276
rect 6788 6264 6794 6316
rect 11793 6307 11851 6313
rect 11793 6273 11805 6307
rect 11839 6304 11851 6307
rect 12986 6304 12992 6316
rect 11839 6276 12992 6304
rect 11839 6273 11851 6276
rect 11793 6267 11851 6273
rect 12986 6264 12992 6276
rect 13044 6264 13050 6316
rect 13357 6307 13415 6313
rect 13357 6273 13369 6307
rect 13403 6304 13415 6307
rect 13832 6304 13860 6403
rect 15654 6400 15660 6412
rect 15712 6400 15718 6452
rect 17586 6440 17592 6452
rect 17547 6412 17592 6440
rect 17586 6400 17592 6412
rect 17644 6400 17650 6452
rect 18509 6443 18567 6449
rect 18509 6409 18521 6443
rect 18555 6440 18567 6443
rect 19426 6440 19432 6452
rect 18555 6412 19432 6440
rect 18555 6409 18567 6412
rect 18509 6403 18567 6409
rect 19426 6400 19432 6412
rect 19484 6400 19490 6452
rect 24578 6400 24584 6452
rect 24636 6440 24642 6452
rect 25961 6443 26019 6449
rect 25961 6440 25973 6443
rect 24636 6412 25973 6440
rect 24636 6400 24642 6412
rect 25961 6409 25973 6412
rect 26007 6409 26019 6443
rect 25961 6403 26019 6409
rect 13998 6304 14004 6316
rect 13403 6276 13860 6304
rect 13959 6276 14004 6304
rect 13403 6273 13415 6276
rect 13357 6267 13415 6273
rect 13998 6264 14004 6276
rect 14056 6264 14062 6316
rect 15562 6304 15568 6316
rect 15523 6276 15568 6304
rect 15562 6264 15568 6276
rect 15620 6264 15626 6316
rect 16574 6264 16580 6316
rect 16632 6304 16638 6316
rect 17497 6307 17555 6313
rect 17497 6304 17509 6307
rect 16632 6276 17509 6304
rect 16632 6264 16638 6276
rect 17497 6273 17509 6276
rect 17543 6304 17555 6307
rect 18417 6307 18475 6313
rect 18417 6304 18429 6307
rect 17543 6276 18429 6304
rect 17543 6273 17555 6276
rect 17497 6267 17555 6273
rect 18417 6273 18429 6276
rect 18463 6273 18475 6307
rect 18417 6267 18475 6273
rect 25225 6307 25283 6313
rect 25225 6273 25237 6307
rect 25271 6304 25283 6307
rect 25314 6304 25320 6316
rect 25271 6276 25320 6304
rect 25271 6273 25283 6276
rect 25225 6267 25283 6273
rect 25314 6264 25320 6276
rect 25372 6264 25378 6316
rect 25869 6307 25927 6313
rect 25869 6273 25881 6307
rect 25915 6304 25927 6307
rect 27522 6304 27528 6316
rect 25915 6276 27528 6304
rect 25915 6273 25927 6276
rect 25869 6267 25927 6273
rect 27522 6264 27528 6276
rect 27580 6264 27586 6316
rect 38286 6304 38292 6316
rect 38247 6276 38292 6304
rect 38286 6264 38292 6276
rect 38344 6264 38350 6316
rect 4062 6060 4068 6112
rect 4120 6100 4126 6112
rect 6549 6103 6607 6109
rect 6549 6100 6561 6103
rect 4120 6072 6561 6100
rect 4120 6060 4126 6072
rect 6549 6069 6561 6072
rect 6595 6069 6607 6103
rect 6549 6063 6607 6069
rect 25317 6103 25375 6109
rect 25317 6069 25329 6103
rect 25363 6100 25375 6103
rect 25682 6100 25688 6112
rect 25363 6072 25688 6100
rect 25363 6069 25375 6072
rect 25317 6063 25375 6069
rect 25682 6060 25688 6072
rect 25740 6060 25746 6112
rect 27430 6060 27436 6112
rect 27488 6100 27494 6112
rect 38105 6103 38163 6109
rect 38105 6100 38117 6103
rect 27488 6072 38117 6100
rect 27488 6060 27494 6072
rect 38105 6069 38117 6072
rect 38151 6069 38163 6103
rect 38105 6063 38163 6069
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 14366 5896 14372 5908
rect 14327 5868 14372 5896
rect 14366 5856 14372 5868
rect 14424 5856 14430 5908
rect 27706 5896 27712 5908
rect 27667 5868 27712 5896
rect 27706 5856 27712 5868
rect 27764 5856 27770 5908
rect 2038 5828 2044 5840
rect 1999 5800 2044 5828
rect 2038 5788 2044 5800
rect 2096 5788 2102 5840
rect 2498 5692 2504 5704
rect 2459 5664 2504 5692
rect 2498 5652 2504 5664
rect 2556 5652 2562 5704
rect 12526 5652 12532 5704
rect 12584 5692 12590 5704
rect 14277 5695 14335 5701
rect 14277 5692 14289 5695
rect 12584 5664 14289 5692
rect 12584 5652 12590 5664
rect 14277 5661 14289 5664
rect 14323 5661 14335 5695
rect 25682 5692 25688 5704
rect 25643 5664 25688 5692
rect 14277 5655 14335 5661
rect 25682 5652 25688 5664
rect 25740 5652 25746 5704
rect 27617 5695 27675 5701
rect 27617 5661 27629 5695
rect 27663 5692 27675 5695
rect 30282 5692 30288 5704
rect 27663 5664 30288 5692
rect 27663 5661 27675 5664
rect 27617 5655 27675 5661
rect 30282 5652 30288 5664
rect 30340 5652 30346 5704
rect 1857 5627 1915 5633
rect 1857 5593 1869 5627
rect 1903 5624 1915 5627
rect 2593 5627 2651 5633
rect 2593 5624 2605 5627
rect 1903 5596 2605 5624
rect 1903 5593 1915 5596
rect 1857 5587 1915 5593
rect 2593 5593 2605 5596
rect 2639 5593 2651 5627
rect 2593 5587 2651 5593
rect 25222 5516 25228 5568
rect 25280 5556 25286 5568
rect 25501 5559 25559 5565
rect 25501 5556 25513 5559
rect 25280 5528 25513 5556
rect 25280 5516 25286 5528
rect 25501 5525 25513 5528
rect 25547 5525 25559 5559
rect 25501 5519 25559 5525
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 6546 5352 6552 5364
rect 1627 5324 6552 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 6546 5312 6552 5324
rect 6604 5312 6610 5364
rect 15746 5312 15752 5364
rect 15804 5352 15810 5364
rect 15804 5324 18736 5352
rect 15804 5312 15810 5324
rect 16022 5244 16028 5296
rect 16080 5284 16086 5296
rect 17773 5287 17831 5293
rect 17773 5284 17785 5287
rect 16080 5256 17785 5284
rect 16080 5244 16086 5256
rect 17773 5253 17785 5256
rect 17819 5253 17831 5287
rect 17773 5247 17831 5253
rect 1762 5216 1768 5228
rect 1723 5188 1768 5216
rect 1762 5176 1768 5188
rect 1820 5176 1826 5228
rect 17681 5151 17739 5157
rect 17681 5117 17693 5151
rect 17727 5148 17739 5151
rect 18506 5148 18512 5160
rect 17727 5120 18512 5148
rect 17727 5117 17739 5120
rect 17681 5111 17739 5117
rect 18506 5108 18512 5120
rect 18564 5108 18570 5160
rect 18708 5157 18736 5324
rect 29914 5216 29920 5228
rect 29875 5188 29920 5216
rect 29914 5176 29920 5188
rect 29972 5176 29978 5228
rect 38010 5216 38016 5228
rect 37971 5188 38016 5216
rect 38010 5176 38016 5188
rect 38068 5176 38074 5228
rect 18693 5151 18751 5157
rect 18693 5117 18705 5151
rect 18739 5148 18751 5151
rect 20530 5148 20536 5160
rect 18739 5120 20536 5148
rect 18739 5117 18751 5120
rect 18693 5111 18751 5117
rect 20530 5108 20536 5120
rect 20588 5108 20594 5160
rect 30009 5015 30067 5021
rect 30009 4981 30021 5015
rect 30055 5012 30067 5015
rect 31662 5012 31668 5024
rect 30055 4984 31668 5012
rect 30055 4981 30067 4984
rect 30009 4975 30067 4981
rect 31662 4972 31668 4984
rect 31720 4972 31726 5024
rect 38194 5012 38200 5024
rect 38155 4984 38200 5012
rect 38194 4972 38200 4984
rect 38252 4972 38258 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 37182 4768 37188 4820
rect 37240 4808 37246 4820
rect 38105 4811 38163 4817
rect 38105 4808 38117 4811
rect 37240 4780 38117 4808
rect 37240 4768 37246 4780
rect 38105 4777 38117 4780
rect 38151 4777 38163 4811
rect 38105 4771 38163 4777
rect 1581 4607 1639 4613
rect 1581 4573 1593 4607
rect 1627 4604 1639 4607
rect 6638 4604 6644 4616
rect 1627 4576 6644 4604
rect 1627 4573 1639 4576
rect 1581 4567 1639 4573
rect 6638 4564 6644 4576
rect 6696 4564 6702 4616
rect 38286 4604 38292 4616
rect 38247 4576 38292 4604
rect 38286 4564 38292 4576
rect 38344 4564 38350 4616
rect 1762 4468 1768 4480
rect 1723 4440 1768 4468
rect 1762 4428 1768 4440
rect 1820 4428 1826 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 37182 4156 37188 4208
rect 37240 4196 37246 4208
rect 38105 4199 38163 4205
rect 38105 4196 38117 4199
rect 37240 4168 38117 4196
rect 37240 4156 37246 4168
rect 38105 4165 38117 4168
rect 38151 4165 38163 4199
rect 38105 4159 38163 4165
rect 1394 4088 1400 4140
rect 1452 4128 1458 4140
rect 1765 4131 1823 4137
rect 1765 4128 1777 4131
rect 1452 4100 1777 4128
rect 1452 4088 1458 4100
rect 1765 4097 1777 4100
rect 1811 4097 1823 4131
rect 1765 4091 1823 4097
rect 5718 4088 5724 4140
rect 5776 4128 5782 4140
rect 6825 4131 6883 4137
rect 6825 4128 6837 4131
rect 5776 4100 6837 4128
rect 5776 4088 5782 4100
rect 6825 4097 6837 4100
rect 6871 4097 6883 4131
rect 6825 4091 6883 4097
rect 18601 4131 18659 4137
rect 18601 4097 18613 4131
rect 18647 4128 18659 4131
rect 19426 4128 19432 4140
rect 18647 4100 19432 4128
rect 18647 4097 18659 4100
rect 18601 4091 18659 4097
rect 19426 4088 19432 4100
rect 19484 4088 19490 4140
rect 20530 4128 20536 4140
rect 20491 4100 20536 4128
rect 20530 4088 20536 4100
rect 20588 4088 20594 4140
rect 36354 4128 36360 4140
rect 36315 4100 36360 4128
rect 36354 4088 36360 4100
rect 36412 4088 36418 4140
rect 18506 4020 18512 4072
rect 18564 4060 18570 4072
rect 18693 4063 18751 4069
rect 18693 4060 18705 4063
rect 18564 4032 18705 4060
rect 18564 4020 18570 4032
rect 18693 4029 18705 4032
rect 18739 4029 18751 4063
rect 18693 4023 18751 4029
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3992 1639 3995
rect 5626 3992 5632 4004
rect 1627 3964 5632 3992
rect 1627 3961 1639 3964
rect 1581 3955 1639 3961
rect 5626 3952 5632 3964
rect 5684 3952 5690 4004
rect 21726 3952 21732 4004
rect 21784 3992 21790 4004
rect 38289 3995 38347 4001
rect 38289 3992 38301 3995
rect 21784 3964 38301 3992
rect 21784 3952 21790 3964
rect 38289 3961 38301 3964
rect 38335 3961 38347 3995
rect 38289 3955 38347 3961
rect 6730 3884 6736 3936
rect 6788 3924 6794 3936
rect 6917 3927 6975 3933
rect 6917 3924 6929 3927
rect 6788 3896 6929 3924
rect 6788 3884 6794 3896
rect 6917 3893 6929 3896
rect 6963 3893 6975 3927
rect 6917 3887 6975 3893
rect 20625 3927 20683 3933
rect 20625 3893 20637 3927
rect 20671 3924 20683 3927
rect 21910 3924 21916 3936
rect 20671 3896 21916 3924
rect 20671 3893 20683 3896
rect 20625 3887 20683 3893
rect 21910 3884 21916 3896
rect 21968 3884 21974 3936
rect 34790 3884 34796 3936
rect 34848 3924 34854 3936
rect 36173 3927 36231 3933
rect 36173 3924 36185 3927
rect 34848 3896 36185 3924
rect 34848 3884 34854 3896
rect 36173 3893 36185 3896
rect 36219 3893 36231 3927
rect 36173 3887 36231 3893
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3516 1915 3519
rect 2225 3519 2283 3525
rect 2225 3516 2237 3519
rect 1903 3488 2237 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 2225 3485 2237 3488
rect 2271 3516 2283 3519
rect 21910 3516 21916 3528
rect 2271 3488 2774 3516
rect 21871 3488 21916 3516
rect 2271 3485 2283 3488
rect 2225 3479 2283 3485
rect 2746 3448 2774 3488
rect 21910 3476 21916 3488
rect 21968 3476 21974 3528
rect 31662 3476 31668 3528
rect 31720 3516 31726 3528
rect 32769 3519 32827 3525
rect 32769 3516 32781 3519
rect 31720 3488 32781 3516
rect 31720 3476 31726 3488
rect 32769 3485 32781 3488
rect 32815 3485 32827 3519
rect 32769 3479 32827 3485
rect 37918 3476 37924 3528
rect 37976 3516 37982 3528
rect 38013 3519 38071 3525
rect 38013 3516 38025 3519
rect 37976 3488 38025 3516
rect 37976 3476 37982 3488
rect 38013 3485 38025 3488
rect 38059 3485 38071 3519
rect 38013 3479 38071 3485
rect 30558 3448 30564 3460
rect 2746 3420 30564 3448
rect 30558 3408 30564 3420
rect 30616 3408 30622 3460
rect 37369 3451 37427 3457
rect 37369 3417 37381 3451
rect 37415 3448 37427 3451
rect 37415 3420 38056 3448
rect 37415 3417 37427 3420
rect 37369 3411 37427 3417
rect 38028 3392 38056 3420
rect 1670 3380 1676 3392
rect 1631 3352 1676 3380
rect 1670 3340 1676 3352
rect 1728 3340 1734 3392
rect 21729 3383 21787 3389
rect 21729 3349 21741 3383
rect 21775 3380 21787 3383
rect 22646 3380 22652 3392
rect 21775 3352 22652 3380
rect 21775 3349 21787 3352
rect 21729 3343 21787 3349
rect 22646 3340 22652 3352
rect 22704 3340 22710 3392
rect 32585 3383 32643 3389
rect 32585 3349 32597 3383
rect 32631 3380 32643 3383
rect 33778 3380 33784 3392
rect 32631 3352 33784 3380
rect 32631 3349 32643 3352
rect 32585 3343 32643 3349
rect 33778 3340 33784 3352
rect 33836 3340 33842 3392
rect 37458 3380 37464 3392
rect 37419 3352 37464 3380
rect 37458 3340 37464 3352
rect 37516 3340 37522 3392
rect 38010 3340 38016 3392
rect 38068 3340 38074 3392
rect 38194 3380 38200 3392
rect 38155 3352 38200 3380
rect 38194 3340 38200 3352
rect 38252 3340 38258 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 3053 3179 3111 3185
rect 3053 3145 3065 3179
rect 3099 3176 3111 3179
rect 3142 3176 3148 3188
rect 3099 3148 3148 3176
rect 3099 3145 3111 3148
rect 3053 3139 3111 3145
rect 3142 3136 3148 3148
rect 3200 3136 3206 3188
rect 9769 3179 9827 3185
rect 9769 3145 9781 3179
rect 9815 3176 9827 3179
rect 9815 3148 12434 3176
rect 9815 3145 9827 3148
rect 9769 3139 9827 3145
rect 4062 3108 4068 3120
rect 1596 3080 4068 3108
rect 1596 3049 1624 3080
rect 4062 3068 4068 3080
rect 4120 3068 4126 3120
rect 12406 3108 12434 3148
rect 35434 3136 35440 3188
rect 35492 3176 35498 3188
rect 36817 3179 36875 3185
rect 36817 3176 36829 3179
rect 35492 3148 36829 3176
rect 35492 3136 35498 3148
rect 36817 3145 36829 3148
rect 36863 3145 36875 3179
rect 36817 3139 36875 3145
rect 37458 3108 37464 3120
rect 12406 3080 13216 3108
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3040 2375 3043
rect 3050 3040 3056 3052
rect 2363 3012 3056 3040
rect 2363 3009 2375 3012
rect 2317 3003 2375 3009
rect 3050 3000 3056 3012
rect 3108 3000 3114 3052
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3009 3295 3043
rect 6730 3040 6736 3052
rect 6691 3012 6736 3040
rect 3237 3003 3295 3009
rect 2774 2932 2780 2984
rect 2832 2972 2838 2984
rect 3252 2972 3280 3003
rect 6730 3000 6736 3012
rect 6788 3000 6794 3052
rect 9674 3000 9680 3052
rect 9732 3040 9738 3052
rect 13188 3049 13216 3080
rect 26206 3080 37464 3108
rect 9953 3043 10011 3049
rect 9953 3040 9965 3043
rect 9732 3012 9965 3040
rect 9732 3000 9738 3012
rect 9953 3009 9965 3012
rect 9999 3009 10011 3043
rect 9953 3003 10011 3009
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3009 13231 3043
rect 13173 3003 13231 3009
rect 14182 3000 14188 3052
rect 14240 3040 14246 3052
rect 14369 3043 14427 3049
rect 14369 3040 14381 3043
rect 14240 3012 14381 3040
rect 14240 3000 14246 3012
rect 14369 3009 14381 3012
rect 14415 3009 14427 3043
rect 14369 3003 14427 3009
rect 17221 3043 17279 3049
rect 17221 3009 17233 3043
rect 17267 3040 17279 3043
rect 17770 3040 17776 3052
rect 17267 3012 17776 3040
rect 17267 3009 17279 3012
rect 17221 3003 17279 3009
rect 17770 3000 17776 3012
rect 17828 3040 17834 3052
rect 26206 3040 26234 3080
rect 37458 3068 37464 3080
rect 37516 3068 37522 3120
rect 17828 3012 26234 3040
rect 36725 3043 36783 3049
rect 17828 3000 17834 3012
rect 36725 3009 36737 3043
rect 36771 3040 36783 3043
rect 37274 3040 37280 3052
rect 36771 3012 37280 3040
rect 36771 3009 36783 3012
rect 36725 3003 36783 3009
rect 37274 3000 37280 3012
rect 37332 3000 37338 3052
rect 39298 3040 39304 3052
rect 37476 3012 39304 3040
rect 37476 2981 37504 3012
rect 39298 3000 39304 3012
rect 39356 3000 39362 3052
rect 2832 2944 3280 2972
rect 37461 2975 37519 2981
rect 2832 2932 2838 2944
rect 37461 2941 37473 2975
rect 37507 2941 37519 2975
rect 37461 2935 37519 2941
rect 37737 2975 37795 2981
rect 37737 2941 37749 2975
rect 37783 2941 37795 2975
rect 37737 2935 37795 2941
rect 14 2864 20 2916
rect 72 2904 78 2916
rect 2501 2907 2559 2913
rect 2501 2904 2513 2907
rect 72 2876 2513 2904
rect 72 2864 78 2876
rect 2501 2873 2513 2876
rect 2547 2873 2559 2907
rect 2501 2867 2559 2873
rect 14553 2907 14611 2913
rect 14553 2873 14565 2907
rect 14599 2904 14611 2907
rect 24486 2904 24492 2916
rect 14599 2876 24492 2904
rect 14599 2873 14611 2876
rect 14553 2867 14611 2873
rect 24486 2864 24492 2876
rect 24544 2864 24550 2916
rect 27246 2864 27252 2916
rect 27304 2904 27310 2916
rect 37752 2904 37780 2935
rect 27304 2876 37780 2904
rect 27304 2864 27310 2876
rect 658 2796 664 2848
rect 716 2836 722 2848
rect 1765 2839 1823 2845
rect 1765 2836 1777 2839
rect 716 2808 1777 2836
rect 716 2796 722 2808
rect 1765 2805 1777 2808
rect 1811 2805 1823 2839
rect 6546 2836 6552 2848
rect 6507 2808 6552 2836
rect 1765 2799 1823 2805
rect 6546 2796 6552 2808
rect 6604 2796 6610 2848
rect 12989 2839 13047 2845
rect 12989 2805 13001 2839
rect 13035 2836 13047 2839
rect 14918 2836 14924 2848
rect 13035 2808 14924 2836
rect 13035 2805 13047 2808
rect 12989 2799 13047 2805
rect 14918 2796 14924 2808
rect 14976 2796 14982 2848
rect 17034 2836 17040 2848
rect 16995 2808 17040 2836
rect 17034 2796 17040 2808
rect 17092 2796 17098 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 7282 2632 7288 2644
rect 7243 2604 7288 2632
rect 7282 2592 7288 2604
rect 7340 2592 7346 2644
rect 11701 2635 11759 2641
rect 11701 2601 11713 2635
rect 11747 2632 11759 2635
rect 12526 2632 12532 2644
rect 11747 2604 12532 2632
rect 11747 2601 11759 2604
rect 11701 2595 11759 2601
rect 12526 2592 12532 2604
rect 12584 2592 12590 2644
rect 12986 2632 12992 2644
rect 12947 2604 12992 2632
rect 12986 2592 12992 2604
rect 13044 2592 13050 2644
rect 16850 2632 16856 2644
rect 16811 2604 16856 2632
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 17494 2632 17500 2644
rect 17455 2604 17500 2632
rect 17494 2592 17500 2604
rect 17552 2592 17558 2644
rect 19426 2632 19432 2644
rect 19387 2604 19432 2632
rect 19426 2592 19432 2604
rect 19484 2592 19490 2644
rect 20714 2632 20720 2644
rect 20675 2604 20720 2632
rect 20714 2592 20720 2604
rect 20772 2592 20778 2644
rect 22002 2632 22008 2644
rect 21963 2604 22008 2632
rect 22002 2592 22008 2604
rect 22060 2592 22066 2644
rect 24581 2635 24639 2641
rect 24581 2601 24593 2635
rect 24627 2632 24639 2635
rect 26234 2632 26240 2644
rect 24627 2604 26240 2632
rect 24627 2601 24639 2604
rect 24581 2595 24639 2601
rect 26234 2592 26240 2604
rect 26292 2592 26298 2644
rect 27157 2635 27215 2641
rect 27157 2601 27169 2635
rect 27203 2632 27215 2635
rect 27338 2632 27344 2644
rect 27203 2604 27344 2632
rect 27203 2601 27215 2604
rect 27157 2595 27215 2601
rect 27338 2592 27344 2604
rect 27396 2592 27402 2644
rect 28445 2635 28503 2641
rect 28445 2632 28457 2635
rect 27448 2604 28457 2632
rect 10410 2564 10416 2576
rect 4264 2536 10416 2564
rect 4264 2505 4292 2536
rect 10410 2524 10416 2536
rect 10468 2524 10474 2576
rect 10965 2567 11023 2573
rect 10965 2533 10977 2567
rect 11011 2564 11023 2567
rect 12342 2564 12348 2576
rect 11011 2536 12348 2564
rect 11011 2533 11023 2536
rect 10965 2527 11023 2533
rect 12342 2524 12348 2536
rect 12400 2524 12406 2576
rect 13262 2524 13268 2576
rect 13320 2564 13326 2576
rect 13320 2536 23336 2564
rect 13320 2524 13326 2536
rect 4249 2499 4307 2505
rect 2056 2468 4200 2496
rect 2056 2437 2084 2468
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2397 2099 2431
rect 2041 2391 2099 2397
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2428 2927 2431
rect 3421 2431 3479 2437
rect 3421 2428 3433 2431
rect 2915 2400 3433 2428
rect 2915 2397 2927 2400
rect 2869 2391 2927 2397
rect 3421 2397 3433 2400
rect 3467 2428 3479 2431
rect 3467 2400 3832 2428
rect 3467 2397 3479 2400
rect 3421 2391 3479 2397
rect 3804 2360 3832 2400
rect 3878 2388 3884 2440
rect 3936 2428 3942 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3936 2400 3985 2428
rect 3936 2388 3942 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 4172 2428 4200 2468
rect 4249 2465 4261 2499
rect 4295 2465 4307 2499
rect 9306 2496 9312 2508
rect 4249 2459 4307 2465
rect 4356 2468 9312 2496
rect 4356 2428 4384 2468
rect 9306 2456 9312 2468
rect 9364 2456 9370 2508
rect 9401 2499 9459 2505
rect 9401 2465 9413 2499
rect 9447 2496 9459 2499
rect 18598 2496 18604 2508
rect 9447 2468 18604 2496
rect 9447 2465 9459 2468
rect 9401 2459 9459 2465
rect 18598 2456 18604 2468
rect 18656 2456 18662 2508
rect 5258 2428 5264 2440
rect 4172 2400 4384 2428
rect 5219 2400 5264 2428
rect 3973 2391 4031 2397
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 6546 2428 6552 2440
rect 6507 2400 6552 2428
rect 6546 2388 6552 2400
rect 6604 2388 6610 2440
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 7156 2400 7481 2428
rect 7156 2388 7162 2400
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8444 2400 9137 2428
rect 8444 2388 8450 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 10962 2388 10968 2440
rect 11020 2428 11026 2440
rect 11149 2431 11207 2437
rect 11149 2428 11161 2431
rect 11020 2400 11161 2428
rect 11020 2388 11026 2400
rect 11149 2397 11161 2400
rect 11195 2397 11207 2431
rect 11149 2391 11207 2397
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 11885 2431 11943 2437
rect 11885 2428 11897 2431
rect 11664 2400 11897 2428
rect 11664 2388 11670 2400
rect 11885 2397 11897 2400
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 12894 2388 12900 2440
rect 12952 2428 12958 2440
rect 13173 2431 13231 2437
rect 13173 2428 13185 2431
rect 12952 2400 13185 2428
rect 12952 2388 12958 2400
rect 13173 2397 13185 2400
rect 13219 2397 13231 2431
rect 14918 2428 14924 2440
rect 14879 2400 14924 2428
rect 13173 2391 13231 2397
rect 14918 2388 14924 2400
rect 14976 2388 14982 2440
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 17037 2431 17095 2437
rect 17037 2428 17049 2431
rect 16172 2400 17049 2428
rect 16172 2388 16178 2400
rect 17037 2397 17049 2400
rect 17083 2397 17095 2431
rect 17037 2391 17095 2397
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 17681 2431 17739 2437
rect 17681 2428 17693 2431
rect 17460 2400 17693 2428
rect 17460 2388 17466 2400
rect 17681 2397 17693 2400
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 17862 2388 17868 2440
rect 17920 2428 17926 2440
rect 18141 2431 18199 2437
rect 18141 2428 18153 2431
rect 17920 2400 18153 2428
rect 17920 2388 17926 2400
rect 18141 2397 18153 2400
rect 18187 2397 18199 2431
rect 18141 2391 18199 2397
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 19392 2400 19625 2428
rect 19392 2388 19398 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 20622 2388 20628 2440
rect 20680 2428 20686 2440
rect 20901 2431 20959 2437
rect 20901 2428 20913 2431
rect 20680 2400 20913 2428
rect 20680 2388 20686 2400
rect 20901 2397 20913 2400
rect 20947 2397 20959 2431
rect 20901 2391 20959 2397
rect 21910 2388 21916 2440
rect 21968 2428 21974 2440
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 21968 2400 22201 2428
rect 21968 2388 21974 2400
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22646 2428 22652 2440
rect 22607 2400 22652 2428
rect 22189 2391 22247 2397
rect 22646 2388 22652 2400
rect 22704 2388 22710 2440
rect 23308 2360 23336 2536
rect 25590 2524 25596 2576
rect 25648 2564 25654 2576
rect 27448 2564 27476 2604
rect 28445 2601 28457 2604
rect 28491 2601 28503 2635
rect 28445 2595 28503 2601
rect 30282 2592 30288 2644
rect 30340 2632 30346 2644
rect 32309 2635 32367 2641
rect 32309 2632 32321 2635
rect 30340 2604 32321 2632
rect 30340 2592 30346 2604
rect 32309 2601 32321 2604
rect 32355 2601 32367 2635
rect 32309 2595 32367 2601
rect 25648 2536 27476 2564
rect 25648 2524 25654 2536
rect 27522 2524 27528 2576
rect 27580 2564 27586 2576
rect 30469 2567 30527 2573
rect 30469 2564 30481 2567
rect 27580 2536 30481 2564
rect 27580 2524 27586 2536
rect 30469 2533 30481 2536
rect 30515 2533 30527 2567
rect 30469 2527 30527 2533
rect 33229 2567 33287 2573
rect 33229 2533 33241 2567
rect 33275 2564 33287 2567
rect 34514 2564 34520 2576
rect 33275 2536 34520 2564
rect 33275 2533 33287 2536
rect 33229 2527 33287 2533
rect 34514 2524 34520 2536
rect 34572 2524 34578 2576
rect 23382 2456 23388 2508
rect 23440 2496 23446 2508
rect 34790 2496 34796 2508
rect 23440 2468 26004 2496
rect 23440 2456 23446 2468
rect 23842 2388 23848 2440
rect 23900 2428 23906 2440
rect 24765 2431 24823 2437
rect 24765 2428 24777 2431
rect 23900 2400 24777 2428
rect 23900 2388 23906 2400
rect 24765 2397 24777 2400
rect 24811 2397 24823 2431
rect 25222 2428 25228 2440
rect 25183 2400 25228 2428
rect 24765 2391 24823 2397
rect 25222 2388 25228 2400
rect 25280 2388 25286 2440
rect 25976 2437 26004 2468
rect 33704 2468 34796 2496
rect 25961 2431 26019 2437
rect 25961 2397 25973 2431
rect 26007 2397 26019 2431
rect 25961 2391 26019 2397
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27341 2431 27399 2437
rect 27341 2428 27353 2431
rect 27120 2400 27353 2428
rect 27120 2388 27126 2400
rect 27341 2397 27353 2400
rect 27387 2397 27399 2431
rect 27341 2391 27399 2397
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 28629 2431 28687 2437
rect 28629 2428 28641 2431
rect 28408 2400 28641 2428
rect 28408 2388 28414 2400
rect 28629 2397 28641 2400
rect 28675 2397 28687 2431
rect 28629 2391 28687 2397
rect 29733 2431 29791 2437
rect 29733 2397 29745 2431
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 29748 2360 29776 2391
rect 30282 2388 30288 2440
rect 30340 2428 30346 2440
rect 30653 2431 30711 2437
rect 30653 2428 30665 2431
rect 30340 2400 30665 2428
rect 30340 2388 30346 2400
rect 30653 2397 30665 2400
rect 30699 2397 30711 2431
rect 30653 2391 30711 2397
rect 31570 2388 31576 2440
rect 31628 2428 31634 2440
rect 33704 2437 33732 2468
rect 34790 2456 34796 2468
rect 34848 2456 34854 2508
rect 37734 2496 37740 2508
rect 37695 2468 37740 2496
rect 37734 2456 37740 2468
rect 37792 2456 37798 2508
rect 32493 2431 32551 2437
rect 32493 2428 32505 2431
rect 31628 2400 32505 2428
rect 31628 2388 31634 2400
rect 32493 2397 32505 2400
rect 32539 2397 32551 2431
rect 32493 2391 32551 2397
rect 33689 2431 33747 2437
rect 33689 2397 33701 2431
rect 33735 2397 33747 2431
rect 33689 2391 33747 2397
rect 33778 2388 33784 2440
rect 33836 2428 33842 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 33836 2400 34897 2428
rect 33836 2388 33842 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 36173 2431 36231 2437
rect 36173 2428 36185 2431
rect 34885 2391 34943 2397
rect 35866 2400 36185 2428
rect 3804 2332 23244 2360
rect 23308 2332 29776 2360
rect 1946 2252 1952 2304
rect 2004 2292 2010 2304
rect 2225 2295 2283 2301
rect 2225 2292 2237 2295
rect 2004 2264 2237 2292
rect 2004 2252 2010 2264
rect 2225 2261 2237 2264
rect 2271 2261 2283 2295
rect 3234 2292 3240 2304
rect 3195 2264 3240 2292
rect 2225 2255 2283 2261
rect 3234 2252 3240 2264
rect 3292 2252 3298 2304
rect 5166 2252 5172 2304
rect 5224 2292 5230 2304
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 5224 2264 5457 2292
rect 5224 2252 5230 2264
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 5445 2255 5503 2261
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 6512 2264 6745 2292
rect 6512 2252 6518 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 14826 2252 14832 2304
rect 14884 2292 14890 2304
rect 15105 2295 15163 2301
rect 15105 2292 15117 2295
rect 14884 2264 15117 2292
rect 14884 2252 14890 2264
rect 15105 2261 15117 2264
rect 15151 2261 15163 2295
rect 15105 2255 15163 2261
rect 18046 2252 18052 2304
rect 18104 2292 18110 2304
rect 18325 2295 18383 2301
rect 18325 2292 18337 2295
rect 18104 2264 18337 2292
rect 18104 2252 18110 2264
rect 18325 2261 18337 2264
rect 18371 2261 18383 2295
rect 18325 2255 18383 2261
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 22833 2295 22891 2301
rect 22833 2292 22845 2295
rect 22612 2264 22845 2292
rect 22612 2252 22618 2264
rect 22833 2261 22845 2264
rect 22879 2261 22891 2295
rect 23216 2292 23244 2332
rect 29822 2320 29828 2372
rect 29880 2360 29886 2372
rect 29880 2332 32444 2360
rect 29880 2320 29886 2332
rect 25038 2292 25044 2304
rect 23216 2264 25044 2292
rect 22833 2255 22891 2261
rect 25038 2252 25044 2264
rect 25096 2252 25102 2304
rect 25130 2252 25136 2304
rect 25188 2292 25194 2304
rect 25409 2295 25467 2301
rect 25409 2292 25421 2295
rect 25188 2264 25421 2292
rect 25188 2252 25194 2264
rect 25409 2261 25421 2264
rect 25455 2261 25467 2295
rect 25409 2255 25467 2261
rect 25774 2252 25780 2304
rect 25832 2292 25838 2304
rect 26145 2295 26203 2301
rect 26145 2292 26157 2295
rect 25832 2264 26157 2292
rect 25832 2252 25838 2264
rect 26145 2261 26157 2264
rect 26191 2261 26203 2295
rect 26145 2255 26203 2261
rect 29638 2252 29644 2304
rect 29696 2292 29702 2304
rect 29917 2295 29975 2301
rect 29917 2292 29929 2295
rect 29696 2264 29929 2292
rect 29696 2252 29702 2264
rect 29917 2261 29929 2264
rect 29963 2261 29975 2295
rect 32416 2292 32444 2332
rect 32858 2320 32864 2372
rect 32916 2360 32922 2372
rect 33045 2363 33103 2369
rect 33045 2360 33057 2363
rect 32916 2332 33057 2360
rect 32916 2320 32922 2332
rect 33045 2329 33057 2332
rect 33091 2329 33103 2363
rect 35866 2360 35894 2400
rect 36173 2397 36185 2400
rect 36219 2397 36231 2431
rect 36173 2391 36231 2397
rect 36722 2388 36728 2440
rect 36780 2428 36786 2440
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 36780 2400 37473 2428
rect 36780 2388 36786 2400
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 33045 2323 33103 2329
rect 33152 2332 35894 2360
rect 33152 2292 33180 2332
rect 32416 2264 33180 2292
rect 29917 2255 29975 2261
rect 33502 2252 33508 2304
rect 33560 2292 33566 2304
rect 33873 2295 33931 2301
rect 33873 2292 33885 2295
rect 33560 2264 33885 2292
rect 33560 2252 33566 2264
rect 33873 2261 33885 2264
rect 33919 2261 33931 2295
rect 33873 2255 33931 2261
rect 34790 2252 34796 2304
rect 34848 2292 34854 2304
rect 35069 2295 35127 2301
rect 35069 2292 35081 2295
rect 34848 2264 35081 2292
rect 34848 2252 34854 2264
rect 35069 2261 35081 2264
rect 35115 2261 35127 2295
rect 35069 2255 35127 2261
rect 36078 2252 36084 2304
rect 36136 2292 36142 2304
rect 36357 2295 36415 2301
rect 36357 2292 36369 2295
rect 36136 2264 36369 2292
rect 36136 2252 36142 2264
rect 36357 2261 36369 2264
rect 36403 2261 36415 2295
rect 36357 2255 36415 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 5258 2048 5264 2100
rect 5316 2088 5322 2100
rect 17034 2088 17040 2100
rect 5316 2060 17040 2088
rect 5316 2048 5322 2060
rect 17034 2048 17040 2060
rect 17092 2048 17098 2100
rect 24394 2048 24400 2100
rect 24452 2088 24458 2100
rect 29822 2088 29828 2100
rect 24452 2060 29828 2088
rect 24452 2048 24458 2060
rect 29822 2048 29828 2060
rect 29880 2048 29886 2100
<< via1 >>
rect 17224 37612 17276 37664
rect 21364 37612 21416 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 5908 37408 5960 37460
rect 24032 37408 24084 37460
rect 6920 37340 6972 37392
rect 8760 37340 8812 37392
rect 17224 37340 17276 37392
rect 17316 37340 17368 37392
rect 19432 37340 19484 37392
rect 21088 37340 21140 37392
rect 1584 37315 1636 37324
rect 1584 37281 1593 37315
rect 1593 37281 1627 37315
rect 1627 37281 1636 37315
rect 1584 37272 1636 37281
rect 11980 37315 12032 37324
rect 2872 37247 2924 37256
rect 2872 37213 2881 37247
rect 2881 37213 2915 37247
rect 2915 37213 2924 37247
rect 2872 37204 2924 37213
rect 3240 37204 3292 37256
rect 4620 37204 4672 37256
rect 5816 37204 5868 37256
rect 6460 37204 6512 37256
rect 8392 37204 8444 37256
rect 11980 37281 11989 37315
rect 11989 37281 12023 37315
rect 12023 37281 12032 37315
rect 11980 37272 12032 37281
rect 9956 37204 10008 37256
rect 10048 37204 10100 37256
rect 12256 37204 12308 37256
rect 4712 37136 4764 37188
rect 2780 37068 2832 37120
rect 4620 37111 4672 37120
rect 4620 37077 4629 37111
rect 4629 37077 4663 37111
rect 4663 37077 4672 37111
rect 10876 37136 10928 37188
rect 11060 37136 11112 37188
rect 14096 37204 14148 37256
rect 15200 37204 15252 37256
rect 15476 37204 15528 37256
rect 16856 37247 16908 37256
rect 16856 37213 16865 37247
rect 16865 37213 16899 37247
rect 16899 37213 16908 37247
rect 16856 37204 16908 37213
rect 17316 37204 17368 37256
rect 17500 37247 17552 37256
rect 17500 37213 17509 37247
rect 17509 37213 17543 37247
rect 17543 37213 17552 37247
rect 17500 37204 17552 37213
rect 18604 37204 18656 37256
rect 18788 37247 18840 37256
rect 18788 37213 18797 37247
rect 18797 37213 18831 37247
rect 18831 37213 18840 37247
rect 18788 37204 18840 37213
rect 19432 37247 19484 37256
rect 19432 37213 19441 37247
rect 19441 37213 19475 37247
rect 19475 37213 19484 37247
rect 20076 37247 20128 37256
rect 19432 37204 19484 37213
rect 20076 37213 20085 37247
rect 20085 37213 20119 37247
rect 20119 37213 20128 37247
rect 20076 37204 20128 37213
rect 4620 37068 4672 37077
rect 6552 37111 6604 37120
rect 6552 37077 6561 37111
rect 6561 37077 6595 37111
rect 6595 37077 6604 37111
rect 6552 37068 6604 37077
rect 7748 37111 7800 37120
rect 7748 37077 7757 37111
rect 7757 37077 7791 37111
rect 7791 37077 7800 37111
rect 7748 37068 7800 37077
rect 9036 37068 9088 37120
rect 9680 37068 9732 37120
rect 12808 37068 12860 37120
rect 13452 37068 13504 37120
rect 13728 37068 13780 37120
rect 13820 37068 13872 37120
rect 15292 37068 15344 37120
rect 16764 37068 16816 37120
rect 16948 37111 17000 37120
rect 16948 37077 16957 37111
rect 16957 37077 16991 37111
rect 16991 37077 17000 37111
rect 16948 37068 17000 37077
rect 17408 37068 17460 37120
rect 21088 37136 21140 37188
rect 19340 37068 19392 37120
rect 19984 37068 20036 37120
rect 23664 37272 23716 37324
rect 25136 37272 25188 37324
rect 21272 37204 21324 37256
rect 21456 37204 21508 37256
rect 22836 37204 22888 37256
rect 23204 37204 23256 37256
rect 23756 37204 23808 37256
rect 25872 37204 25924 37256
rect 27436 37204 27488 37256
rect 27804 37247 27856 37256
rect 27804 37213 27813 37247
rect 27813 37213 27847 37247
rect 27847 37213 27856 37247
rect 27804 37204 27856 37213
rect 28356 37272 28408 37324
rect 29644 37272 29696 37324
rect 34152 37272 34204 37324
rect 37924 37272 37976 37324
rect 30932 37204 30984 37256
rect 32864 37204 32916 37256
rect 36176 37247 36228 37256
rect 36176 37213 36185 37247
rect 36185 37213 36219 37247
rect 36219 37213 36228 37247
rect 36176 37204 36228 37213
rect 38108 37247 38160 37256
rect 38108 37213 38117 37247
rect 38117 37213 38151 37247
rect 38151 37213 38160 37247
rect 38108 37204 38160 37213
rect 21456 37068 21508 37120
rect 21916 37068 21968 37120
rect 22008 37068 22060 37120
rect 24400 37068 24452 37120
rect 24492 37068 24544 37120
rect 25504 37068 25556 37120
rect 36820 37136 36872 37188
rect 27712 37068 27764 37120
rect 28540 37111 28592 37120
rect 28540 37077 28549 37111
rect 28549 37077 28583 37111
rect 28583 37077 28592 37111
rect 28540 37068 28592 37077
rect 28908 37068 28960 37120
rect 29828 37068 29880 37120
rect 31024 37111 31076 37120
rect 31024 37077 31033 37111
rect 31033 37077 31067 37111
rect 31067 37077 31076 37111
rect 31024 37068 31076 37077
rect 32220 37068 32272 37120
rect 33048 37111 33100 37120
rect 33048 37077 33057 37111
rect 33057 37077 33091 37111
rect 33091 37077 33100 37111
rect 33048 37068 33100 37077
rect 35900 37068 35952 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 1768 36907 1820 36916
rect 1768 36873 1777 36907
rect 1777 36873 1811 36907
rect 1811 36873 1820 36907
rect 1768 36864 1820 36873
rect 20 36796 72 36848
rect 6552 36864 6604 36916
rect 1584 36771 1636 36780
rect 1584 36737 1593 36771
rect 1593 36737 1627 36771
rect 1627 36737 1636 36771
rect 1584 36728 1636 36737
rect 2964 36771 3016 36780
rect 2964 36737 2973 36771
rect 2973 36737 3007 36771
rect 3007 36737 3016 36771
rect 2964 36728 3016 36737
rect 3976 36728 4028 36780
rect 7932 36796 7984 36848
rect 13360 36796 13412 36848
rect 8300 36728 8352 36780
rect 9680 36728 9732 36780
rect 4804 36660 4856 36712
rect 8760 36660 8812 36712
rect 3056 36567 3108 36576
rect 3056 36533 3065 36567
rect 3065 36533 3099 36567
rect 3099 36533 3108 36567
rect 3056 36524 3108 36533
rect 4896 36524 4948 36576
rect 6460 36524 6512 36576
rect 6920 36524 6972 36576
rect 10876 36660 10928 36712
rect 12348 36728 12400 36780
rect 13636 36864 13688 36916
rect 13728 36796 13780 36848
rect 15384 36796 15436 36848
rect 18512 36864 18564 36916
rect 21732 36864 21784 36916
rect 21824 36864 21876 36916
rect 22008 36864 22060 36916
rect 22100 36864 22152 36916
rect 27804 36864 27856 36916
rect 28724 36864 28776 36916
rect 31024 36864 31076 36916
rect 22744 36796 22796 36848
rect 25136 36839 25188 36848
rect 14188 36771 14240 36780
rect 14188 36737 14197 36771
rect 14197 36737 14231 36771
rect 14231 36737 14240 36771
rect 14188 36728 14240 36737
rect 15200 36728 15252 36780
rect 16764 36728 16816 36780
rect 19340 36771 19392 36780
rect 19340 36737 19349 36771
rect 19349 36737 19383 36771
rect 19383 36737 19392 36771
rect 19340 36728 19392 36737
rect 19524 36728 19576 36780
rect 21088 36728 21140 36780
rect 21456 36728 21508 36780
rect 21548 36728 21600 36780
rect 22100 36728 22152 36780
rect 22928 36771 22980 36780
rect 22928 36737 22937 36771
rect 22937 36737 22971 36771
rect 22971 36737 22980 36771
rect 25136 36805 25145 36839
rect 25145 36805 25179 36839
rect 25179 36805 25188 36839
rect 25136 36796 25188 36805
rect 25228 36796 25280 36848
rect 27436 36796 27488 36848
rect 28816 36796 28868 36848
rect 39304 36864 39356 36916
rect 22928 36728 22980 36737
rect 26976 36728 27028 36780
rect 28632 36728 28684 36780
rect 38660 36796 38712 36848
rect 12716 36592 12768 36644
rect 14556 36660 14608 36712
rect 16488 36660 16540 36712
rect 14464 36592 14516 36644
rect 17592 36660 17644 36712
rect 17684 36660 17736 36712
rect 20904 36660 20956 36712
rect 25044 36703 25096 36712
rect 25044 36669 25053 36703
rect 25053 36669 25087 36703
rect 25087 36669 25096 36703
rect 25044 36660 25096 36669
rect 25228 36660 25280 36712
rect 20720 36592 20772 36644
rect 25136 36592 25188 36644
rect 27252 36592 27304 36644
rect 27528 36660 27580 36712
rect 28356 36703 28408 36712
rect 27988 36592 28040 36644
rect 12992 36567 13044 36576
rect 12992 36533 13001 36567
rect 13001 36533 13035 36567
rect 13035 36533 13044 36567
rect 12992 36524 13044 36533
rect 13636 36567 13688 36576
rect 13636 36533 13645 36567
rect 13645 36533 13679 36567
rect 13679 36533 13688 36567
rect 13636 36524 13688 36533
rect 14832 36524 14884 36576
rect 14924 36567 14976 36576
rect 14924 36533 14933 36567
rect 14933 36533 14967 36567
rect 14967 36533 14976 36567
rect 16212 36567 16264 36576
rect 14924 36524 14976 36533
rect 16212 36533 16221 36567
rect 16221 36533 16255 36567
rect 16255 36533 16264 36567
rect 16212 36524 16264 36533
rect 17132 36567 17184 36576
rect 17132 36533 17162 36567
rect 17162 36533 17184 36567
rect 17132 36524 17184 36533
rect 18604 36567 18656 36576
rect 18604 36533 18613 36567
rect 18613 36533 18647 36567
rect 18647 36533 18656 36567
rect 18604 36524 18656 36533
rect 20444 36567 20496 36576
rect 20444 36533 20453 36567
rect 20453 36533 20487 36567
rect 20487 36533 20496 36567
rect 20444 36524 20496 36533
rect 20996 36524 21048 36576
rect 21180 36524 21232 36576
rect 22468 36524 22520 36576
rect 23020 36524 23072 36576
rect 28356 36669 28365 36703
rect 28365 36669 28399 36703
rect 28399 36669 28408 36703
rect 28356 36660 28408 36669
rect 29736 36592 29788 36644
rect 38200 36567 38252 36576
rect 38200 36533 38209 36567
rect 38209 36533 38243 36567
rect 38243 36533 38252 36567
rect 38200 36524 38252 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2964 36320 3016 36372
rect 3976 36363 4028 36372
rect 3976 36329 3985 36363
rect 3985 36329 4019 36363
rect 4019 36329 4028 36363
rect 3976 36320 4028 36329
rect 4620 36320 4672 36372
rect 7932 36363 7984 36372
rect 3056 36252 3108 36304
rect 4804 36227 4856 36236
rect 4804 36193 4813 36227
rect 4813 36193 4847 36227
rect 4847 36193 4856 36227
rect 4804 36184 4856 36193
rect 5908 36184 5960 36236
rect 7932 36329 7941 36363
rect 7941 36329 7975 36363
rect 7975 36329 7984 36363
rect 7932 36320 7984 36329
rect 8484 36320 8536 36372
rect 12348 36320 12400 36372
rect 12716 36320 12768 36372
rect 14740 36320 14792 36372
rect 14832 36320 14884 36372
rect 22928 36320 22980 36372
rect 24400 36320 24452 36372
rect 17500 36252 17552 36304
rect 21180 36252 21232 36304
rect 21640 36252 21692 36304
rect 25872 36320 25924 36372
rect 27436 36320 27488 36372
rect 37188 36320 37240 36372
rect 1308 36116 1360 36168
rect 4160 36159 4212 36168
rect 2688 36023 2740 36032
rect 2688 35989 2697 36023
rect 2697 35989 2731 36023
rect 2731 35989 2740 36023
rect 2688 35980 2740 35989
rect 4160 36125 4169 36159
rect 4169 36125 4203 36159
rect 4203 36125 4212 36159
rect 4160 36116 4212 36125
rect 4896 36091 4948 36100
rect 4896 36057 4905 36091
rect 4905 36057 4939 36091
rect 4939 36057 4948 36091
rect 4896 36048 4948 36057
rect 4988 36048 5040 36100
rect 5908 35980 5960 36032
rect 6460 36091 6512 36100
rect 6460 36057 6469 36091
rect 6469 36057 6503 36091
rect 6503 36057 6512 36091
rect 7380 36091 7432 36100
rect 6460 36048 6512 36057
rect 7380 36057 7389 36091
rect 7389 36057 7423 36091
rect 7423 36057 7432 36091
rect 7380 36048 7432 36057
rect 8300 36048 8352 36100
rect 9404 36048 9456 36100
rect 9220 35980 9272 36032
rect 14464 36184 14516 36236
rect 16488 36184 16540 36236
rect 16764 36184 16816 36236
rect 20444 36184 20496 36236
rect 11704 36159 11756 36168
rect 11704 36125 11713 36159
rect 11713 36125 11747 36159
rect 11747 36125 11756 36159
rect 11704 36116 11756 36125
rect 14372 36116 14424 36168
rect 15016 36116 15068 36168
rect 15200 36159 15252 36168
rect 15200 36125 15209 36159
rect 15209 36125 15243 36159
rect 15243 36125 15252 36159
rect 15200 36116 15252 36125
rect 13728 36091 13780 36100
rect 13728 36057 13737 36091
rect 13737 36057 13771 36091
rect 13771 36057 13780 36091
rect 13728 36048 13780 36057
rect 18512 36116 18564 36168
rect 20168 36116 20220 36168
rect 21088 36116 21140 36168
rect 13912 35980 13964 36032
rect 14096 35980 14148 36032
rect 15200 35980 15252 36032
rect 15384 35980 15436 36032
rect 16028 36048 16080 36100
rect 16120 36091 16172 36100
rect 16120 36057 16129 36091
rect 16129 36057 16163 36091
rect 16163 36057 16172 36091
rect 16120 36048 16172 36057
rect 16856 35980 16908 36032
rect 17960 35980 18012 36032
rect 19984 36023 20036 36032
rect 19984 35989 19993 36023
rect 19993 35989 20027 36023
rect 20027 35989 20036 36023
rect 19984 35980 20036 35989
rect 20720 36023 20772 36032
rect 20720 35989 20729 36023
rect 20729 35989 20763 36023
rect 20763 35989 20772 36023
rect 20720 35980 20772 35989
rect 22560 36184 22612 36236
rect 22744 36184 22796 36236
rect 25504 36227 25556 36236
rect 25504 36193 25513 36227
rect 25513 36193 25547 36227
rect 25547 36193 25556 36227
rect 25504 36184 25556 36193
rect 27528 36227 27580 36236
rect 27528 36193 27537 36227
rect 27537 36193 27571 36227
rect 27571 36193 27580 36227
rect 27528 36184 27580 36193
rect 27620 36184 27672 36236
rect 21364 36091 21416 36100
rect 21364 36057 21373 36091
rect 21373 36057 21407 36091
rect 21407 36057 21416 36091
rect 21364 36048 21416 36057
rect 21640 36048 21692 36100
rect 22284 36048 22336 36100
rect 25596 36091 25648 36100
rect 21732 35980 21784 36032
rect 23480 35980 23532 36032
rect 25596 36057 25605 36091
rect 25605 36057 25639 36091
rect 25639 36057 25648 36091
rect 25596 36048 25648 36057
rect 26792 35980 26844 36032
rect 26976 35980 27028 36032
rect 27528 35980 27580 36032
rect 27988 36048 28040 36100
rect 33048 36252 33100 36304
rect 38200 36252 38252 36304
rect 36084 36116 36136 36168
rect 37280 36159 37332 36168
rect 37280 36125 37289 36159
rect 37289 36125 37323 36159
rect 37323 36125 37332 36159
rect 37280 36116 37332 36125
rect 36544 36048 36596 36100
rect 34520 35980 34572 36032
rect 38200 36023 38252 36032
rect 38200 35989 38209 36023
rect 38209 35989 38243 36023
rect 38243 35989 38252 36023
rect 38200 35980 38252 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 5908 35819 5960 35828
rect 3240 35708 3292 35760
rect 5908 35785 5917 35819
rect 5917 35785 5951 35819
rect 5951 35785 5960 35819
rect 5908 35776 5960 35785
rect 9404 35751 9456 35760
rect 9404 35717 9413 35751
rect 9413 35717 9447 35751
rect 9447 35717 9456 35751
rect 9404 35708 9456 35717
rect 6828 35640 6880 35692
rect 1584 35615 1636 35624
rect 1584 35581 1593 35615
rect 1593 35581 1627 35615
rect 1627 35581 1636 35615
rect 1584 35572 1636 35581
rect 4160 35572 4212 35624
rect 4620 35572 4672 35624
rect 5448 35572 5500 35624
rect 10508 35640 10560 35692
rect 9128 35615 9180 35624
rect 9128 35581 9137 35615
rect 9137 35581 9171 35615
rect 9171 35581 9180 35615
rect 9128 35572 9180 35581
rect 9404 35572 9456 35624
rect 10876 35572 10928 35624
rect 12440 35776 12492 35828
rect 13728 35776 13780 35828
rect 14004 35819 14056 35828
rect 14004 35785 14013 35819
rect 14013 35785 14047 35819
rect 14047 35785 14056 35819
rect 14004 35776 14056 35785
rect 15200 35776 15252 35828
rect 18696 35776 18748 35828
rect 22008 35776 22060 35828
rect 11336 35708 11388 35760
rect 15108 35708 15160 35760
rect 16304 35708 16356 35760
rect 17224 35708 17276 35760
rect 17408 35708 17460 35760
rect 19800 35708 19852 35760
rect 20352 35708 20404 35760
rect 20812 35751 20864 35760
rect 20812 35717 20821 35751
rect 20821 35717 20855 35751
rect 20855 35717 20864 35751
rect 20812 35708 20864 35717
rect 22192 35708 22244 35760
rect 22652 35708 22704 35760
rect 25136 35708 25188 35760
rect 25412 35751 25464 35760
rect 25412 35717 25421 35751
rect 25421 35717 25455 35751
rect 25455 35717 25464 35751
rect 25412 35708 25464 35717
rect 26424 35776 26476 35828
rect 28632 35776 28684 35828
rect 28816 35819 28868 35828
rect 28816 35785 28825 35819
rect 28825 35785 28859 35819
rect 28859 35785 28868 35819
rect 28816 35776 28868 35785
rect 27252 35751 27304 35760
rect 11428 35640 11480 35692
rect 13912 35683 13964 35692
rect 13912 35649 13921 35683
rect 13921 35649 13955 35683
rect 13955 35649 13964 35683
rect 13912 35640 13964 35649
rect 14096 35572 14148 35624
rect 14832 35615 14884 35624
rect 4160 35436 4212 35488
rect 7012 35436 7064 35488
rect 8208 35436 8260 35488
rect 8668 35479 8720 35488
rect 8668 35445 8677 35479
rect 8677 35445 8711 35479
rect 8711 35445 8720 35479
rect 8668 35436 8720 35445
rect 12440 35504 12492 35556
rect 14464 35504 14516 35556
rect 13452 35436 13504 35488
rect 14832 35581 14841 35615
rect 14841 35581 14875 35615
rect 14875 35581 14884 35615
rect 14832 35572 14884 35581
rect 15200 35572 15252 35624
rect 16488 35640 16540 35692
rect 18696 35640 18748 35692
rect 20168 35640 20220 35692
rect 20536 35640 20588 35692
rect 21640 35640 21692 35692
rect 21824 35640 21876 35692
rect 27252 35717 27261 35751
rect 27261 35717 27295 35751
rect 27295 35717 27304 35751
rect 27252 35708 27304 35717
rect 17132 35615 17184 35624
rect 15200 35436 15252 35488
rect 16304 35547 16356 35556
rect 16304 35513 16313 35547
rect 16313 35513 16347 35547
rect 16347 35513 16356 35547
rect 16304 35504 16356 35513
rect 16672 35436 16724 35488
rect 17132 35581 17141 35615
rect 17141 35581 17175 35615
rect 17175 35581 17184 35615
rect 17132 35572 17184 35581
rect 17224 35572 17276 35624
rect 20904 35504 20956 35556
rect 21272 35504 21324 35556
rect 23296 35572 23348 35624
rect 18880 35436 18932 35488
rect 19340 35479 19392 35488
rect 19340 35445 19349 35479
rect 19349 35445 19383 35479
rect 19383 35445 19392 35479
rect 19340 35436 19392 35445
rect 20352 35436 20404 35488
rect 22376 35436 22428 35488
rect 24768 35436 24820 35488
rect 25228 35436 25280 35488
rect 28908 35708 28960 35760
rect 25780 35504 25832 35556
rect 28448 35640 28500 35692
rect 38016 35683 38068 35692
rect 38016 35649 38025 35683
rect 38025 35649 38059 35683
rect 38059 35649 38068 35683
rect 38016 35640 38068 35649
rect 26332 35436 26384 35488
rect 27344 35436 27396 35488
rect 38200 35479 38252 35488
rect 38200 35445 38209 35479
rect 38209 35445 38243 35479
rect 38243 35445 38252 35479
rect 38200 35436 38252 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 1768 35275 1820 35284
rect 1768 35241 1777 35275
rect 1777 35241 1811 35275
rect 1811 35241 1820 35275
rect 1768 35232 1820 35241
rect 6828 35232 6880 35284
rect 10508 35232 10560 35284
rect 17408 35232 17460 35284
rect 17592 35232 17644 35284
rect 18880 35232 18932 35284
rect 21180 35232 21232 35284
rect 25596 35232 25648 35284
rect 36544 35232 36596 35284
rect 4620 35139 4672 35148
rect 4620 35105 4629 35139
rect 4629 35105 4663 35139
rect 4663 35105 4672 35139
rect 4620 35096 4672 35105
rect 2688 35028 2740 35080
rect 8484 35096 8536 35148
rect 9220 35139 9272 35148
rect 9220 35105 9229 35139
rect 9229 35105 9263 35139
rect 9263 35105 9272 35139
rect 9220 35096 9272 35105
rect 9864 35164 9916 35216
rect 11152 35164 11204 35216
rect 11612 35096 11664 35148
rect 15016 35164 15068 35216
rect 17132 35164 17184 35216
rect 18604 35164 18656 35216
rect 18696 35164 18748 35216
rect 19892 35164 19944 35216
rect 22560 35164 22612 35216
rect 23388 35164 23440 35216
rect 24492 35164 24544 35216
rect 15200 35096 15252 35148
rect 16488 35096 16540 35148
rect 16672 35096 16724 35148
rect 8576 35071 8628 35080
rect 8576 35037 8585 35071
rect 8585 35037 8619 35071
rect 8619 35037 8628 35071
rect 8576 35028 8628 35037
rect 11704 35071 11756 35080
rect 11704 35037 11713 35071
rect 11713 35037 11747 35071
rect 11747 35037 11756 35071
rect 11704 35028 11756 35037
rect 14280 35028 14332 35080
rect 17316 35096 17368 35148
rect 19708 35096 19760 35148
rect 20444 35096 20496 35148
rect 25136 35164 25188 35216
rect 26332 35139 26384 35148
rect 19800 35028 19852 35080
rect 19892 35071 19944 35080
rect 19892 35037 19901 35071
rect 19901 35037 19935 35071
rect 19935 35037 19944 35071
rect 19892 35028 19944 35037
rect 20168 35028 20220 35080
rect 26332 35105 26341 35139
rect 26341 35105 26375 35139
rect 26375 35105 26384 35139
rect 26332 35096 26384 35105
rect 26792 35096 26844 35148
rect 27068 35096 27120 35148
rect 29736 35096 29788 35148
rect 25320 35071 25372 35080
rect 25320 35037 25329 35071
rect 25329 35037 25363 35071
rect 25363 35037 25372 35071
rect 25320 35028 25372 35037
rect 4896 35003 4948 35012
rect 4896 34969 4905 35003
rect 4905 34969 4939 35003
rect 4939 34969 4948 35003
rect 4896 34960 4948 34969
rect 9312 35003 9364 35012
rect 9312 34969 9321 35003
rect 9321 34969 9355 35003
rect 9355 34969 9364 35003
rect 9312 34960 9364 34969
rect 9864 34960 9916 35012
rect 8944 34892 8996 34944
rect 9220 34892 9272 34944
rect 12072 34892 12124 34944
rect 13544 34960 13596 35012
rect 13636 34960 13688 35012
rect 15936 34960 15988 35012
rect 16120 34960 16172 35012
rect 17684 34960 17736 35012
rect 17776 35003 17828 35012
rect 17776 34969 17785 35003
rect 17785 34969 17819 35003
rect 17819 34969 17828 35003
rect 17776 34960 17828 34969
rect 14464 34892 14516 34944
rect 20076 34960 20128 35012
rect 22560 34960 22612 35012
rect 23112 35003 23164 35012
rect 23112 34969 23121 35003
rect 23121 34969 23155 35003
rect 23155 34969 23164 35003
rect 24032 35003 24084 35012
rect 23112 34960 23164 34969
rect 24032 34969 24041 35003
rect 24041 34969 24075 35003
rect 24075 34969 24084 35003
rect 24032 34960 24084 34969
rect 26424 35003 26476 35012
rect 26424 34969 26433 35003
rect 26433 34969 26467 35003
rect 26467 34969 26476 35003
rect 26424 34960 26476 34969
rect 28172 35003 28224 35012
rect 28172 34969 28181 35003
rect 28181 34969 28215 35003
rect 28215 34969 28224 35003
rect 28172 34960 28224 34969
rect 28264 35003 28316 35012
rect 28264 34969 28273 35003
rect 28273 34969 28307 35003
rect 28307 34969 28316 35003
rect 28264 34960 28316 34969
rect 18328 34892 18380 34944
rect 18880 34892 18932 34944
rect 20628 34935 20680 34944
rect 20628 34901 20637 34935
rect 20637 34901 20671 34935
rect 20671 34901 20680 34935
rect 20628 34892 20680 34901
rect 21272 34935 21324 34944
rect 21272 34901 21281 34935
rect 21281 34901 21315 34935
rect 21315 34901 21324 34935
rect 21272 34892 21324 34901
rect 21916 34935 21968 34944
rect 21916 34901 21925 34935
rect 21925 34901 21959 34935
rect 21959 34901 21968 34935
rect 21916 34892 21968 34901
rect 26516 34892 26568 34944
rect 37372 35028 37424 35080
rect 37464 34935 37516 34944
rect 37464 34901 37473 34935
rect 37473 34901 37507 34935
rect 37507 34901 37516 34935
rect 37464 34892 37516 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 1768 34595 1820 34604
rect 1768 34561 1777 34595
rect 1777 34561 1811 34595
rect 1811 34561 1820 34595
rect 1768 34552 1820 34561
rect 8576 34688 8628 34740
rect 13360 34620 13412 34672
rect 1584 34484 1636 34536
rect 8668 34552 8720 34604
rect 13544 34688 13596 34740
rect 22100 34688 22152 34740
rect 13728 34620 13780 34672
rect 17684 34620 17736 34672
rect 18052 34620 18104 34672
rect 11336 34484 11388 34536
rect 8208 34416 8260 34468
rect 15568 34552 15620 34604
rect 11704 34527 11756 34536
rect 11704 34493 11713 34527
rect 11713 34493 11747 34527
rect 11747 34493 11756 34527
rect 11704 34484 11756 34493
rect 13912 34484 13964 34536
rect 17408 34595 17460 34604
rect 17408 34561 17417 34595
rect 17417 34561 17451 34595
rect 17451 34561 17460 34595
rect 18696 34620 18748 34672
rect 18972 34620 19024 34672
rect 20260 34620 20312 34672
rect 23388 34688 23440 34740
rect 17408 34552 17460 34561
rect 19248 34595 19300 34604
rect 19248 34561 19257 34595
rect 19257 34561 19291 34595
rect 19291 34561 19300 34595
rect 19248 34552 19300 34561
rect 20536 34552 20588 34604
rect 25136 34688 25188 34740
rect 26516 34731 26568 34740
rect 26516 34697 26525 34731
rect 26525 34697 26559 34731
rect 26559 34697 26568 34731
rect 26516 34688 26568 34697
rect 28172 34688 28224 34740
rect 24768 34663 24820 34672
rect 24768 34629 24777 34663
rect 24777 34629 24811 34663
rect 24811 34629 24820 34663
rect 24768 34620 24820 34629
rect 24952 34620 25004 34672
rect 27344 34663 27396 34672
rect 22284 34552 22336 34604
rect 23940 34595 23992 34604
rect 17316 34416 17368 34468
rect 17500 34484 17552 34536
rect 18144 34484 18196 34536
rect 18696 34527 18748 34536
rect 18696 34493 18705 34527
rect 18705 34493 18739 34527
rect 18739 34493 18748 34527
rect 18696 34484 18748 34493
rect 19340 34484 19392 34536
rect 20904 34484 20956 34536
rect 19524 34416 19576 34468
rect 20720 34416 20772 34468
rect 21180 34416 21232 34468
rect 4988 34391 5040 34400
rect 4988 34357 4997 34391
rect 4997 34357 5031 34391
rect 5031 34357 5040 34391
rect 4988 34348 5040 34357
rect 6920 34348 6972 34400
rect 11796 34348 11848 34400
rect 14372 34348 14424 34400
rect 18144 34348 18196 34400
rect 18236 34348 18288 34400
rect 21272 34348 21324 34400
rect 22008 34348 22060 34400
rect 23940 34561 23949 34595
rect 23949 34561 23983 34595
rect 23983 34561 23992 34595
rect 23940 34552 23992 34561
rect 24492 34552 24544 34604
rect 27344 34629 27353 34663
rect 27353 34629 27387 34663
rect 27387 34629 27396 34663
rect 27344 34620 27396 34629
rect 36636 34552 36688 34604
rect 23388 34416 23440 34468
rect 27896 34527 27948 34536
rect 27896 34493 27905 34527
rect 27905 34493 27939 34527
rect 27939 34493 27948 34527
rect 27896 34484 27948 34493
rect 28356 34416 28408 34468
rect 24124 34348 24176 34400
rect 28724 34348 28776 34400
rect 38200 34391 38252 34400
rect 38200 34357 38209 34391
rect 38209 34357 38243 34391
rect 38243 34357 38252 34391
rect 38200 34348 38252 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 3240 34144 3292 34196
rect 6920 34144 6972 34196
rect 5448 34008 5500 34060
rect 2412 33940 2464 33992
rect 2504 33983 2556 33992
rect 2504 33949 2513 33983
rect 2513 33949 2547 33983
rect 2547 33949 2556 33983
rect 9128 34008 9180 34060
rect 9680 34051 9732 34060
rect 9680 34017 9689 34051
rect 9689 34017 9723 34051
rect 9723 34017 9732 34051
rect 9680 34008 9732 34017
rect 11704 34008 11756 34060
rect 12164 34144 12216 34196
rect 13728 34144 13780 34196
rect 15292 34144 15344 34196
rect 16856 34144 16908 34196
rect 17132 34144 17184 34196
rect 18236 34144 18288 34196
rect 18512 34144 18564 34196
rect 19064 34144 19116 34196
rect 20260 34144 20312 34196
rect 28264 34144 28316 34196
rect 36636 34187 36688 34196
rect 36636 34153 36645 34187
rect 36645 34153 36679 34187
rect 36679 34153 36688 34187
rect 36636 34144 36688 34153
rect 16580 34076 16632 34128
rect 20628 34076 20680 34128
rect 22744 34076 22796 34128
rect 23480 34076 23532 34128
rect 24032 34076 24084 34128
rect 14924 34008 14976 34060
rect 15200 34008 15252 34060
rect 17132 34008 17184 34060
rect 17408 34008 17460 34060
rect 23020 34008 23072 34060
rect 24492 34008 24544 34060
rect 27252 34051 27304 34060
rect 27252 34017 27261 34051
rect 27261 34017 27295 34051
rect 27295 34017 27304 34051
rect 27252 34008 27304 34017
rect 2504 33940 2556 33949
rect 13268 33940 13320 33992
rect 18052 33983 18104 33992
rect 18052 33949 18061 33983
rect 18061 33949 18095 33983
rect 18095 33949 18104 33983
rect 18052 33940 18104 33949
rect 18144 33983 18196 33992
rect 18144 33949 18153 33983
rect 18153 33949 18187 33983
rect 18187 33949 18196 33983
rect 18144 33940 18196 33949
rect 19432 33940 19484 33992
rect 19524 33983 19576 33992
rect 19524 33949 19533 33983
rect 19533 33949 19567 33983
rect 19567 33949 19576 33983
rect 19524 33940 19576 33949
rect 20628 33940 20680 33992
rect 5908 33915 5960 33924
rect 5908 33881 5917 33915
rect 5917 33881 5951 33915
rect 5951 33881 5960 33915
rect 5908 33872 5960 33881
rect 1768 33847 1820 33856
rect 1768 33813 1777 33847
rect 1777 33813 1811 33847
rect 1811 33813 1820 33847
rect 1768 33804 1820 33813
rect 1860 33804 1912 33856
rect 9588 33804 9640 33856
rect 11152 33847 11204 33856
rect 11152 33813 11161 33847
rect 11161 33813 11195 33847
rect 11195 33813 11204 33847
rect 11152 33804 11204 33813
rect 12256 33872 12308 33924
rect 15292 33804 15344 33856
rect 15844 33872 15896 33924
rect 16948 33872 17000 33924
rect 17040 33872 17092 33924
rect 19340 33872 19392 33924
rect 21088 33940 21140 33992
rect 23572 33940 23624 33992
rect 22744 33915 22796 33924
rect 16580 33804 16632 33856
rect 19248 33804 19300 33856
rect 22744 33881 22753 33915
rect 22753 33881 22787 33915
rect 22787 33881 22796 33915
rect 22744 33872 22796 33881
rect 24308 33940 24360 33992
rect 28356 33983 28408 33992
rect 28356 33949 28365 33983
rect 28365 33949 28399 33983
rect 28399 33949 28408 33983
rect 28356 33940 28408 33949
rect 36820 33983 36872 33992
rect 36820 33949 36829 33983
rect 36829 33949 36863 33983
rect 36863 33949 36872 33983
rect 36820 33940 36872 33949
rect 19984 33804 20036 33856
rect 20444 33804 20496 33856
rect 20904 33847 20956 33856
rect 20904 33813 20913 33847
rect 20913 33813 20947 33847
rect 20947 33813 20956 33847
rect 20904 33804 20956 33813
rect 27712 33872 27764 33924
rect 29644 33872 29696 33924
rect 28448 33847 28500 33856
rect 28448 33813 28457 33847
rect 28457 33813 28491 33847
rect 28491 33813 28500 33847
rect 28448 33804 28500 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 1584 33464 1636 33516
rect 4068 33532 4120 33584
rect 5448 33600 5500 33652
rect 5908 33600 5960 33652
rect 13268 33600 13320 33652
rect 17040 33600 17092 33652
rect 9128 33532 9180 33584
rect 11152 33532 11204 33584
rect 7472 33507 7524 33516
rect 5264 33396 5316 33448
rect 4988 33260 5040 33312
rect 7472 33473 7481 33507
rect 7481 33473 7515 33507
rect 7515 33473 7524 33507
rect 7472 33464 7524 33473
rect 8484 33396 8536 33448
rect 9036 33464 9088 33516
rect 9496 33464 9548 33516
rect 11980 33464 12032 33516
rect 11612 33396 11664 33448
rect 9036 33328 9088 33380
rect 11888 33328 11940 33380
rect 13084 33532 13136 33584
rect 17408 33532 17460 33584
rect 18788 33532 18840 33584
rect 20076 33532 20128 33584
rect 20444 33575 20496 33584
rect 20444 33541 20453 33575
rect 20453 33541 20487 33575
rect 20487 33541 20496 33575
rect 20444 33532 20496 33541
rect 23572 33600 23624 33652
rect 23848 33643 23900 33652
rect 23848 33609 23857 33643
rect 23857 33609 23891 33643
rect 23891 33609 23900 33643
rect 23848 33600 23900 33609
rect 25136 33643 25188 33652
rect 25136 33609 25145 33643
rect 25145 33609 25179 33643
rect 25179 33609 25188 33643
rect 25136 33600 25188 33609
rect 26424 33600 26476 33652
rect 22192 33532 22244 33584
rect 24124 33532 24176 33584
rect 27344 33575 27396 33584
rect 15200 33464 15252 33516
rect 16488 33464 16540 33516
rect 19156 33464 19208 33516
rect 19432 33464 19484 33516
rect 22744 33507 22796 33516
rect 22744 33473 22753 33507
rect 22753 33473 22787 33507
rect 22787 33473 22796 33507
rect 22744 33464 22796 33473
rect 27344 33541 27353 33575
rect 27353 33541 27387 33575
rect 27387 33541 27396 33575
rect 27344 33532 27396 33541
rect 27712 33600 27764 33652
rect 28540 33532 28592 33584
rect 25044 33507 25096 33516
rect 25044 33473 25053 33507
rect 25053 33473 25087 33507
rect 25087 33473 25096 33507
rect 25044 33464 25096 33473
rect 25964 33464 26016 33516
rect 29828 33532 29880 33584
rect 29644 33507 29696 33516
rect 12348 33396 12400 33448
rect 15844 33396 15896 33448
rect 17592 33396 17644 33448
rect 17684 33396 17736 33448
rect 12164 33260 12216 33312
rect 21088 33328 21140 33380
rect 27252 33439 27304 33448
rect 27252 33405 27261 33439
rect 27261 33405 27295 33439
rect 27295 33405 27304 33439
rect 27252 33396 27304 33405
rect 27896 33439 27948 33448
rect 27896 33405 27905 33439
rect 27905 33405 27939 33439
rect 27939 33405 27948 33439
rect 27896 33396 27948 33405
rect 18512 33260 18564 33312
rect 19340 33260 19392 33312
rect 19708 33260 19760 33312
rect 21824 33260 21876 33312
rect 26148 33328 26200 33380
rect 26240 33328 26292 33380
rect 29644 33473 29653 33507
rect 29653 33473 29687 33507
rect 29687 33473 29696 33507
rect 29644 33464 29696 33473
rect 23480 33260 23532 33312
rect 23940 33260 23992 33312
rect 29092 33303 29144 33312
rect 29092 33269 29101 33303
rect 29101 33269 29135 33303
rect 29135 33269 29144 33303
rect 29092 33260 29144 33269
rect 29184 33260 29236 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 2504 33056 2556 33108
rect 9680 33056 9732 33108
rect 11060 33056 11112 33108
rect 12256 33056 12308 33108
rect 14740 33056 14792 33108
rect 17684 33056 17736 33108
rect 19156 33056 19208 33108
rect 7472 32920 7524 32972
rect 5816 32852 5868 32904
rect 13452 32988 13504 33040
rect 14924 32988 14976 33040
rect 15200 32963 15252 32972
rect 10784 32852 10836 32904
rect 10876 32784 10928 32836
rect 12624 32784 12676 32836
rect 12992 32827 13044 32836
rect 12992 32793 13001 32827
rect 13001 32793 13035 32827
rect 13035 32793 13044 32827
rect 12992 32784 13044 32793
rect 11888 32716 11940 32768
rect 11980 32716 12032 32768
rect 15200 32929 15209 32963
rect 15209 32929 15243 32963
rect 15243 32929 15252 32963
rect 15200 32920 15252 32929
rect 16212 32920 16264 32972
rect 19524 32988 19576 33040
rect 17316 32920 17368 32972
rect 19616 32920 19668 32972
rect 17408 32852 17460 32904
rect 19892 33031 19944 33040
rect 19892 32997 19901 33031
rect 19901 32997 19935 33031
rect 19935 32997 19944 33031
rect 19892 32988 19944 32997
rect 23572 32988 23624 33040
rect 19984 32920 20036 32972
rect 20260 32920 20312 32972
rect 20536 32963 20588 32972
rect 20536 32929 20545 32963
rect 20545 32929 20579 32963
rect 20579 32929 20588 32963
rect 20536 32920 20588 32929
rect 21456 32920 21508 32972
rect 20076 32852 20128 32904
rect 15292 32784 15344 32836
rect 16396 32784 16448 32836
rect 17960 32784 18012 32836
rect 18604 32784 18656 32836
rect 20536 32784 20588 32836
rect 23204 32852 23256 32904
rect 24584 32895 24636 32904
rect 24584 32861 24593 32895
rect 24593 32861 24627 32895
rect 24627 32861 24636 32895
rect 24584 32852 24636 32861
rect 25044 32852 25096 32904
rect 17132 32716 17184 32768
rect 17592 32759 17644 32768
rect 17592 32725 17601 32759
rect 17601 32725 17635 32759
rect 17635 32725 17644 32759
rect 17592 32716 17644 32725
rect 17776 32716 17828 32768
rect 21088 32716 21140 32768
rect 23848 32784 23900 32836
rect 27344 33056 27396 33108
rect 26148 32920 26200 32972
rect 29092 32920 29144 32972
rect 34152 32852 34204 32904
rect 25504 32784 25556 32836
rect 26148 32827 26200 32836
rect 26148 32793 26157 32827
rect 26157 32793 26191 32827
rect 26191 32793 26200 32827
rect 26148 32784 26200 32793
rect 26056 32716 26108 32768
rect 27344 32784 27396 32836
rect 27988 32784 28040 32836
rect 28448 32716 28500 32768
rect 38200 32759 38252 32768
rect 38200 32725 38209 32759
rect 38209 32725 38243 32759
rect 38243 32725 38252 32759
rect 38200 32716 38252 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 10508 32512 10560 32564
rect 20260 32512 20312 32564
rect 20628 32512 20680 32564
rect 22192 32512 22244 32564
rect 5448 32444 5500 32496
rect 9588 32444 9640 32496
rect 11980 32487 12032 32496
rect 11980 32453 11989 32487
rect 11989 32453 12023 32487
rect 12023 32453 12032 32487
rect 11980 32444 12032 32453
rect 14740 32487 14792 32496
rect 14740 32453 14749 32487
rect 14749 32453 14783 32487
rect 14783 32453 14792 32487
rect 14740 32444 14792 32453
rect 16764 32444 16816 32496
rect 17040 32444 17092 32496
rect 17408 32444 17460 32496
rect 19616 32444 19668 32496
rect 1676 32419 1728 32428
rect 1676 32385 1685 32419
rect 1685 32385 1719 32419
rect 1719 32385 1728 32419
rect 1676 32376 1728 32385
rect 6552 32419 6604 32428
rect 6552 32385 6561 32419
rect 6561 32385 6595 32419
rect 6595 32385 6604 32419
rect 6552 32376 6604 32385
rect 9128 32376 9180 32428
rect 13820 32376 13872 32428
rect 14464 32419 14516 32428
rect 14464 32385 14473 32419
rect 14473 32385 14507 32419
rect 14507 32385 14516 32419
rect 14464 32376 14516 32385
rect 16488 32376 16540 32428
rect 9680 32308 9732 32360
rect 2228 32240 2280 32292
rect 11704 32308 11756 32360
rect 11888 32308 11940 32360
rect 12348 32308 12400 32360
rect 16212 32308 16264 32360
rect 16304 32308 16356 32360
rect 17224 32308 17276 32360
rect 17776 32308 17828 32360
rect 19064 32376 19116 32428
rect 19248 32376 19300 32428
rect 19616 32308 19668 32360
rect 19892 32351 19944 32360
rect 19892 32317 19901 32351
rect 19901 32317 19935 32351
rect 19935 32317 19944 32351
rect 19892 32308 19944 32317
rect 20260 32351 20312 32360
rect 20260 32317 20269 32351
rect 20269 32317 20303 32351
rect 20303 32317 20312 32351
rect 20260 32308 20312 32317
rect 23204 32444 23256 32496
rect 23572 32487 23624 32496
rect 23572 32453 23581 32487
rect 23581 32453 23615 32487
rect 23615 32453 23624 32487
rect 23572 32444 23624 32453
rect 25136 32487 25188 32496
rect 25136 32453 25145 32487
rect 25145 32453 25179 32487
rect 25179 32453 25188 32487
rect 25136 32444 25188 32453
rect 22008 32419 22060 32428
rect 22008 32385 22017 32419
rect 22017 32385 22051 32419
rect 22051 32385 22060 32419
rect 22008 32376 22060 32385
rect 23296 32376 23348 32428
rect 34520 32512 34572 32564
rect 27252 32487 27304 32496
rect 27252 32453 27261 32487
rect 27261 32453 27295 32487
rect 27295 32453 27304 32487
rect 27252 32444 27304 32453
rect 27436 32376 27488 32428
rect 22468 32308 22520 32360
rect 23940 32308 23992 32360
rect 5540 32172 5592 32224
rect 11060 32172 11112 32224
rect 14372 32172 14424 32224
rect 14464 32172 14516 32224
rect 15844 32172 15896 32224
rect 16212 32215 16264 32224
rect 16212 32181 16221 32215
rect 16221 32181 16255 32215
rect 16255 32181 16264 32215
rect 16212 32172 16264 32181
rect 16396 32172 16448 32224
rect 16948 32172 17000 32224
rect 17132 32172 17184 32224
rect 23020 32240 23072 32292
rect 24860 32308 24912 32360
rect 26148 32308 26200 32360
rect 28724 32376 28776 32428
rect 35440 32376 35492 32428
rect 29000 32308 29052 32360
rect 19248 32215 19300 32224
rect 19248 32181 19257 32215
rect 19257 32181 19291 32215
rect 19291 32181 19300 32215
rect 19248 32172 19300 32181
rect 19892 32172 19944 32224
rect 20812 32172 20864 32224
rect 21088 32172 21140 32224
rect 25412 32240 25464 32292
rect 29920 32240 29972 32292
rect 25228 32172 25280 32224
rect 26700 32172 26752 32224
rect 27068 32172 27120 32224
rect 28080 32172 28132 32224
rect 38200 32215 38252 32224
rect 38200 32181 38209 32215
rect 38209 32181 38243 32215
rect 38243 32181 38252 32215
rect 38200 32172 38252 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 6092 31968 6144 32020
rect 5540 31875 5592 31884
rect 5540 31841 5549 31875
rect 5549 31841 5583 31875
rect 5583 31841 5592 31875
rect 5540 31832 5592 31841
rect 1860 31764 1912 31816
rect 2320 31807 2372 31816
rect 2320 31773 2329 31807
rect 2329 31773 2363 31807
rect 2363 31773 2372 31807
rect 2320 31764 2372 31773
rect 2412 31807 2464 31816
rect 2412 31773 2421 31807
rect 2421 31773 2455 31807
rect 2455 31773 2464 31807
rect 7012 31943 7064 31952
rect 7012 31909 7021 31943
rect 7021 31909 7055 31943
rect 7055 31909 7064 31943
rect 7012 31900 7064 31909
rect 9128 31875 9180 31884
rect 9128 31841 9137 31875
rect 9137 31841 9171 31875
rect 9171 31841 9180 31875
rect 9128 31832 9180 31841
rect 11796 31832 11848 31884
rect 13820 31968 13872 32020
rect 15384 31968 15436 32020
rect 15936 31968 15988 32020
rect 19340 31968 19392 32020
rect 13820 31832 13872 31884
rect 14556 31832 14608 31884
rect 14740 31832 14792 31884
rect 16396 31832 16448 31884
rect 16672 31832 16724 31884
rect 18512 31900 18564 31952
rect 17776 31875 17828 31884
rect 17776 31841 17785 31875
rect 17785 31841 17819 31875
rect 17819 31841 17828 31875
rect 17776 31832 17828 31841
rect 17868 31832 17920 31884
rect 20260 31900 20312 31952
rect 24952 31900 25004 31952
rect 25136 31968 25188 32020
rect 29000 32011 29052 32020
rect 29000 31977 29009 32011
rect 29009 31977 29043 32011
rect 29043 31977 29052 32011
rect 29000 31968 29052 31977
rect 25412 31900 25464 31952
rect 25688 31832 25740 31884
rect 25872 31832 25924 31884
rect 2412 31764 2464 31773
rect 10508 31764 10560 31816
rect 10784 31764 10836 31816
rect 11888 31764 11940 31816
rect 17684 31764 17736 31816
rect 19064 31764 19116 31816
rect 20536 31764 20588 31816
rect 25780 31764 25832 31816
rect 27068 31875 27120 31884
rect 27068 31841 27077 31875
rect 27077 31841 27111 31875
rect 27111 31841 27120 31875
rect 27068 31832 27120 31841
rect 27620 31832 27672 31884
rect 28264 31764 28316 31816
rect 30012 31764 30064 31816
rect 11612 31696 11664 31748
rect 12256 31739 12308 31748
rect 12256 31705 12265 31739
rect 12265 31705 12299 31739
rect 12299 31705 12308 31739
rect 12256 31696 12308 31705
rect 15936 31696 15988 31748
rect 16580 31696 16632 31748
rect 23204 31696 23256 31748
rect 26056 31696 26108 31748
rect 1768 31671 1820 31680
rect 1768 31637 1777 31671
rect 1777 31637 1811 31671
rect 1811 31637 1820 31671
rect 1768 31628 1820 31637
rect 3608 31628 3660 31680
rect 13636 31628 13688 31680
rect 13728 31671 13780 31680
rect 13728 31637 13737 31671
rect 13737 31637 13771 31671
rect 13771 31637 13780 31671
rect 13728 31628 13780 31637
rect 14188 31628 14240 31680
rect 14924 31628 14976 31680
rect 17960 31628 18012 31680
rect 19340 31628 19392 31680
rect 20076 31628 20128 31680
rect 22928 31628 22980 31680
rect 25320 31628 25372 31680
rect 28172 31671 28224 31680
rect 28172 31637 28181 31671
rect 28181 31637 28215 31671
rect 28215 31637 28224 31671
rect 28172 31628 28224 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 5448 31424 5500 31476
rect 3608 31356 3660 31408
rect 5356 31356 5408 31408
rect 12072 31356 12124 31408
rect 14832 31356 14884 31408
rect 14924 31356 14976 31408
rect 17776 31356 17828 31408
rect 19616 31356 19668 31408
rect 19984 31424 20036 31476
rect 20720 31424 20772 31476
rect 23480 31424 23532 31476
rect 23756 31424 23808 31476
rect 23848 31424 23900 31476
rect 28080 31467 28132 31476
rect 28080 31433 28089 31467
rect 28089 31433 28123 31467
rect 28123 31433 28132 31467
rect 28080 31424 28132 31433
rect 11704 31331 11756 31340
rect 11704 31297 11713 31331
rect 11713 31297 11747 31331
rect 11747 31297 11756 31331
rect 11704 31288 11756 31297
rect 4712 31084 4764 31136
rect 9312 31220 9364 31272
rect 11152 31220 11204 31272
rect 11612 31220 11664 31272
rect 12072 31220 12124 31272
rect 9128 31084 9180 31136
rect 9772 31084 9824 31136
rect 14740 31288 14792 31340
rect 17500 31288 17552 31340
rect 19984 31288 20036 31340
rect 20168 31288 20220 31340
rect 24124 31356 24176 31408
rect 25320 31399 25372 31408
rect 25320 31365 25329 31399
rect 25329 31365 25363 31399
rect 25363 31365 25372 31399
rect 25320 31356 25372 31365
rect 17868 31220 17920 31272
rect 18788 31263 18840 31272
rect 18788 31229 18797 31263
rect 18797 31229 18831 31263
rect 18831 31229 18840 31263
rect 18788 31220 18840 31229
rect 19064 31220 19116 31272
rect 20720 31220 20772 31272
rect 20996 31152 21048 31204
rect 16396 31084 16448 31136
rect 16488 31084 16540 31136
rect 20536 31084 20588 31136
rect 21456 31288 21508 31340
rect 22008 31331 22060 31340
rect 22008 31297 22017 31331
rect 22017 31297 22051 31331
rect 22051 31297 22060 31331
rect 22008 31288 22060 31297
rect 23756 31288 23808 31340
rect 23848 31331 23900 31340
rect 23848 31297 23857 31331
rect 23857 31297 23891 31331
rect 23891 31297 23900 31331
rect 23848 31288 23900 31297
rect 28172 31288 28224 31340
rect 29828 31288 29880 31340
rect 30012 31331 30064 31340
rect 30012 31297 30021 31331
rect 30021 31297 30055 31331
rect 30055 31297 30064 31331
rect 30012 31288 30064 31297
rect 25228 31263 25280 31272
rect 25228 31229 25237 31263
rect 25237 31229 25271 31263
rect 25271 31229 25280 31263
rect 25228 31220 25280 31229
rect 27252 31220 27304 31272
rect 22560 31127 22612 31136
rect 22560 31093 22569 31127
rect 22569 31093 22603 31127
rect 22603 31093 22612 31127
rect 22560 31084 22612 31093
rect 24768 31084 24820 31136
rect 38016 31084 38068 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 12992 30880 13044 30932
rect 13820 30880 13872 30932
rect 20168 30880 20220 30932
rect 23756 30923 23808 30932
rect 15568 30812 15620 30864
rect 17132 30812 17184 30864
rect 5448 30744 5500 30796
rect 6092 30744 6144 30796
rect 9588 30744 9640 30796
rect 10784 30744 10836 30796
rect 15844 30787 15896 30796
rect 15844 30753 15853 30787
rect 15853 30753 15887 30787
rect 15887 30753 15896 30787
rect 15844 30744 15896 30753
rect 16580 30744 16632 30796
rect 16672 30744 16724 30796
rect 17684 30812 17736 30864
rect 23756 30889 23765 30923
rect 23765 30889 23799 30923
rect 23799 30889 23808 30923
rect 23756 30880 23808 30889
rect 2780 30676 2832 30728
rect 5356 30676 5408 30728
rect 20352 30744 20404 30796
rect 21640 30787 21692 30796
rect 21640 30753 21649 30787
rect 21649 30753 21683 30787
rect 21683 30753 21692 30787
rect 21640 30744 21692 30753
rect 22100 30787 22152 30796
rect 22100 30753 22109 30787
rect 22109 30753 22143 30787
rect 22143 30753 22152 30787
rect 22100 30744 22152 30753
rect 23020 30744 23072 30796
rect 18328 30676 18380 30728
rect 19340 30676 19392 30728
rect 4620 30540 4672 30592
rect 8484 30540 8536 30592
rect 10784 30608 10836 30660
rect 15108 30540 15160 30592
rect 17960 30608 18012 30660
rect 18052 30608 18104 30660
rect 20168 30608 20220 30660
rect 20720 30676 20772 30728
rect 21088 30676 21140 30728
rect 23112 30719 23164 30728
rect 23112 30685 23121 30719
rect 23121 30685 23155 30719
rect 23155 30685 23164 30719
rect 23112 30676 23164 30685
rect 28080 30812 28132 30864
rect 27160 30744 27212 30796
rect 29276 30676 29328 30728
rect 38292 30719 38344 30728
rect 38292 30685 38301 30719
rect 38301 30685 38335 30719
rect 38335 30685 38344 30719
rect 38292 30676 38344 30685
rect 21180 30608 21232 30660
rect 21732 30651 21784 30660
rect 21732 30617 21741 30651
rect 21741 30617 21775 30651
rect 21775 30617 21784 30651
rect 21732 30608 21784 30617
rect 17132 30540 17184 30592
rect 17776 30540 17828 30592
rect 18788 30583 18840 30592
rect 18788 30549 18797 30583
rect 18797 30549 18831 30583
rect 18831 30549 18840 30583
rect 18788 30540 18840 30549
rect 19156 30540 19208 30592
rect 20536 30540 20588 30592
rect 20996 30583 21048 30592
rect 20996 30549 21005 30583
rect 21005 30549 21039 30583
rect 21039 30549 21048 30583
rect 20996 30540 21048 30549
rect 26608 30608 26660 30660
rect 28540 30583 28592 30592
rect 28540 30549 28549 30583
rect 28549 30549 28583 30583
rect 28583 30549 28592 30583
rect 28540 30540 28592 30549
rect 38108 30583 38160 30592
rect 38108 30549 38117 30583
rect 38117 30549 38151 30583
rect 38151 30549 38160 30583
rect 38108 30540 38160 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 6184 30268 6236 30320
rect 6552 30268 6604 30320
rect 11336 30268 11388 30320
rect 11980 30268 12032 30320
rect 15844 30268 15896 30320
rect 16764 30336 16816 30388
rect 17224 30336 17276 30388
rect 18972 30336 19024 30388
rect 19340 30336 19392 30388
rect 20076 30336 20128 30388
rect 1584 30243 1636 30252
rect 1584 30209 1593 30243
rect 1593 30209 1627 30243
rect 1627 30209 1636 30243
rect 1584 30200 1636 30209
rect 6092 30200 6144 30252
rect 12348 30200 12400 30252
rect 9680 30132 9732 30184
rect 11704 30132 11756 30184
rect 12072 30132 12124 30184
rect 15292 30200 15344 30252
rect 19248 30268 19300 30320
rect 19432 30243 19484 30252
rect 19432 30209 19441 30243
rect 19441 30209 19475 30243
rect 19475 30209 19484 30243
rect 19432 30200 19484 30209
rect 19524 30200 19576 30252
rect 19984 30200 20036 30252
rect 21364 30336 21416 30388
rect 29276 30379 29328 30388
rect 20812 30268 20864 30320
rect 21272 30200 21324 30252
rect 22192 30243 22244 30252
rect 22192 30209 22201 30243
rect 22201 30209 22235 30243
rect 22235 30209 22244 30243
rect 22192 30200 22244 30209
rect 22284 30243 22336 30252
rect 22284 30209 22293 30243
rect 22293 30209 22327 30243
rect 22327 30209 22336 30243
rect 23572 30268 23624 30320
rect 24400 30268 24452 30320
rect 24952 30311 25004 30320
rect 24952 30277 24961 30311
rect 24961 30277 24995 30311
rect 24995 30277 25004 30311
rect 24952 30268 25004 30277
rect 29276 30345 29285 30379
rect 29285 30345 29319 30379
rect 29319 30345 29328 30379
rect 29276 30336 29328 30345
rect 27344 30268 27396 30320
rect 22284 30200 22336 30209
rect 16212 30132 16264 30184
rect 17224 30132 17276 30184
rect 17500 30132 17552 30184
rect 1768 30039 1820 30048
rect 1768 30005 1777 30039
rect 1777 30005 1811 30039
rect 1811 30005 1820 30039
rect 1768 29996 1820 30005
rect 7840 30039 7892 30048
rect 7840 30005 7870 30039
rect 7870 30005 7892 30039
rect 7840 29996 7892 30005
rect 9312 30039 9364 30048
rect 9312 30005 9321 30039
rect 9321 30005 9355 30039
rect 9355 30005 9364 30039
rect 9312 29996 9364 30005
rect 11980 29996 12032 30048
rect 18144 30064 18196 30116
rect 22928 30132 22980 30184
rect 23204 30132 23256 30184
rect 24216 30132 24268 30184
rect 25780 30175 25832 30184
rect 21640 30064 21692 30116
rect 25780 30141 25789 30175
rect 25789 30141 25823 30175
rect 25823 30141 25832 30175
rect 25780 30132 25832 30141
rect 27528 30200 27580 30252
rect 29736 30200 29788 30252
rect 36820 30268 36872 30320
rect 27988 30064 28040 30116
rect 14556 30039 14608 30048
rect 14556 30005 14565 30039
rect 14565 30005 14599 30039
rect 14599 30005 14608 30039
rect 14556 29996 14608 30005
rect 15200 29996 15252 30048
rect 16396 29996 16448 30048
rect 16580 29996 16632 30048
rect 18604 30039 18656 30048
rect 18604 30005 18613 30039
rect 18613 30005 18647 30039
rect 18647 30005 18656 30039
rect 18604 29996 18656 30005
rect 18696 29996 18748 30048
rect 20812 30039 20864 30048
rect 20812 30005 20821 30039
rect 20821 30005 20855 30039
rect 20855 30005 20864 30039
rect 20812 29996 20864 30005
rect 20904 29996 20956 30048
rect 23940 29996 23992 30048
rect 24308 29996 24360 30048
rect 28172 29996 28224 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 20904 29792 20956 29844
rect 21732 29792 21784 29844
rect 23940 29792 23992 29844
rect 24860 29792 24912 29844
rect 28540 29835 28592 29844
rect 28540 29801 28549 29835
rect 28549 29801 28583 29835
rect 28583 29801 28592 29835
rect 28540 29792 28592 29801
rect 29736 29835 29788 29844
rect 29736 29801 29745 29835
rect 29745 29801 29779 29835
rect 29779 29801 29788 29835
rect 29736 29792 29788 29801
rect 35440 29792 35492 29844
rect 8208 29656 8260 29708
rect 13544 29656 13596 29708
rect 15200 29656 15252 29708
rect 15844 29656 15896 29708
rect 17316 29724 17368 29776
rect 18144 29724 18196 29776
rect 18604 29724 18656 29776
rect 26332 29724 26384 29776
rect 4804 29588 4856 29640
rect 9128 29631 9180 29640
rect 9128 29597 9137 29631
rect 9137 29597 9171 29631
rect 9171 29597 9180 29631
rect 9128 29588 9180 29597
rect 11336 29631 11388 29640
rect 11336 29597 11345 29631
rect 11345 29597 11379 29631
rect 11379 29597 11388 29631
rect 11336 29588 11388 29597
rect 9404 29563 9456 29572
rect 9404 29529 9413 29563
rect 9413 29529 9447 29563
rect 9447 29529 9456 29563
rect 9404 29520 9456 29529
rect 13912 29588 13964 29640
rect 14464 29588 14516 29640
rect 15936 29588 15988 29640
rect 18052 29588 18104 29640
rect 20628 29656 20680 29708
rect 22008 29656 22060 29708
rect 24308 29656 24360 29708
rect 24768 29656 24820 29708
rect 25320 29656 25372 29708
rect 26240 29656 26292 29708
rect 18972 29588 19024 29640
rect 19524 29588 19576 29640
rect 20260 29631 20312 29640
rect 20260 29597 20269 29631
rect 20269 29597 20303 29631
rect 20303 29597 20312 29631
rect 20260 29588 20312 29597
rect 20996 29631 21048 29640
rect 20996 29597 21005 29631
rect 21005 29597 21039 29631
rect 21039 29597 21048 29631
rect 20996 29588 21048 29597
rect 21180 29588 21232 29640
rect 21640 29631 21692 29640
rect 21640 29597 21649 29631
rect 21649 29597 21683 29631
rect 21683 29597 21692 29631
rect 21640 29588 21692 29597
rect 22744 29588 22796 29640
rect 22928 29631 22980 29640
rect 22928 29597 22937 29631
rect 22937 29597 22971 29631
rect 22971 29597 22980 29631
rect 22928 29588 22980 29597
rect 26424 29631 26476 29640
rect 12072 29563 12124 29572
rect 12072 29529 12081 29563
rect 12081 29529 12115 29563
rect 12115 29529 12124 29563
rect 12072 29520 12124 29529
rect 13452 29520 13504 29572
rect 11520 29452 11572 29504
rect 21916 29520 21968 29572
rect 26424 29597 26433 29631
rect 26433 29597 26467 29631
rect 26467 29597 26476 29631
rect 26424 29588 26476 29597
rect 37464 29724 37516 29776
rect 28172 29699 28224 29708
rect 28172 29665 28181 29699
rect 28181 29665 28215 29699
rect 28215 29665 28224 29699
rect 28172 29656 28224 29665
rect 28540 29656 28592 29708
rect 28448 29588 28500 29640
rect 34612 29656 34664 29708
rect 37464 29631 37516 29640
rect 29184 29520 29236 29572
rect 17684 29452 17736 29504
rect 18052 29452 18104 29504
rect 18788 29452 18840 29504
rect 18880 29452 18932 29504
rect 21548 29452 21600 29504
rect 23020 29495 23072 29504
rect 23020 29461 23029 29495
rect 23029 29461 23063 29495
rect 23063 29461 23072 29495
rect 23020 29452 23072 29461
rect 26148 29452 26200 29504
rect 26516 29495 26568 29504
rect 26516 29461 26525 29495
rect 26525 29461 26559 29495
rect 26559 29461 26568 29495
rect 26516 29452 26568 29461
rect 27160 29495 27212 29504
rect 27160 29461 27169 29495
rect 27169 29461 27203 29495
rect 27203 29461 27212 29495
rect 27160 29452 27212 29461
rect 27528 29452 27580 29504
rect 37464 29597 37473 29631
rect 37473 29597 37507 29631
rect 37507 29597 37516 29631
rect 37464 29588 37516 29597
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 9404 29248 9456 29300
rect 13544 29248 13596 29300
rect 1768 29155 1820 29164
rect 1768 29121 1777 29155
rect 1777 29121 1811 29155
rect 1811 29121 1820 29155
rect 1768 29112 1820 29121
rect 2780 29180 2832 29232
rect 4068 29180 4120 29232
rect 6184 29180 6236 29232
rect 11520 29180 11572 29232
rect 7012 29112 7064 29164
rect 9128 29112 9180 29164
rect 4896 29044 4948 29096
rect 11612 29112 11664 29164
rect 12072 29180 12124 29232
rect 15752 29248 15804 29300
rect 16028 29248 16080 29300
rect 16488 29180 16540 29232
rect 17132 29248 17184 29300
rect 21916 29248 21968 29300
rect 17868 29180 17920 29232
rect 18144 29223 18196 29232
rect 18144 29189 18153 29223
rect 18153 29189 18187 29223
rect 18187 29189 18196 29223
rect 18144 29180 18196 29189
rect 18236 29180 18288 29232
rect 19340 29180 19392 29232
rect 11060 29087 11112 29096
rect 11060 29053 11069 29087
rect 11069 29053 11103 29087
rect 11103 29053 11112 29087
rect 11060 29044 11112 29053
rect 11428 29044 11480 29096
rect 20260 29180 20312 29232
rect 21272 29180 21324 29232
rect 24860 29248 24912 29300
rect 22928 29180 22980 29232
rect 23020 29180 23072 29232
rect 24492 29180 24544 29232
rect 14464 28976 14516 29028
rect 1860 28908 1912 28960
rect 4712 28908 4764 28960
rect 5264 28908 5316 28960
rect 10968 28908 11020 28960
rect 12072 28908 12124 28960
rect 14740 28951 14792 28960
rect 14740 28917 14770 28951
rect 14770 28917 14792 28951
rect 14740 28908 14792 28917
rect 16304 28976 16356 29028
rect 16488 28976 16540 29028
rect 18236 29044 18288 29096
rect 18420 29087 18472 29096
rect 18420 29053 18429 29087
rect 18429 29053 18463 29087
rect 18463 29053 18472 29087
rect 18420 29044 18472 29053
rect 18512 29044 18564 29096
rect 19708 29155 19760 29164
rect 19708 29121 19717 29155
rect 19717 29121 19751 29155
rect 19751 29121 19760 29155
rect 19708 29112 19760 29121
rect 19340 29044 19392 29096
rect 19708 28976 19760 29028
rect 20260 29044 20312 29096
rect 22376 29112 22428 29164
rect 20168 28976 20220 29028
rect 23940 29044 23992 29096
rect 25044 29112 25096 29164
rect 25596 29180 25648 29232
rect 32956 29180 33008 29232
rect 26976 29112 27028 29164
rect 25228 29044 25280 29096
rect 26608 29087 26660 29096
rect 26608 29053 26617 29087
rect 26617 29053 26651 29087
rect 26651 29053 26660 29087
rect 26608 29044 26660 29053
rect 27252 29087 27304 29096
rect 27252 29053 27261 29087
rect 27261 29053 27295 29087
rect 27295 29053 27304 29087
rect 27252 29044 27304 29053
rect 27988 29087 28040 29096
rect 27988 29053 27997 29087
rect 27997 29053 28031 29087
rect 28031 29053 28040 29087
rect 27988 29044 28040 29053
rect 18236 28908 18288 28960
rect 20076 28908 20128 28960
rect 27620 28976 27672 29028
rect 28448 29019 28500 29028
rect 28448 28985 28457 29019
rect 28457 28985 28491 29019
rect 28491 28985 28500 29019
rect 28448 28976 28500 28985
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 13084 28704 13136 28756
rect 9312 28636 9364 28688
rect 16212 28704 16264 28756
rect 17316 28704 17368 28756
rect 17684 28704 17736 28756
rect 11612 28611 11664 28620
rect 11612 28577 11621 28611
rect 11621 28577 11655 28611
rect 11655 28577 11664 28611
rect 11612 28568 11664 28577
rect 13636 28636 13688 28688
rect 15752 28568 15804 28620
rect 18144 28636 18196 28688
rect 20352 28704 20404 28756
rect 22652 28704 22704 28756
rect 1860 28543 1912 28552
rect 1860 28509 1869 28543
rect 1869 28509 1903 28543
rect 1903 28509 1912 28543
rect 1860 28500 1912 28509
rect 4896 28543 4948 28552
rect 4896 28509 4905 28543
rect 4905 28509 4939 28543
rect 4939 28509 4948 28543
rect 4896 28500 4948 28509
rect 18512 28500 18564 28552
rect 19524 28500 19576 28552
rect 20168 28500 20220 28552
rect 21180 28500 21232 28552
rect 21732 28543 21784 28552
rect 21732 28509 21741 28543
rect 21741 28509 21775 28543
rect 21775 28509 21784 28543
rect 21732 28500 21784 28509
rect 21916 28543 21968 28552
rect 21916 28509 21925 28543
rect 21925 28509 21959 28543
rect 21959 28509 21968 28543
rect 21916 28500 21968 28509
rect 3424 28432 3476 28484
rect 6460 28432 6512 28484
rect 11888 28475 11940 28484
rect 11888 28441 11897 28475
rect 11897 28441 11931 28475
rect 11931 28441 11940 28475
rect 11888 28432 11940 28441
rect 2136 28364 2188 28416
rect 16212 28432 16264 28484
rect 18880 28432 18932 28484
rect 19248 28432 19300 28484
rect 20536 28432 20588 28484
rect 23848 28636 23900 28688
rect 24584 28636 24636 28688
rect 25412 28704 25464 28756
rect 25964 28704 26016 28756
rect 27528 28704 27580 28756
rect 26332 28636 26384 28688
rect 23020 28611 23072 28620
rect 23020 28577 23029 28611
rect 23029 28577 23063 28611
rect 23063 28577 23072 28611
rect 23020 28568 23072 28577
rect 26240 28568 26292 28620
rect 27160 28568 27212 28620
rect 27804 28611 27856 28620
rect 27804 28577 27813 28611
rect 27813 28577 27847 28611
rect 27847 28577 27856 28611
rect 27804 28568 27856 28577
rect 24584 28543 24636 28552
rect 24584 28509 24593 28543
rect 24593 28509 24627 28543
rect 24627 28509 24636 28543
rect 24584 28500 24636 28509
rect 24952 28500 25004 28552
rect 25136 28500 25188 28552
rect 26516 28432 26568 28484
rect 17500 28364 17552 28416
rect 19156 28364 19208 28416
rect 21088 28364 21140 28416
rect 22284 28364 22336 28416
rect 22376 28364 22428 28416
rect 24768 28364 24820 28416
rect 25964 28364 26016 28416
rect 27344 28432 27396 28484
rect 27620 28475 27672 28484
rect 27620 28441 27629 28475
rect 27629 28441 27663 28475
rect 27663 28441 27672 28475
rect 27620 28432 27672 28441
rect 38108 28568 38160 28620
rect 32956 28475 33008 28484
rect 32956 28441 32965 28475
rect 32965 28441 32999 28475
rect 32999 28441 33008 28475
rect 32956 28432 33008 28441
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 9588 28160 9640 28212
rect 4988 28092 5040 28144
rect 9680 28092 9732 28144
rect 20996 28160 21048 28212
rect 21272 28203 21324 28212
rect 21272 28169 21281 28203
rect 21281 28169 21315 28203
rect 21315 28169 21324 28203
rect 21272 28160 21324 28169
rect 22284 28160 22336 28212
rect 18696 28092 18748 28144
rect 23204 28092 23256 28144
rect 23388 28092 23440 28144
rect 24952 28203 25004 28212
rect 24952 28169 24961 28203
rect 24961 28169 24995 28203
rect 24995 28169 25004 28203
rect 25596 28203 25648 28212
rect 24952 28160 25004 28169
rect 25596 28169 25605 28203
rect 25605 28169 25639 28203
rect 25639 28169 25648 28203
rect 25596 28160 25648 28169
rect 26148 28160 26200 28212
rect 10692 28024 10744 28076
rect 15844 28067 15896 28076
rect 15844 28033 15853 28067
rect 15853 28033 15887 28067
rect 15887 28033 15896 28067
rect 15844 28024 15896 28033
rect 18420 28024 18472 28076
rect 19248 28067 19300 28076
rect 19248 28033 19257 28067
rect 19257 28033 19291 28067
rect 19291 28033 19300 28067
rect 19248 28024 19300 28033
rect 20168 28024 20220 28076
rect 21180 28067 21232 28076
rect 2780 27956 2832 28008
rect 3516 27999 3568 28008
rect 3516 27965 3525 27999
rect 3525 27965 3559 27999
rect 3559 27965 3568 27999
rect 3516 27956 3568 27965
rect 3884 27956 3936 28008
rect 9588 27999 9640 28008
rect 9588 27965 9597 27999
rect 9597 27965 9631 27999
rect 9631 27965 9640 27999
rect 9588 27956 9640 27965
rect 15476 27956 15528 28008
rect 4896 27820 4948 27872
rect 8024 27820 8076 27872
rect 9404 27820 9456 27872
rect 13728 27820 13780 27872
rect 17684 27956 17736 28008
rect 18328 27956 18380 28008
rect 21180 28033 21189 28067
rect 21189 28033 21223 28067
rect 21223 28033 21232 28067
rect 21180 28024 21232 28033
rect 22652 28024 22704 28076
rect 23020 28024 23072 28076
rect 23572 28024 23624 28076
rect 24952 28024 25004 28076
rect 38292 28067 38344 28076
rect 38292 28033 38301 28067
rect 38301 28033 38335 28067
rect 38335 28033 38344 28067
rect 38292 28024 38344 28033
rect 21088 27956 21140 28008
rect 21824 27956 21876 28008
rect 22376 27999 22428 28008
rect 22376 27965 22385 27999
rect 22385 27965 22419 27999
rect 22419 27965 22428 27999
rect 22376 27956 22428 27965
rect 24308 27999 24360 28008
rect 24308 27965 24317 27999
rect 24317 27965 24351 27999
rect 24351 27965 24360 27999
rect 24308 27956 24360 27965
rect 27712 27956 27764 28008
rect 23388 27931 23440 27940
rect 23388 27897 23397 27931
rect 23397 27897 23431 27931
rect 23431 27897 23440 27931
rect 23388 27888 23440 27897
rect 27804 27931 27856 27940
rect 27804 27897 27813 27931
rect 27813 27897 27847 27931
rect 27847 27897 27856 27931
rect 27804 27888 27856 27897
rect 17960 27820 18012 27872
rect 20628 27863 20680 27872
rect 20628 27829 20637 27863
rect 20637 27829 20671 27863
rect 20671 27829 20680 27863
rect 20628 27820 20680 27829
rect 25780 27820 25832 27872
rect 35900 27820 35952 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 2872 27616 2924 27668
rect 8024 27616 8076 27668
rect 8116 27616 8168 27668
rect 10692 27616 10744 27668
rect 20628 27616 20680 27668
rect 20904 27616 20956 27668
rect 24952 27616 25004 27668
rect 7104 27548 7156 27600
rect 9588 27548 9640 27600
rect 4896 27480 4948 27532
rect 9680 27480 9732 27532
rect 1584 27455 1636 27464
rect 1584 27421 1593 27455
rect 1593 27421 1627 27455
rect 1627 27421 1636 27455
rect 1584 27412 1636 27421
rect 18144 27548 18196 27600
rect 22192 27548 22244 27600
rect 24032 27548 24084 27600
rect 11796 27480 11848 27532
rect 12348 27523 12400 27532
rect 12348 27489 12357 27523
rect 12357 27489 12391 27523
rect 12391 27489 12400 27523
rect 12348 27480 12400 27489
rect 21916 27480 21968 27532
rect 20628 27412 20680 27464
rect 21640 27412 21692 27464
rect 5632 27344 5684 27396
rect 1768 27319 1820 27328
rect 1768 27285 1777 27319
rect 1777 27285 1811 27319
rect 1811 27285 1820 27319
rect 1768 27276 1820 27285
rect 12348 27344 12400 27396
rect 13176 27276 13228 27328
rect 17684 27387 17736 27396
rect 17684 27353 17693 27387
rect 17693 27353 17727 27387
rect 17727 27353 17736 27387
rect 17684 27344 17736 27353
rect 18696 27344 18748 27396
rect 18972 27276 19024 27328
rect 19800 27387 19852 27396
rect 19800 27353 19809 27387
rect 19809 27353 19843 27387
rect 19843 27353 19852 27387
rect 19800 27344 19852 27353
rect 20536 27344 20588 27396
rect 26700 27548 26752 27600
rect 27988 27548 28040 27600
rect 26240 27480 26292 27532
rect 23572 27455 23624 27464
rect 23572 27421 23581 27455
rect 23581 27421 23615 27455
rect 23615 27421 23624 27455
rect 23572 27412 23624 27421
rect 24584 27455 24636 27464
rect 24584 27421 24593 27455
rect 24593 27421 24627 27455
rect 24627 27421 24636 27455
rect 24584 27412 24636 27421
rect 29736 27455 29788 27464
rect 29736 27421 29745 27455
rect 29745 27421 29779 27455
rect 29779 27421 29788 27455
rect 29736 27412 29788 27421
rect 38016 27455 38068 27464
rect 38016 27421 38025 27455
rect 38025 27421 38059 27455
rect 38059 27421 38068 27455
rect 38016 27412 38068 27421
rect 20904 27276 20956 27328
rect 21272 27319 21324 27328
rect 21272 27285 21281 27319
rect 21281 27285 21315 27319
rect 21315 27285 21324 27319
rect 21272 27276 21324 27285
rect 24676 27319 24728 27328
rect 24676 27285 24685 27319
rect 24685 27285 24719 27319
rect 24719 27285 24728 27319
rect 24676 27276 24728 27285
rect 25964 27387 26016 27396
rect 25964 27353 25973 27387
rect 25973 27353 26007 27387
rect 26007 27353 26016 27387
rect 26884 27387 26936 27396
rect 25964 27344 26016 27353
rect 26884 27353 26893 27387
rect 26893 27353 26927 27387
rect 26927 27353 26936 27387
rect 26884 27344 26936 27353
rect 28080 27276 28132 27328
rect 38200 27319 38252 27328
rect 38200 27285 38209 27319
rect 38209 27285 38243 27319
rect 38243 27285 38252 27319
rect 38200 27276 38252 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 2320 27072 2372 27124
rect 3332 27072 3384 27124
rect 4620 27004 4672 27056
rect 16488 27072 16540 27124
rect 11336 27004 11388 27056
rect 13728 27004 13780 27056
rect 17684 27072 17736 27124
rect 20904 27115 20956 27124
rect 18144 27047 18196 27056
rect 1768 26979 1820 26988
rect 1768 26945 1777 26979
rect 1777 26945 1811 26979
rect 1811 26945 1820 26979
rect 1768 26936 1820 26945
rect 16488 26936 16540 26988
rect 18144 27013 18153 27047
rect 18153 27013 18187 27047
rect 18187 27013 18196 27047
rect 18144 27004 18196 27013
rect 20904 27081 20913 27115
rect 20913 27081 20947 27115
rect 20947 27081 20956 27115
rect 20904 27072 20956 27081
rect 21732 27072 21784 27124
rect 23572 27072 23624 27124
rect 24032 27072 24084 27124
rect 24400 27072 24452 27124
rect 24584 27072 24636 27124
rect 34152 27115 34204 27124
rect 22468 27004 22520 27056
rect 23848 27047 23900 27056
rect 23848 27013 23857 27047
rect 23857 27013 23891 27047
rect 23891 27013 23900 27047
rect 23848 27004 23900 27013
rect 17592 26936 17644 26988
rect 4620 26868 4672 26920
rect 4896 26868 4948 26920
rect 5080 26868 5132 26920
rect 5724 26868 5776 26920
rect 6736 26868 6788 26920
rect 7564 26868 7616 26920
rect 11612 26868 11664 26920
rect 17684 26868 17736 26920
rect 19432 26936 19484 26988
rect 19984 26936 20036 26988
rect 20168 26979 20220 26988
rect 20168 26945 20177 26979
rect 20177 26945 20211 26979
rect 20211 26945 20220 26979
rect 20168 26936 20220 26945
rect 21640 26936 21692 26988
rect 23388 26936 23440 26988
rect 24400 26936 24452 26988
rect 34152 27081 34161 27115
rect 34161 27081 34195 27115
rect 34195 27081 34204 27115
rect 34152 27072 34204 27081
rect 34612 27004 34664 27056
rect 25780 26979 25832 26988
rect 25780 26945 25789 26979
rect 25789 26945 25823 26979
rect 25823 26945 25832 26979
rect 25780 26936 25832 26945
rect 28356 26979 28408 26988
rect 28356 26945 28365 26979
rect 28365 26945 28399 26979
rect 28399 26945 28408 26979
rect 28356 26936 28408 26945
rect 4620 26732 4672 26784
rect 5172 26732 5224 26784
rect 22100 26868 22152 26920
rect 22468 26868 22520 26920
rect 31944 26936 31996 26988
rect 12072 26732 12124 26784
rect 17132 26732 17184 26784
rect 19984 26732 20036 26784
rect 21088 26800 21140 26852
rect 23112 26800 23164 26852
rect 38108 26868 38160 26920
rect 24768 26800 24820 26852
rect 27712 26800 27764 26852
rect 24492 26732 24544 26784
rect 25044 26775 25096 26784
rect 25044 26741 25053 26775
rect 25053 26741 25087 26775
rect 25087 26741 25096 26775
rect 25044 26732 25096 26741
rect 27896 26732 27948 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 2964 26528 3016 26580
rect 3516 26528 3568 26580
rect 8944 26528 8996 26580
rect 17776 26528 17828 26580
rect 17868 26528 17920 26580
rect 20352 26528 20404 26580
rect 21088 26528 21140 26580
rect 23848 26528 23900 26580
rect 25964 26528 26016 26580
rect 13268 26460 13320 26512
rect 19432 26460 19484 26512
rect 19524 26460 19576 26512
rect 24676 26460 24728 26512
rect 2136 26435 2188 26444
rect 2136 26401 2145 26435
rect 2145 26401 2179 26435
rect 2179 26401 2188 26435
rect 2136 26392 2188 26401
rect 7012 26435 7064 26444
rect 7012 26401 7021 26435
rect 7021 26401 7055 26435
rect 7055 26401 7064 26435
rect 7012 26392 7064 26401
rect 6736 26367 6788 26376
rect 6736 26333 6745 26367
rect 6745 26333 6779 26367
rect 6779 26333 6788 26367
rect 6736 26324 6788 26333
rect 11612 26324 11664 26376
rect 11704 26324 11756 26376
rect 21272 26392 21324 26444
rect 29460 26528 29512 26580
rect 31944 26571 31996 26580
rect 31944 26537 31953 26571
rect 31953 26537 31987 26571
rect 31987 26537 31996 26571
rect 31944 26528 31996 26537
rect 38108 26571 38160 26580
rect 38108 26537 38117 26571
rect 38117 26537 38151 26571
rect 38151 26537 38160 26571
rect 38108 26528 38160 26537
rect 27804 26460 27856 26512
rect 33232 26460 33284 26512
rect 15752 26367 15804 26376
rect 15752 26333 15761 26367
rect 15761 26333 15795 26367
rect 15795 26333 15804 26367
rect 15752 26324 15804 26333
rect 17132 26324 17184 26376
rect 17592 26324 17644 26376
rect 3056 26256 3108 26308
rect 5080 26256 5132 26308
rect 8392 26256 8444 26308
rect 12256 26299 12308 26308
rect 12256 26265 12265 26299
rect 12265 26265 12299 26299
rect 12299 26265 12308 26299
rect 12256 26256 12308 26265
rect 17776 26299 17828 26308
rect 17776 26265 17785 26299
rect 17785 26265 17819 26299
rect 17819 26265 17828 26299
rect 17776 26256 17828 26265
rect 19064 26324 19116 26376
rect 19248 26324 19300 26376
rect 19524 26299 19576 26308
rect 12992 26188 13044 26240
rect 15108 26188 15160 26240
rect 18880 26188 18932 26240
rect 19524 26265 19533 26299
rect 19533 26265 19567 26299
rect 19567 26265 19576 26299
rect 19524 26256 19576 26265
rect 20812 26324 20864 26376
rect 23112 26367 23164 26376
rect 23112 26333 23121 26367
rect 23121 26333 23155 26367
rect 23155 26333 23164 26367
rect 23112 26324 23164 26333
rect 23756 26367 23808 26376
rect 23756 26333 23765 26367
rect 23765 26333 23799 26367
rect 23799 26333 23808 26367
rect 23756 26324 23808 26333
rect 24400 26324 24452 26376
rect 20536 26299 20588 26308
rect 20536 26265 20545 26299
rect 20545 26265 20579 26299
rect 20579 26265 20588 26299
rect 20536 26256 20588 26265
rect 21088 26256 21140 26308
rect 21456 26188 21508 26240
rect 23296 26188 23348 26240
rect 25412 26324 25464 26376
rect 25872 26324 25924 26376
rect 31852 26367 31904 26376
rect 31852 26333 31861 26367
rect 31861 26333 31895 26367
rect 31895 26333 31904 26367
rect 31852 26324 31904 26333
rect 38292 26367 38344 26376
rect 38292 26333 38301 26367
rect 38301 26333 38335 26367
rect 38335 26333 38344 26367
rect 38292 26324 38344 26333
rect 26424 26299 26476 26308
rect 26424 26265 26433 26299
rect 26433 26265 26467 26299
rect 26467 26265 26476 26299
rect 26424 26256 26476 26265
rect 32588 26299 32640 26308
rect 32588 26265 32597 26299
rect 32597 26265 32631 26299
rect 32631 26265 32640 26299
rect 32588 26256 32640 26265
rect 33232 26299 33284 26308
rect 33232 26265 33241 26299
rect 33241 26265 33275 26299
rect 33275 26265 33284 26299
rect 33232 26256 33284 26265
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 3056 26027 3108 26036
rect 3056 25993 3065 26027
rect 3065 25993 3099 26027
rect 3099 25993 3108 26027
rect 3056 25984 3108 25993
rect 1952 25916 2004 25968
rect 17960 25984 18012 26036
rect 18144 25984 18196 26036
rect 21180 25984 21232 26036
rect 26424 25984 26476 26036
rect 32588 25984 32640 26036
rect 14648 25916 14700 25968
rect 17224 25916 17276 25968
rect 19156 25916 19208 25968
rect 2964 25891 3016 25900
rect 2964 25857 2973 25891
rect 2973 25857 3007 25891
rect 3007 25857 3016 25891
rect 2964 25848 3016 25857
rect 4988 25848 5040 25900
rect 7932 25891 7984 25900
rect 7932 25857 7941 25891
rect 7941 25857 7975 25891
rect 7975 25857 7984 25891
rect 7932 25848 7984 25857
rect 3884 25823 3936 25832
rect 3884 25789 3893 25823
rect 3893 25789 3927 25823
rect 3927 25789 3936 25823
rect 3884 25780 3936 25789
rect 6736 25780 6788 25832
rect 8392 25780 8444 25832
rect 9128 25780 9180 25832
rect 10968 25780 11020 25832
rect 11704 25823 11756 25832
rect 11704 25789 11713 25823
rect 11713 25789 11747 25823
rect 11747 25789 11756 25823
rect 11704 25780 11756 25789
rect 10876 25712 10928 25764
rect 4620 25644 4672 25696
rect 11060 25687 11112 25696
rect 11060 25653 11069 25687
rect 11069 25653 11103 25687
rect 11103 25653 11112 25687
rect 11060 25644 11112 25653
rect 14832 25848 14884 25900
rect 16764 25848 16816 25900
rect 18604 25848 18656 25900
rect 22376 25916 22428 25968
rect 13452 25823 13504 25832
rect 13452 25789 13461 25823
rect 13461 25789 13495 25823
rect 13495 25789 13504 25823
rect 13452 25780 13504 25789
rect 15752 25780 15804 25832
rect 17132 25823 17184 25832
rect 17132 25789 17141 25823
rect 17141 25789 17175 25823
rect 17175 25789 17184 25823
rect 17132 25780 17184 25789
rect 17224 25780 17276 25832
rect 20168 25848 20220 25900
rect 21180 25848 21232 25900
rect 21364 25848 21416 25900
rect 21640 25848 21692 25900
rect 22192 25848 22244 25900
rect 23296 25848 23348 25900
rect 23940 25848 23992 25900
rect 28264 25891 28316 25900
rect 28264 25857 28273 25891
rect 28273 25857 28307 25891
rect 28307 25857 28316 25891
rect 28264 25848 28316 25857
rect 20812 25780 20864 25832
rect 29920 25823 29972 25832
rect 29920 25789 29929 25823
rect 29929 25789 29963 25823
rect 29963 25789 29972 25823
rect 29920 25780 29972 25789
rect 30104 25823 30156 25832
rect 30104 25789 30113 25823
rect 30113 25789 30147 25823
rect 30147 25789 30156 25823
rect 30104 25780 30156 25789
rect 30472 25780 30524 25832
rect 16672 25644 16724 25696
rect 20996 25712 21048 25764
rect 29092 25712 29144 25764
rect 29184 25712 29236 25764
rect 18604 25687 18656 25696
rect 18604 25653 18613 25687
rect 18613 25653 18647 25687
rect 18647 25653 18656 25687
rect 18604 25644 18656 25653
rect 19432 25644 19484 25696
rect 21364 25687 21416 25696
rect 21364 25653 21373 25687
rect 21373 25653 21407 25687
rect 21407 25653 21416 25687
rect 21364 25644 21416 25653
rect 28540 25644 28592 25696
rect 31852 25712 31904 25764
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 10876 25483 10928 25492
rect 10876 25449 10885 25483
rect 10885 25449 10919 25483
rect 10919 25449 10928 25483
rect 10876 25440 10928 25449
rect 6736 25347 6788 25356
rect 6736 25313 6745 25347
rect 6745 25313 6779 25347
rect 6779 25313 6788 25347
rect 6736 25304 6788 25313
rect 9128 25347 9180 25356
rect 1676 25279 1728 25288
rect 1676 25245 1685 25279
rect 1685 25245 1719 25279
rect 1719 25245 1728 25279
rect 1676 25236 1728 25245
rect 2688 25168 2740 25220
rect 8024 25168 8076 25220
rect 3976 25100 4028 25152
rect 8668 25100 8720 25152
rect 9128 25313 9137 25347
rect 9137 25313 9171 25347
rect 9171 25313 9180 25347
rect 9128 25304 9180 25313
rect 13728 25440 13780 25492
rect 14832 25304 14884 25356
rect 10508 25236 10560 25288
rect 11796 25279 11848 25288
rect 11796 25245 11805 25279
rect 11805 25245 11839 25279
rect 11839 25245 11848 25279
rect 11796 25236 11848 25245
rect 19340 25440 19392 25492
rect 19524 25440 19576 25492
rect 20536 25440 20588 25492
rect 22560 25440 22612 25492
rect 30104 25440 30156 25492
rect 16580 25304 16632 25356
rect 25872 25372 25924 25424
rect 20076 25304 20128 25356
rect 15384 25236 15436 25288
rect 15752 25236 15804 25288
rect 18788 25236 18840 25288
rect 19340 25236 19392 25288
rect 19984 25236 20036 25288
rect 20444 25236 20496 25288
rect 20628 25279 20680 25288
rect 20628 25245 20637 25279
rect 20637 25245 20671 25279
rect 20671 25245 20680 25279
rect 20628 25236 20680 25245
rect 20720 25236 20772 25288
rect 21456 25279 21508 25288
rect 21456 25245 21465 25279
rect 21465 25245 21499 25279
rect 21499 25245 21508 25279
rect 21456 25236 21508 25245
rect 22928 25236 22980 25288
rect 23756 25236 23808 25288
rect 27160 25236 27212 25288
rect 28540 25279 28592 25288
rect 28540 25245 28549 25279
rect 28549 25245 28583 25279
rect 28583 25245 28592 25279
rect 28540 25236 28592 25245
rect 29184 25279 29236 25288
rect 29184 25245 29193 25279
rect 29193 25245 29227 25279
rect 29227 25245 29236 25279
rect 29184 25236 29236 25245
rect 9680 25100 9732 25152
rect 15752 25100 15804 25152
rect 18604 25100 18656 25152
rect 18880 25100 18932 25152
rect 20720 25143 20772 25152
rect 20720 25109 20729 25143
rect 20729 25109 20763 25143
rect 20763 25109 20772 25143
rect 20720 25100 20772 25109
rect 28632 25100 28684 25152
rect 36176 25168 36228 25220
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 1768 24803 1820 24812
rect 1768 24769 1777 24803
rect 1777 24769 1811 24803
rect 1811 24769 1820 24803
rect 1768 24760 1820 24769
rect 6920 24760 6972 24812
rect 8392 24803 8444 24812
rect 8392 24769 8401 24803
rect 8401 24769 8435 24803
rect 8435 24769 8444 24803
rect 8392 24760 8444 24769
rect 9772 24760 9824 24812
rect 4620 24692 4672 24744
rect 6000 24692 6052 24744
rect 1216 24556 1268 24608
rect 4068 24556 4120 24608
rect 4712 24556 4764 24608
rect 6920 24556 6972 24608
rect 7932 24556 7984 24608
rect 11336 24692 11388 24744
rect 11796 24692 11848 24744
rect 13176 24803 13228 24812
rect 13176 24769 13185 24803
rect 13185 24769 13219 24803
rect 13219 24769 13228 24803
rect 13176 24760 13228 24769
rect 15476 24760 15528 24812
rect 15752 24896 15804 24948
rect 29184 24896 29236 24948
rect 16764 24828 16816 24880
rect 18972 24828 19024 24880
rect 27528 24871 27580 24880
rect 10140 24667 10192 24676
rect 10140 24633 10149 24667
rect 10149 24633 10183 24667
rect 10183 24633 10192 24667
rect 10140 24624 10192 24633
rect 12992 24624 13044 24676
rect 10600 24556 10652 24608
rect 17224 24735 17276 24744
rect 16764 24624 16816 24676
rect 17224 24701 17233 24735
rect 17233 24701 17267 24735
rect 17267 24701 17276 24735
rect 17224 24692 17276 24701
rect 17592 24692 17644 24744
rect 18880 24760 18932 24812
rect 19984 24760 20036 24812
rect 20168 24760 20220 24812
rect 20628 24760 20680 24812
rect 20996 24803 21048 24812
rect 20996 24769 21005 24803
rect 21005 24769 21039 24803
rect 21039 24769 21048 24803
rect 20996 24760 21048 24769
rect 20812 24692 20864 24744
rect 21916 24692 21968 24744
rect 27528 24837 27537 24871
rect 27537 24837 27571 24871
rect 27571 24837 27580 24871
rect 27528 24828 27580 24837
rect 23940 24803 23992 24812
rect 23940 24769 23949 24803
rect 23949 24769 23983 24803
rect 23983 24769 23992 24803
rect 23940 24760 23992 24769
rect 25412 24760 25464 24812
rect 27160 24760 27212 24812
rect 29092 24760 29144 24812
rect 17132 24624 17184 24676
rect 17408 24624 17460 24676
rect 21364 24624 21416 24676
rect 21640 24624 21692 24676
rect 22928 24624 22980 24676
rect 15384 24556 15436 24608
rect 15936 24556 15988 24608
rect 18236 24556 18288 24608
rect 20536 24556 20588 24608
rect 22008 24556 22060 24608
rect 27252 24692 27304 24744
rect 28356 24735 28408 24744
rect 28356 24701 28365 24735
rect 28365 24701 28399 24735
rect 28399 24701 28408 24735
rect 28356 24692 28408 24701
rect 28540 24692 28592 24744
rect 23848 24624 23900 24676
rect 24216 24556 24268 24608
rect 25596 24556 25648 24608
rect 38200 24599 38252 24608
rect 38200 24565 38209 24599
rect 38209 24565 38243 24599
rect 38243 24565 38252 24599
rect 38200 24556 38252 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 2688 24352 2740 24404
rect 6460 24352 6512 24404
rect 9588 24352 9640 24404
rect 9772 24352 9824 24404
rect 13912 24352 13964 24404
rect 4252 24216 4304 24268
rect 4620 24216 4672 24268
rect 7748 24284 7800 24336
rect 11704 24284 11756 24336
rect 12992 24284 13044 24336
rect 21732 24352 21784 24404
rect 25412 24352 25464 24404
rect 22008 24284 22060 24336
rect 22652 24284 22704 24336
rect 29644 24352 29696 24404
rect 6276 24148 6328 24200
rect 18880 24216 18932 24268
rect 19340 24216 19392 24268
rect 19432 24216 19484 24268
rect 15384 24191 15436 24200
rect 15384 24157 15393 24191
rect 15393 24157 15427 24191
rect 15427 24157 15436 24191
rect 15384 24148 15436 24157
rect 21548 24148 21600 24200
rect 22836 24259 22888 24268
rect 22836 24225 22845 24259
rect 22845 24225 22879 24259
rect 22879 24225 22888 24259
rect 22836 24216 22888 24225
rect 23204 24216 23256 24268
rect 29736 24284 29788 24336
rect 28540 24259 28592 24268
rect 28540 24225 28549 24259
rect 28549 24225 28583 24259
rect 28583 24225 28592 24259
rect 28540 24216 28592 24225
rect 29920 24216 29972 24268
rect 1124 24080 1176 24132
rect 1952 24123 2004 24132
rect 1952 24089 1961 24123
rect 1961 24089 1995 24123
rect 1995 24089 2004 24123
rect 1952 24080 2004 24089
rect 2504 24080 2556 24132
rect 4528 24080 4580 24132
rect 4804 24080 4856 24132
rect 6368 24080 6420 24132
rect 9220 24080 9272 24132
rect 2044 24012 2096 24064
rect 8208 24055 8260 24064
rect 8208 24021 8217 24055
rect 8217 24021 8251 24055
rect 8251 24021 8260 24055
rect 8208 24012 8260 24021
rect 9588 24012 9640 24064
rect 10784 24012 10836 24064
rect 13728 24012 13780 24064
rect 19432 24080 19484 24132
rect 20628 24080 20680 24132
rect 34704 24148 34756 24200
rect 16580 24012 16632 24064
rect 17132 24055 17184 24064
rect 17132 24021 17141 24055
rect 17141 24021 17175 24055
rect 17175 24021 17184 24055
rect 17132 24012 17184 24021
rect 18144 24012 18196 24064
rect 19984 24012 20036 24064
rect 21732 24012 21784 24064
rect 27712 24080 27764 24132
rect 28632 24123 28684 24132
rect 28632 24089 28641 24123
rect 28641 24089 28675 24123
rect 28675 24089 28684 24123
rect 28632 24080 28684 24089
rect 28908 24012 28960 24064
rect 38200 24055 38252 24064
rect 38200 24021 38209 24055
rect 38209 24021 38243 24055
rect 38243 24021 38252 24055
rect 38200 24012 38252 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 4712 23808 4764 23860
rect 5172 23808 5224 23860
rect 4160 23740 4212 23792
rect 7748 23740 7800 23792
rect 2780 23672 2832 23724
rect 4252 23715 4304 23724
rect 4252 23681 4261 23715
rect 4261 23681 4295 23715
rect 4295 23681 4304 23715
rect 4252 23672 4304 23681
rect 11796 23808 11848 23860
rect 16488 23808 16540 23860
rect 8668 23740 8720 23792
rect 11336 23740 11388 23792
rect 18144 23783 18196 23792
rect 13728 23672 13780 23724
rect 16856 23715 16908 23724
rect 16856 23681 16865 23715
rect 16865 23681 16899 23715
rect 16899 23681 16908 23715
rect 16856 23672 16908 23681
rect 2872 23604 2924 23656
rect 1492 23468 1544 23520
rect 2688 23468 2740 23520
rect 6368 23468 6420 23520
rect 10140 23604 10192 23656
rect 15384 23604 15436 23656
rect 18144 23749 18153 23783
rect 18153 23749 18187 23783
rect 18187 23749 18196 23783
rect 18144 23740 18196 23749
rect 24032 23808 24084 23860
rect 20168 23740 20220 23792
rect 21456 23740 21508 23792
rect 23020 23740 23072 23792
rect 25596 23783 25648 23792
rect 25596 23749 25605 23783
rect 25605 23749 25639 23783
rect 25639 23749 25648 23783
rect 25596 23740 25648 23749
rect 29092 23808 29144 23860
rect 27896 23740 27948 23792
rect 19156 23672 19208 23724
rect 20812 23672 20864 23724
rect 22652 23715 22704 23724
rect 22652 23681 22661 23715
rect 22661 23681 22695 23715
rect 22695 23681 22704 23715
rect 22652 23672 22704 23681
rect 24124 23672 24176 23724
rect 21640 23604 21692 23656
rect 27528 23672 27580 23724
rect 33232 23672 33284 23724
rect 26884 23604 26936 23656
rect 27988 23647 28040 23656
rect 27988 23613 27997 23647
rect 27997 23613 28031 23647
rect 28031 23613 28040 23647
rect 27988 23604 28040 23613
rect 29828 23604 29880 23656
rect 14740 23536 14792 23588
rect 17224 23536 17276 23588
rect 20168 23536 20220 23588
rect 22192 23536 22244 23588
rect 22468 23536 22520 23588
rect 29920 23536 29972 23588
rect 13912 23468 13964 23520
rect 20352 23468 20404 23520
rect 24400 23511 24452 23520
rect 24400 23477 24409 23511
rect 24409 23477 24443 23511
rect 24443 23477 24452 23511
rect 24400 23468 24452 23477
rect 34428 23468 34480 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 4620 23128 4672 23180
rect 5080 23128 5132 23180
rect 15200 23264 15252 23316
rect 12992 23196 13044 23248
rect 20720 23264 20772 23316
rect 28448 23264 28500 23316
rect 16948 23196 17000 23248
rect 20536 23196 20588 23248
rect 1584 23060 1636 23112
rect 9312 23060 9364 23112
rect 14832 23128 14884 23180
rect 25596 23128 25648 23180
rect 29828 23171 29880 23180
rect 29828 23137 29837 23171
rect 29837 23137 29871 23171
rect 29871 23137 29880 23171
rect 29828 23128 29880 23137
rect 12348 23060 12400 23112
rect 12808 23060 12860 23112
rect 12900 23060 12952 23112
rect 15292 23060 15344 23112
rect 15476 23103 15528 23112
rect 15476 23069 15485 23103
rect 15485 23069 15519 23103
rect 15519 23069 15528 23103
rect 15476 23060 15528 23069
rect 18236 23060 18288 23112
rect 18972 23060 19024 23112
rect 20352 23060 20404 23112
rect 21548 23060 21600 23112
rect 26148 23103 26200 23112
rect 26148 23069 26157 23103
rect 26157 23069 26191 23103
rect 26191 23069 26200 23103
rect 26148 23060 26200 23069
rect 28172 23103 28224 23112
rect 28172 23069 28181 23103
rect 28181 23069 28215 23103
rect 28215 23069 28224 23103
rect 28172 23060 28224 23069
rect 28724 23060 28776 23112
rect 2044 22992 2096 23044
rect 3792 22992 3844 23044
rect 6736 22992 6788 23044
rect 12716 22992 12768 23044
rect 13544 22992 13596 23044
rect 15752 23035 15804 23044
rect 15752 23001 15761 23035
rect 15761 23001 15795 23035
rect 15795 23001 15804 23035
rect 15752 22992 15804 23001
rect 17408 22992 17460 23044
rect 18512 22992 18564 23044
rect 29920 23035 29972 23044
rect 29920 23001 29929 23035
rect 29929 23001 29963 23035
rect 29963 23001 29972 23035
rect 29920 22992 29972 23001
rect 32956 22992 33008 23044
rect 35992 22992 36044 23044
rect 3424 22967 3476 22976
rect 3424 22933 3433 22967
rect 3433 22933 3467 22967
rect 3467 22933 3476 22967
rect 3424 22924 3476 22933
rect 7564 22924 7616 22976
rect 12256 22967 12308 22976
rect 12256 22933 12265 22967
rect 12265 22933 12299 22967
rect 12299 22933 12308 22967
rect 12256 22924 12308 22933
rect 17224 22924 17276 22976
rect 17684 22924 17736 22976
rect 28448 22924 28500 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 7472 22720 7524 22772
rect 1400 22652 1452 22704
rect 3148 22652 3200 22704
rect 5540 22652 5592 22704
rect 1584 22559 1636 22568
rect 1584 22525 1593 22559
rect 1593 22525 1627 22559
rect 1627 22525 1636 22559
rect 1584 22516 1636 22525
rect 6828 22516 6880 22568
rect 4712 22380 4764 22432
rect 6000 22423 6052 22432
rect 6000 22389 6009 22423
rect 6009 22389 6043 22423
rect 6043 22389 6052 22423
rect 6000 22380 6052 22389
rect 11060 22720 11112 22772
rect 15476 22720 15528 22772
rect 17224 22720 17276 22772
rect 24584 22720 24636 22772
rect 26148 22720 26200 22772
rect 28724 22763 28776 22772
rect 28724 22729 28733 22763
rect 28733 22729 28767 22763
rect 28767 22729 28776 22763
rect 28724 22720 28776 22729
rect 34704 22720 34756 22772
rect 15292 22695 15344 22704
rect 15292 22661 15301 22695
rect 15301 22661 15335 22695
rect 15335 22661 15344 22695
rect 15292 22652 15344 22661
rect 16580 22652 16632 22704
rect 9128 22516 9180 22568
rect 14648 22584 14700 22636
rect 11888 22448 11940 22500
rect 13268 22448 13320 22500
rect 11428 22380 11480 22432
rect 11520 22380 11572 22432
rect 13176 22380 13228 22432
rect 13544 22559 13596 22568
rect 13544 22525 13553 22559
rect 13553 22525 13587 22559
rect 13587 22525 13596 22559
rect 17040 22584 17092 22636
rect 18512 22627 18564 22636
rect 18512 22593 18521 22627
rect 18521 22593 18555 22627
rect 18555 22593 18564 22627
rect 18512 22584 18564 22593
rect 18972 22584 19024 22636
rect 20628 22652 20680 22704
rect 22192 22695 22244 22704
rect 22192 22661 22201 22695
rect 22201 22661 22235 22695
rect 22235 22661 22244 22695
rect 22192 22652 22244 22661
rect 27804 22652 27856 22704
rect 28080 22652 28132 22704
rect 20812 22584 20864 22636
rect 13544 22516 13596 22525
rect 17776 22516 17828 22568
rect 18420 22516 18472 22568
rect 19156 22516 19208 22568
rect 19616 22559 19668 22568
rect 19616 22525 19625 22559
rect 19625 22525 19659 22559
rect 19659 22525 19668 22559
rect 19616 22516 19668 22525
rect 20536 22516 20588 22568
rect 25964 22627 26016 22636
rect 25964 22593 25973 22627
rect 25973 22593 26007 22627
rect 26007 22593 26016 22627
rect 25964 22584 26016 22593
rect 28908 22627 28960 22636
rect 19984 22448 20036 22500
rect 20996 22516 21048 22568
rect 25780 22516 25832 22568
rect 28908 22593 28917 22627
rect 28917 22593 28951 22627
rect 28951 22593 28960 22627
rect 28908 22584 28960 22593
rect 31300 22627 31352 22636
rect 31300 22593 31309 22627
rect 31309 22593 31343 22627
rect 31343 22593 31352 22627
rect 31300 22584 31352 22593
rect 34428 22627 34480 22636
rect 34428 22593 34437 22627
rect 34437 22593 34471 22627
rect 34471 22593 34480 22627
rect 34428 22584 34480 22593
rect 28080 22516 28132 22568
rect 22468 22448 22520 22500
rect 22652 22491 22704 22500
rect 22652 22457 22661 22491
rect 22661 22457 22695 22491
rect 22695 22457 22704 22491
rect 22652 22448 22704 22457
rect 38200 22491 38252 22500
rect 38200 22457 38209 22491
rect 38209 22457 38243 22491
rect 38243 22457 38252 22491
rect 38200 22448 38252 22457
rect 15844 22380 15896 22432
rect 16488 22380 16540 22432
rect 19340 22380 19392 22432
rect 20168 22380 20220 22432
rect 22100 22380 22152 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 8300 22176 8352 22228
rect 11520 22176 11572 22228
rect 12900 22176 12952 22228
rect 13268 22176 13320 22228
rect 25136 22176 25188 22228
rect 25780 22176 25832 22228
rect 25964 22176 26016 22228
rect 5080 22083 5132 22092
rect 5080 22049 5089 22083
rect 5089 22049 5123 22083
rect 5123 22049 5132 22083
rect 5080 22040 5132 22049
rect 6828 22083 6880 22092
rect 6828 22049 6837 22083
rect 6837 22049 6871 22083
rect 6871 22049 6880 22083
rect 6828 22040 6880 22049
rect 10784 22040 10836 22092
rect 1676 21947 1728 21956
rect 1676 21913 1685 21947
rect 1685 21913 1719 21947
rect 1719 21913 1728 21947
rect 1676 21904 1728 21913
rect 3332 21904 3384 21956
rect 5264 21904 5316 21956
rect 9312 21904 9364 21956
rect 9680 21904 9732 21956
rect 4896 21836 4948 21888
rect 5080 21836 5132 21888
rect 7748 21836 7800 21888
rect 11796 22040 11848 22092
rect 13176 22108 13228 22160
rect 16304 22108 16356 22160
rect 16488 22108 16540 22160
rect 19616 22108 19668 22160
rect 22100 22108 22152 22160
rect 22284 22108 22336 22160
rect 13636 22083 13688 22092
rect 13636 22049 13645 22083
rect 13645 22049 13679 22083
rect 13679 22049 13688 22083
rect 13636 22040 13688 22049
rect 17316 22040 17368 22092
rect 19064 22040 19116 22092
rect 13820 21972 13872 22024
rect 18512 21972 18564 22024
rect 18972 21972 19024 22024
rect 20352 22040 20404 22092
rect 20812 22040 20864 22092
rect 21364 22083 21416 22092
rect 21364 22049 21373 22083
rect 21373 22049 21407 22083
rect 21407 22049 21416 22083
rect 21364 22040 21416 22049
rect 23756 22040 23808 22092
rect 12624 21904 12676 21956
rect 11796 21836 11848 21888
rect 20536 21972 20588 22024
rect 22468 21972 22520 22024
rect 23204 22015 23256 22024
rect 23204 21981 23213 22015
rect 23213 21981 23247 22015
rect 23247 21981 23256 22015
rect 23204 21972 23256 21981
rect 23848 22015 23900 22024
rect 23848 21981 23857 22015
rect 23857 21981 23891 22015
rect 23891 21981 23900 22015
rect 23848 21972 23900 21981
rect 26332 22015 26384 22024
rect 26332 21981 26341 22015
rect 26341 21981 26375 22015
rect 26375 21981 26384 22015
rect 26332 21972 26384 21981
rect 31300 22040 31352 22092
rect 20260 21904 20312 21956
rect 21088 21947 21140 21956
rect 21088 21913 21097 21947
rect 21097 21913 21131 21947
rect 21131 21913 21140 21947
rect 21088 21904 21140 21913
rect 24676 21947 24728 21956
rect 24676 21913 24685 21947
rect 24685 21913 24719 21947
rect 24719 21913 24728 21947
rect 24676 21904 24728 21913
rect 17960 21836 18012 21888
rect 20628 21836 20680 21888
rect 25320 21904 25372 21956
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 5816 21632 5868 21684
rect 6920 21564 6972 21616
rect 7748 21607 7800 21616
rect 7748 21573 7757 21607
rect 7757 21573 7791 21607
rect 7791 21573 7800 21607
rect 7748 21564 7800 21573
rect 10140 21632 10192 21684
rect 16212 21632 16264 21684
rect 16120 21564 16172 21616
rect 20812 21632 20864 21684
rect 21088 21632 21140 21684
rect 21364 21632 21416 21684
rect 23756 21632 23808 21684
rect 24032 21675 24084 21684
rect 24032 21641 24041 21675
rect 24041 21641 24075 21675
rect 24075 21641 24084 21675
rect 24032 21632 24084 21641
rect 38016 21632 38068 21684
rect 16396 21564 16448 21616
rect 23204 21564 23256 21616
rect 15844 21496 15896 21548
rect 18328 21539 18380 21548
rect 18328 21505 18337 21539
rect 18337 21505 18371 21539
rect 18371 21505 18380 21539
rect 18328 21496 18380 21505
rect 18972 21539 19024 21548
rect 18972 21505 18981 21539
rect 18981 21505 19015 21539
rect 19015 21505 19024 21539
rect 18972 21496 19024 21505
rect 20352 21496 20404 21548
rect 20536 21496 20588 21548
rect 23296 21539 23348 21548
rect 4804 21428 4856 21480
rect 6552 21428 6604 21480
rect 9128 21428 9180 21480
rect 14464 21471 14516 21480
rect 14464 21437 14473 21471
rect 14473 21437 14507 21471
rect 14507 21437 14516 21471
rect 14464 21428 14516 21437
rect 15200 21428 15252 21480
rect 18880 21428 18932 21480
rect 19064 21428 19116 21480
rect 19248 21428 19300 21480
rect 20720 21428 20772 21480
rect 23296 21505 23305 21539
rect 23305 21505 23339 21539
rect 23339 21505 23348 21539
rect 23296 21496 23348 21505
rect 24584 21539 24636 21548
rect 22284 21471 22336 21480
rect 22284 21437 22293 21471
rect 22293 21437 22327 21471
rect 22327 21437 22336 21471
rect 22284 21428 22336 21437
rect 24584 21505 24593 21539
rect 24593 21505 24627 21539
rect 24627 21505 24636 21539
rect 24584 21496 24636 21505
rect 28080 21539 28132 21548
rect 28080 21505 28089 21539
rect 28089 21505 28123 21539
rect 28123 21505 28132 21539
rect 28080 21496 28132 21505
rect 35900 21564 35952 21616
rect 31668 21539 31720 21548
rect 31668 21505 31677 21539
rect 31677 21505 31711 21539
rect 31711 21505 31720 21539
rect 31668 21496 31720 21505
rect 37832 21496 37884 21548
rect 26240 21428 26292 21480
rect 22744 21360 22796 21412
rect 28448 21403 28500 21412
rect 28448 21369 28457 21403
rect 28457 21369 28491 21403
rect 28491 21369 28500 21403
rect 28448 21360 28500 21369
rect 9772 21292 9824 21344
rect 17132 21292 17184 21344
rect 18420 21335 18472 21344
rect 18420 21301 18429 21335
rect 18429 21301 18463 21335
rect 18463 21301 18472 21335
rect 18420 21292 18472 21301
rect 19708 21292 19760 21344
rect 20812 21292 20864 21344
rect 20904 21292 20956 21344
rect 23664 21292 23716 21344
rect 27436 21292 27488 21344
rect 38200 21335 38252 21344
rect 38200 21301 38209 21335
rect 38209 21301 38243 21335
rect 38243 21301 38252 21335
rect 38200 21292 38252 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 8208 21088 8260 21140
rect 12440 21088 12492 21140
rect 15844 21088 15896 21140
rect 28080 21088 28132 21140
rect 29092 21131 29144 21140
rect 29092 21097 29101 21131
rect 29101 21097 29135 21131
rect 29135 21097 29144 21131
rect 29092 21088 29144 21097
rect 6552 20952 6604 21004
rect 6644 20952 6696 21004
rect 9128 20995 9180 21004
rect 9128 20961 9137 20995
rect 9137 20961 9171 20995
rect 9171 20961 9180 20995
rect 9128 20952 9180 20961
rect 14832 21020 14884 21072
rect 16764 21020 16816 21072
rect 20720 21020 20772 21072
rect 9036 20884 9088 20936
rect 1676 20859 1728 20868
rect 1676 20825 1685 20859
rect 1685 20825 1719 20859
rect 1719 20825 1728 20859
rect 1676 20816 1728 20825
rect 10416 20816 10468 20868
rect 12164 20748 12216 20800
rect 20168 20952 20220 21004
rect 20536 20995 20588 21004
rect 20536 20961 20545 20995
rect 20545 20961 20579 20995
rect 20579 20961 20588 20995
rect 27344 21020 27396 21072
rect 20536 20952 20588 20961
rect 23756 20952 23808 21004
rect 24676 20952 24728 21004
rect 27436 20952 27488 21004
rect 14464 20884 14516 20936
rect 17776 20884 17828 20936
rect 21180 20927 21232 20936
rect 21180 20893 21189 20927
rect 21189 20893 21223 20927
rect 21223 20893 21232 20927
rect 21180 20884 21232 20893
rect 28632 20884 28684 20936
rect 38108 21020 38160 21072
rect 30932 20927 30984 20936
rect 15108 20816 15160 20868
rect 17684 20816 17736 20868
rect 19708 20859 19760 20868
rect 17040 20748 17092 20800
rect 17132 20748 17184 20800
rect 18328 20748 18380 20800
rect 19708 20825 19717 20859
rect 19717 20825 19751 20859
rect 19751 20825 19760 20859
rect 19708 20816 19760 20825
rect 20628 20816 20680 20868
rect 23020 20816 23072 20868
rect 23112 20816 23164 20868
rect 21180 20748 21232 20800
rect 22284 20748 22336 20800
rect 23572 20748 23624 20800
rect 24860 20748 24912 20800
rect 26792 20816 26844 20868
rect 28448 20816 28500 20868
rect 30932 20893 30941 20927
rect 30941 20893 30975 20927
rect 30975 20893 30984 20927
rect 30932 20884 30984 20893
rect 31760 20927 31812 20936
rect 31760 20893 31769 20927
rect 31769 20893 31803 20927
rect 31803 20893 31812 20927
rect 31760 20884 31812 20893
rect 37188 20884 37240 20936
rect 37740 20927 37792 20936
rect 37740 20893 37749 20927
rect 37749 20893 37783 20927
rect 37783 20893 37792 20927
rect 37740 20884 37792 20893
rect 31852 20816 31904 20868
rect 31576 20791 31628 20800
rect 31576 20757 31585 20791
rect 31585 20757 31619 20791
rect 31619 20757 31628 20791
rect 31576 20748 31628 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 10692 20544 10744 20596
rect 17960 20544 18012 20596
rect 20444 20544 20496 20596
rect 20628 20544 20680 20596
rect 22192 20544 22244 20596
rect 26240 20544 26292 20596
rect 26792 20544 26844 20596
rect 31760 20544 31812 20596
rect 6920 20476 6972 20528
rect 1768 20451 1820 20460
rect 1768 20417 1777 20451
rect 1777 20417 1811 20451
rect 1811 20417 1820 20451
rect 1768 20408 1820 20417
rect 7472 20408 7524 20460
rect 9128 20476 9180 20528
rect 17408 20476 17460 20528
rect 17040 20408 17092 20460
rect 18144 20408 18196 20460
rect 20352 20451 20404 20460
rect 20352 20417 20361 20451
rect 20361 20417 20395 20451
rect 20395 20417 20404 20451
rect 20352 20408 20404 20417
rect 1584 20340 1636 20392
rect 3056 20340 3108 20392
rect 11980 20340 12032 20392
rect 15108 20340 15160 20392
rect 17500 20340 17552 20392
rect 20628 20383 20680 20392
rect 20628 20349 20637 20383
rect 20637 20349 20671 20383
rect 20671 20349 20680 20383
rect 20628 20340 20680 20349
rect 21916 20340 21968 20392
rect 26332 20408 26384 20460
rect 27252 20451 27304 20460
rect 27252 20417 27261 20451
rect 27261 20417 27295 20451
rect 27295 20417 27304 20451
rect 27252 20408 27304 20417
rect 27896 20451 27948 20460
rect 27896 20417 27897 20451
rect 27897 20417 27931 20451
rect 27931 20417 27948 20451
rect 27896 20408 27948 20417
rect 28632 20451 28684 20460
rect 28632 20417 28641 20451
rect 28641 20417 28675 20451
rect 28675 20417 28684 20451
rect 28632 20408 28684 20417
rect 30932 20408 30984 20460
rect 31576 20408 31628 20460
rect 31852 20408 31904 20460
rect 31116 20383 31168 20392
rect 31116 20349 31125 20383
rect 31125 20349 31159 20383
rect 31159 20349 31168 20383
rect 31116 20340 31168 20349
rect 9404 20272 9456 20324
rect 2136 20204 2188 20256
rect 5356 20204 5408 20256
rect 5632 20204 5684 20256
rect 8484 20204 8536 20256
rect 27528 20204 27580 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 3332 20000 3384 20052
rect 19984 20000 20036 20052
rect 3976 19864 4028 19916
rect 1584 19796 1636 19848
rect 5540 19728 5592 19780
rect 6552 19864 6604 19916
rect 11980 19864 12032 19916
rect 9312 19839 9364 19848
rect 9312 19805 9321 19839
rect 9321 19805 9355 19839
rect 9355 19805 9364 19839
rect 9312 19796 9364 19805
rect 10692 19796 10744 19848
rect 14556 19932 14608 19984
rect 21916 19932 21968 19984
rect 26884 20000 26936 20052
rect 27712 19932 27764 19984
rect 27436 19907 27488 19916
rect 6092 19728 6144 19780
rect 6920 19728 6972 19780
rect 4160 19660 4212 19712
rect 7748 19728 7800 19780
rect 9588 19771 9640 19780
rect 9588 19737 9597 19771
rect 9597 19737 9631 19771
rect 9631 19737 9640 19771
rect 9588 19728 9640 19737
rect 10968 19728 11020 19780
rect 7656 19703 7708 19712
rect 7656 19669 7665 19703
rect 7665 19669 7699 19703
rect 7699 19669 7708 19703
rect 7656 19660 7708 19669
rect 8116 19660 8168 19712
rect 11060 19703 11112 19712
rect 11060 19669 11069 19703
rect 11069 19669 11103 19703
rect 11103 19669 11112 19703
rect 11060 19660 11112 19669
rect 12164 19728 12216 19780
rect 15108 19839 15160 19848
rect 15108 19805 15117 19839
rect 15117 19805 15151 19839
rect 15151 19805 15160 19839
rect 15108 19796 15160 19805
rect 15384 19771 15436 19780
rect 15384 19737 15393 19771
rect 15393 19737 15427 19771
rect 15427 19737 15436 19771
rect 15384 19728 15436 19737
rect 16764 19728 16816 19780
rect 17960 19728 18012 19780
rect 16856 19703 16908 19712
rect 16856 19669 16865 19703
rect 16865 19669 16899 19703
rect 16899 19669 16908 19703
rect 16856 19660 16908 19669
rect 20352 19660 20404 19712
rect 27436 19873 27445 19907
rect 27445 19873 27479 19907
rect 27479 19873 27488 19907
rect 27436 19864 27488 19873
rect 27804 19907 27856 19916
rect 27804 19873 27813 19907
rect 27813 19873 27847 19907
rect 27847 19873 27856 19907
rect 27804 19864 27856 19873
rect 31116 19864 31168 19916
rect 23204 19796 23256 19848
rect 22560 19771 22612 19780
rect 22560 19737 22569 19771
rect 22569 19737 22603 19771
rect 22603 19737 22612 19771
rect 22560 19728 22612 19737
rect 27528 19771 27580 19780
rect 27528 19737 27537 19771
rect 27537 19737 27571 19771
rect 27571 19737 27580 19771
rect 27528 19728 27580 19737
rect 21640 19660 21692 19712
rect 23572 19660 23624 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 3240 19456 3292 19508
rect 4252 19456 4304 19508
rect 5356 19456 5408 19508
rect 4160 19388 4212 19440
rect 4068 19320 4120 19372
rect 4804 19388 4856 19440
rect 8208 19456 8260 19508
rect 9588 19456 9640 19508
rect 11520 19456 11572 19508
rect 11704 19456 11756 19508
rect 16764 19456 16816 19508
rect 31668 19456 31720 19508
rect 38108 19499 38160 19508
rect 38108 19465 38117 19499
rect 38117 19465 38151 19499
rect 38151 19465 38160 19499
rect 38108 19456 38160 19465
rect 7380 19388 7432 19440
rect 9772 19388 9824 19440
rect 9956 19388 10008 19440
rect 11060 19388 11112 19440
rect 12348 19388 12400 19440
rect 6552 19363 6604 19372
rect 6552 19329 6561 19363
rect 6561 19329 6595 19363
rect 6595 19329 6604 19363
rect 6552 19320 6604 19329
rect 8116 19320 8168 19372
rect 1584 19295 1636 19304
rect 1584 19261 1593 19295
rect 1593 19261 1627 19295
rect 1627 19261 1636 19295
rect 1584 19252 1636 19261
rect 4160 19252 4212 19304
rect 5724 19252 5776 19304
rect 7196 19252 7248 19304
rect 9128 19320 9180 19372
rect 12256 19320 12308 19372
rect 15108 19388 15160 19440
rect 16488 19388 16540 19440
rect 22192 19431 22244 19440
rect 22192 19397 22201 19431
rect 22201 19397 22235 19431
rect 22235 19397 22244 19431
rect 22192 19388 22244 19397
rect 23020 19388 23072 19440
rect 27896 19388 27948 19440
rect 19984 19320 20036 19372
rect 21916 19320 21968 19372
rect 23572 19363 23624 19372
rect 23572 19329 23581 19363
rect 23581 19329 23615 19363
rect 23615 19329 23624 19363
rect 23572 19320 23624 19329
rect 30840 19363 30892 19372
rect 30840 19329 30849 19363
rect 30849 19329 30883 19363
rect 30883 19329 30892 19363
rect 30840 19320 30892 19329
rect 31852 19320 31904 19372
rect 33324 19320 33376 19372
rect 38292 19363 38344 19372
rect 38292 19329 38301 19363
rect 38301 19329 38335 19363
rect 38335 19329 38344 19363
rect 38292 19320 38344 19329
rect 10140 19252 10192 19304
rect 11060 19252 11112 19304
rect 17592 19252 17644 19304
rect 4712 19116 4764 19168
rect 7564 19116 7616 19168
rect 8116 19116 8168 19168
rect 8300 19159 8352 19168
rect 8300 19125 8309 19159
rect 8309 19125 8343 19159
rect 8343 19125 8352 19159
rect 8300 19116 8352 19125
rect 16212 19184 16264 19236
rect 19708 19184 19760 19236
rect 20720 19184 20772 19236
rect 14464 19116 14516 19168
rect 16396 19116 16448 19168
rect 19524 19116 19576 19168
rect 20260 19116 20312 19168
rect 22100 19116 22152 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1308 18912 1360 18964
rect 6644 18912 6696 18964
rect 10324 18912 10376 18964
rect 4436 18844 4488 18896
rect 5724 18844 5776 18896
rect 6460 18844 6512 18896
rect 3056 18776 3108 18828
rect 4804 18776 4856 18828
rect 6552 18776 6604 18828
rect 8484 18844 8536 18896
rect 8392 18776 8444 18828
rect 18052 18912 18104 18964
rect 19984 18912 20036 18964
rect 17684 18844 17736 18896
rect 21640 18844 21692 18896
rect 22192 18912 22244 18964
rect 11980 18819 12032 18828
rect 11980 18785 11989 18819
rect 11989 18785 12023 18819
rect 12023 18785 12032 18819
rect 11980 18776 12032 18785
rect 1584 18751 1636 18760
rect 1584 18717 1593 18751
rect 1593 18717 1627 18751
rect 1627 18717 1636 18751
rect 1584 18708 1636 18717
rect 4160 18708 4212 18760
rect 8760 18708 8812 18760
rect 9312 18708 9364 18760
rect 14464 18776 14516 18828
rect 4712 18683 4764 18692
rect 4712 18649 4721 18683
rect 4721 18649 4755 18683
rect 4755 18649 4764 18683
rect 4712 18640 4764 18649
rect 5724 18640 5776 18692
rect 7564 18640 7616 18692
rect 6644 18572 6696 18624
rect 7288 18572 7340 18624
rect 9404 18640 9456 18692
rect 9864 18683 9916 18692
rect 9864 18649 9873 18683
rect 9873 18649 9907 18683
rect 9907 18649 9916 18683
rect 9864 18640 9916 18649
rect 8852 18572 8904 18624
rect 14372 18640 14424 18692
rect 15108 18708 15160 18760
rect 17500 18708 17552 18760
rect 22928 18751 22980 18760
rect 22928 18717 22937 18751
rect 22937 18717 22971 18751
rect 22971 18717 22980 18751
rect 22928 18708 22980 18717
rect 23388 18708 23440 18760
rect 27252 18708 27304 18760
rect 15568 18640 15620 18692
rect 11336 18615 11388 18624
rect 11336 18581 11345 18615
rect 11345 18581 11379 18615
rect 11379 18581 11388 18615
rect 11336 18572 11388 18581
rect 13176 18572 13228 18624
rect 17684 18640 17736 18692
rect 19524 18683 19576 18692
rect 19524 18649 19533 18683
rect 19533 18649 19567 18683
rect 19567 18649 19576 18683
rect 19524 18640 19576 18649
rect 16396 18572 16448 18624
rect 19340 18572 19392 18624
rect 20076 18640 20128 18692
rect 20536 18683 20588 18692
rect 20536 18649 20545 18683
rect 20545 18649 20579 18683
rect 20579 18649 20588 18683
rect 20536 18640 20588 18649
rect 21088 18683 21140 18692
rect 21088 18649 21097 18683
rect 21097 18649 21131 18683
rect 21131 18649 21140 18683
rect 21088 18640 21140 18649
rect 19708 18572 19760 18624
rect 30380 18615 30432 18624
rect 30380 18581 30389 18615
rect 30389 18581 30423 18615
rect 30423 18581 30432 18615
rect 30380 18572 30432 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 3700 18368 3752 18420
rect 4712 18368 4764 18420
rect 7196 18368 7248 18420
rect 1676 18343 1728 18352
rect 1676 18309 1685 18343
rect 1685 18309 1719 18343
rect 1719 18309 1728 18343
rect 1676 18300 1728 18309
rect 3332 18300 3384 18352
rect 4436 18300 4488 18352
rect 6552 18300 6604 18352
rect 2596 18207 2648 18216
rect 2596 18173 2605 18207
rect 2605 18173 2639 18207
rect 2639 18173 2648 18207
rect 2596 18164 2648 18173
rect 2872 18207 2924 18216
rect 2872 18173 2881 18207
rect 2881 18173 2915 18207
rect 2915 18173 2924 18207
rect 2872 18164 2924 18173
rect 3424 18164 3476 18216
rect 7564 18232 7616 18284
rect 7840 18232 7892 18284
rect 8760 18300 8812 18352
rect 9404 18368 9456 18420
rect 11336 18368 11388 18420
rect 25688 18368 25740 18420
rect 29460 18368 29512 18420
rect 10324 18300 10376 18352
rect 12808 18300 12860 18352
rect 15476 18300 15528 18352
rect 16764 18300 16816 18352
rect 18696 18300 18748 18352
rect 19892 18343 19944 18352
rect 19892 18309 19901 18343
rect 19901 18309 19935 18343
rect 19935 18309 19944 18343
rect 19892 18300 19944 18309
rect 20996 18300 21048 18352
rect 23848 18343 23900 18352
rect 23848 18309 23857 18343
rect 23857 18309 23891 18343
rect 23891 18309 23900 18343
rect 23848 18300 23900 18309
rect 15108 18232 15160 18284
rect 33324 18275 33376 18284
rect 4712 18164 4764 18216
rect 33324 18241 33333 18275
rect 33333 18241 33367 18275
rect 33367 18241 33376 18275
rect 33324 18232 33376 18241
rect 11336 18164 11388 18216
rect 12900 18207 12952 18216
rect 12900 18173 12909 18207
rect 12909 18173 12943 18207
rect 12943 18173 12952 18207
rect 12900 18164 12952 18173
rect 13176 18207 13228 18216
rect 13176 18173 13185 18207
rect 13185 18173 13219 18207
rect 13219 18173 13228 18207
rect 13176 18164 13228 18173
rect 15384 18164 15436 18216
rect 15568 18164 15620 18216
rect 16212 18164 16264 18216
rect 17132 18207 17184 18216
rect 17132 18173 17141 18207
rect 17141 18173 17175 18207
rect 17175 18173 17184 18207
rect 17132 18164 17184 18173
rect 17500 18164 17552 18216
rect 18144 18164 18196 18216
rect 18604 18207 18656 18216
rect 18604 18173 18613 18207
rect 18613 18173 18647 18207
rect 18647 18173 18656 18207
rect 18604 18164 18656 18173
rect 23756 18207 23808 18216
rect 5356 18096 5408 18148
rect 7564 18096 7616 18148
rect 19892 18096 19944 18148
rect 19156 18028 19208 18080
rect 23756 18173 23765 18207
rect 23765 18173 23799 18207
rect 23799 18173 23808 18207
rect 23756 18164 23808 18173
rect 21456 18096 21508 18148
rect 22008 18096 22060 18148
rect 30196 18164 30248 18216
rect 37924 18164 37976 18216
rect 38200 18071 38252 18080
rect 38200 18037 38209 18071
rect 38209 18037 38243 18071
rect 38243 18037 38252 18071
rect 38200 18028 38252 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 9220 17867 9272 17876
rect 9220 17833 9229 17867
rect 9229 17833 9263 17867
rect 9263 17833 9272 17867
rect 9220 17824 9272 17833
rect 10416 17824 10468 17876
rect 15936 17824 15988 17876
rect 16672 17824 16724 17876
rect 17868 17824 17920 17876
rect 17684 17756 17736 17808
rect 1584 17731 1636 17740
rect 1584 17697 1593 17731
rect 1593 17697 1627 17731
rect 1627 17697 1636 17731
rect 1584 17688 1636 17697
rect 2596 17688 2648 17740
rect 4068 17688 4120 17740
rect 12900 17688 12952 17740
rect 15108 17731 15160 17740
rect 15108 17697 15117 17731
rect 15117 17697 15151 17731
rect 15151 17697 15160 17731
rect 15108 17688 15160 17697
rect 16856 17688 16908 17740
rect 19892 17756 19944 17808
rect 19984 17688 20036 17740
rect 23756 17756 23808 17808
rect 27528 17756 27580 17808
rect 27804 17756 27856 17808
rect 9128 17663 9180 17672
rect 9128 17629 9137 17663
rect 9137 17629 9171 17663
rect 9171 17629 9180 17663
rect 9128 17620 9180 17629
rect 5080 17552 5132 17604
rect 3240 17484 3292 17536
rect 3516 17484 3568 17536
rect 7012 17552 7064 17604
rect 8116 17552 8168 17604
rect 21548 17663 21600 17672
rect 21548 17629 21557 17663
rect 21557 17629 21591 17663
rect 21591 17629 21600 17663
rect 21548 17620 21600 17629
rect 24584 17663 24636 17672
rect 24584 17629 24593 17663
rect 24593 17629 24627 17663
rect 24627 17629 24636 17663
rect 24584 17620 24636 17629
rect 12532 17552 12584 17604
rect 9864 17484 9916 17536
rect 14004 17552 14056 17604
rect 17040 17552 17092 17604
rect 17592 17552 17644 17604
rect 12992 17527 13044 17536
rect 12992 17493 13001 17527
rect 13001 17493 13035 17527
rect 13035 17493 13044 17527
rect 12992 17484 13044 17493
rect 13360 17484 13412 17536
rect 19616 17552 19668 17604
rect 19892 17595 19944 17604
rect 19892 17561 19901 17595
rect 19901 17561 19935 17595
rect 19935 17561 19944 17595
rect 19892 17552 19944 17561
rect 20444 17552 20496 17604
rect 21640 17595 21692 17604
rect 21640 17561 21649 17595
rect 21649 17561 21683 17595
rect 21683 17561 21692 17595
rect 22284 17595 22336 17604
rect 21640 17552 21692 17561
rect 22284 17561 22293 17595
rect 22293 17561 22327 17595
rect 22327 17561 22336 17595
rect 22284 17552 22336 17561
rect 22376 17595 22428 17604
rect 22376 17561 22385 17595
rect 22385 17561 22419 17595
rect 22419 17561 22428 17595
rect 22376 17552 22428 17561
rect 23204 17552 23256 17604
rect 27160 17620 27212 17672
rect 28264 17620 28316 17672
rect 29368 17620 29420 17672
rect 30196 17663 30248 17672
rect 30196 17629 30205 17663
rect 30205 17629 30239 17663
rect 30239 17629 30248 17663
rect 30196 17620 30248 17629
rect 18420 17484 18472 17536
rect 19708 17484 19760 17536
rect 23480 17484 23532 17536
rect 30564 17552 30616 17604
rect 27252 17484 27304 17536
rect 28080 17484 28132 17536
rect 29920 17484 29972 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 8300 17280 8352 17332
rect 3240 17212 3292 17264
rect 10416 17212 10468 17264
rect 1676 17187 1728 17196
rect 1676 17153 1685 17187
rect 1685 17153 1719 17187
rect 1719 17153 1728 17187
rect 1676 17144 1728 17153
rect 2504 17187 2556 17196
rect 2504 17153 2513 17187
rect 2513 17153 2547 17187
rect 2547 17153 2556 17187
rect 2504 17144 2556 17153
rect 7840 17144 7892 17196
rect 11980 17212 12032 17264
rect 10784 17144 10836 17196
rect 14188 17187 14240 17196
rect 14188 17153 14197 17187
rect 14197 17153 14231 17187
rect 14231 17153 14240 17187
rect 17960 17280 18012 17332
rect 20996 17323 21048 17332
rect 20996 17289 21005 17323
rect 21005 17289 21039 17323
rect 21039 17289 21048 17323
rect 20996 17280 21048 17289
rect 28356 17280 28408 17332
rect 17224 17212 17276 17264
rect 22376 17212 22428 17264
rect 14188 17144 14240 17153
rect 17776 17187 17828 17196
rect 17776 17153 17785 17187
rect 17785 17153 17819 17187
rect 17819 17153 17828 17187
rect 17776 17144 17828 17153
rect 17868 17144 17920 17196
rect 9220 17076 9272 17128
rect 25228 17212 25280 17264
rect 27620 17212 27672 17264
rect 27344 17187 27396 17196
rect 1860 17051 1912 17060
rect 1860 17017 1869 17051
rect 1869 17017 1903 17051
rect 1903 17017 1912 17051
rect 1860 17008 1912 17017
rect 1952 17008 2004 17060
rect 8484 17008 8536 17060
rect 8760 17008 8812 17060
rect 11888 17008 11940 17060
rect 11980 17008 12032 17060
rect 17224 17008 17276 17060
rect 27344 17153 27353 17187
rect 27353 17153 27387 17187
rect 27387 17153 27396 17187
rect 27344 17144 27396 17153
rect 28080 17187 28132 17196
rect 28080 17153 28089 17187
rect 28089 17153 28123 17187
rect 28123 17153 28132 17187
rect 28080 17144 28132 17153
rect 26148 17119 26200 17128
rect 26148 17085 26157 17119
rect 26157 17085 26191 17119
rect 26191 17085 26200 17119
rect 26148 17076 26200 17085
rect 29460 17076 29512 17128
rect 3240 16940 3292 16992
rect 8300 16940 8352 16992
rect 9128 16940 9180 16992
rect 15752 16940 15804 16992
rect 16396 16940 16448 16992
rect 26240 17008 26292 17060
rect 29736 17008 29788 17060
rect 17776 16940 17828 16992
rect 17960 16940 18012 16992
rect 20444 16940 20496 16992
rect 24768 16983 24820 16992
rect 24768 16949 24777 16983
rect 24777 16949 24811 16983
rect 24811 16949 24820 16983
rect 24768 16940 24820 16949
rect 26332 16983 26384 16992
rect 26332 16949 26341 16983
rect 26341 16949 26375 16983
rect 26375 16949 26384 16983
rect 26332 16940 26384 16949
rect 26976 16940 27028 16992
rect 28540 16983 28592 16992
rect 28540 16949 28549 16983
rect 28549 16949 28583 16983
rect 28583 16949 28592 16983
rect 28540 16940 28592 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2780 16779 2832 16788
rect 2780 16745 2789 16779
rect 2789 16745 2823 16779
rect 2823 16745 2832 16779
rect 2780 16736 2832 16745
rect 3608 16736 3660 16788
rect 8116 16736 8168 16788
rect 17224 16736 17276 16788
rect 27988 16736 28040 16788
rect 2136 16668 2188 16720
rect 1952 16643 2004 16652
rect 1952 16609 1961 16643
rect 1961 16609 1995 16643
rect 1995 16609 2004 16643
rect 1952 16600 2004 16609
rect 2780 16600 2832 16652
rect 8484 16668 8536 16720
rect 4068 16532 4120 16584
rect 6184 16532 6236 16584
rect 8300 16600 8352 16652
rect 8392 16600 8444 16652
rect 13360 16668 13412 16720
rect 7472 16575 7524 16584
rect 7472 16541 7481 16575
rect 7481 16541 7515 16575
rect 7515 16541 7524 16575
rect 8116 16575 8168 16584
rect 7472 16532 7524 16541
rect 8116 16541 8125 16575
rect 8125 16541 8159 16575
rect 8159 16541 8168 16575
rect 8116 16532 8168 16541
rect 10324 16532 10376 16584
rect 11796 16600 11848 16652
rect 11888 16600 11940 16652
rect 12532 16532 12584 16584
rect 13728 16600 13780 16652
rect 14280 16668 14332 16720
rect 19064 16668 19116 16720
rect 20628 16600 20680 16652
rect 21088 16600 21140 16652
rect 14280 16575 14332 16584
rect 14280 16541 14289 16575
rect 14289 16541 14323 16575
rect 14323 16541 14332 16575
rect 14280 16532 14332 16541
rect 14372 16575 14424 16584
rect 14372 16541 14381 16575
rect 14381 16541 14415 16575
rect 14415 16541 14424 16575
rect 14372 16532 14424 16541
rect 16304 16532 16356 16584
rect 17500 16532 17552 16584
rect 20444 16532 20496 16584
rect 21732 16600 21784 16652
rect 22376 16643 22428 16652
rect 22376 16609 22385 16643
rect 22385 16609 22419 16643
rect 22419 16609 22428 16643
rect 22376 16600 22428 16609
rect 22560 16575 22612 16584
rect 22560 16541 22569 16575
rect 22569 16541 22603 16575
rect 22603 16541 22612 16575
rect 22560 16532 22612 16541
rect 23572 16600 23624 16652
rect 24492 16600 24544 16652
rect 29000 16600 29052 16652
rect 29920 16643 29972 16652
rect 29920 16609 29929 16643
rect 29929 16609 29963 16643
rect 29963 16609 29972 16643
rect 29920 16600 29972 16609
rect 25412 16575 25464 16584
rect 25412 16541 25421 16575
rect 25421 16541 25455 16575
rect 25455 16541 25464 16575
rect 25412 16532 25464 16541
rect 26240 16575 26292 16584
rect 26240 16541 26249 16575
rect 26249 16541 26283 16575
rect 26283 16541 26292 16575
rect 26240 16532 26292 16541
rect 27896 16532 27948 16584
rect 29736 16575 29788 16584
rect 29736 16541 29745 16575
rect 29745 16541 29779 16575
rect 29779 16541 29788 16575
rect 29736 16532 29788 16541
rect 30472 16532 30524 16584
rect 38016 16575 38068 16584
rect 38016 16541 38025 16575
rect 38025 16541 38059 16575
rect 38059 16541 38068 16575
rect 38016 16532 38068 16541
rect 2596 16464 2648 16516
rect 4620 16464 4672 16516
rect 6276 16464 6328 16516
rect 6644 16464 6696 16516
rect 8208 16507 8260 16516
rect 8208 16473 8217 16507
rect 8217 16473 8251 16507
rect 8251 16473 8260 16507
rect 9220 16507 9272 16516
rect 8208 16464 8260 16473
rect 9220 16473 9229 16507
rect 9229 16473 9263 16507
rect 9263 16473 9272 16507
rect 9220 16464 9272 16473
rect 9588 16464 9640 16516
rect 14648 16464 14700 16516
rect 17040 16464 17092 16516
rect 2964 16439 3016 16448
rect 2964 16405 2973 16439
rect 2973 16405 3007 16439
rect 3007 16405 3016 16439
rect 2964 16396 3016 16405
rect 3976 16439 4028 16448
rect 3976 16405 3985 16439
rect 3985 16405 4019 16439
rect 4019 16405 4028 16439
rect 3976 16396 4028 16405
rect 5540 16396 5592 16448
rect 5908 16396 5960 16448
rect 10600 16396 10652 16448
rect 10968 16439 11020 16448
rect 10968 16405 10977 16439
rect 10977 16405 11011 16439
rect 11011 16405 11020 16439
rect 10968 16396 11020 16405
rect 13636 16439 13688 16448
rect 13636 16405 13645 16439
rect 13645 16405 13679 16439
rect 13679 16405 13688 16439
rect 13636 16396 13688 16405
rect 16672 16396 16724 16448
rect 21824 16464 21876 16516
rect 22008 16464 22060 16516
rect 22928 16464 22980 16516
rect 26332 16464 26384 16516
rect 20812 16396 20864 16448
rect 21272 16439 21324 16448
rect 21272 16405 21281 16439
rect 21281 16405 21315 16439
rect 21315 16405 21324 16439
rect 21272 16396 21324 16405
rect 23572 16439 23624 16448
rect 23572 16405 23581 16439
rect 23581 16405 23615 16439
rect 23615 16405 23624 16439
rect 23572 16396 23624 16405
rect 24676 16439 24728 16448
rect 24676 16405 24685 16439
rect 24685 16405 24719 16439
rect 24719 16405 24728 16439
rect 24676 16396 24728 16405
rect 25780 16396 25832 16448
rect 27344 16396 27396 16448
rect 27436 16396 27488 16448
rect 38200 16439 38252 16448
rect 38200 16405 38209 16439
rect 38209 16405 38243 16439
rect 38243 16405 38252 16439
rect 38200 16396 38252 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 3976 16192 4028 16244
rect 5264 16235 5316 16244
rect 5264 16201 5273 16235
rect 5273 16201 5307 16235
rect 5307 16201 5316 16235
rect 5264 16192 5316 16201
rect 7380 16192 7432 16244
rect 7748 16235 7800 16244
rect 7748 16201 7757 16235
rect 7757 16201 7791 16235
rect 7791 16201 7800 16235
rect 7748 16192 7800 16201
rect 7932 16192 7984 16244
rect 9496 16192 9548 16244
rect 10508 16192 10560 16244
rect 10968 16192 11020 16244
rect 12624 16192 12676 16244
rect 16396 16192 16448 16244
rect 2964 16031 3016 16040
rect 2964 15997 2973 16031
rect 2973 15997 3007 16031
rect 3007 15997 3016 16031
rect 2964 15988 3016 15997
rect 3608 16031 3660 16040
rect 3608 15997 3617 16031
rect 3617 15997 3651 16031
rect 3651 15997 3660 16031
rect 3608 15988 3660 15997
rect 5448 16124 5500 16176
rect 6276 16124 6328 16176
rect 5264 16056 5316 16108
rect 5632 16056 5684 16108
rect 6184 16056 6236 16108
rect 9404 16124 9456 16176
rect 7656 16099 7708 16108
rect 4712 15988 4764 16040
rect 5080 15988 5132 16040
rect 7656 16065 7665 16099
rect 7665 16065 7699 16099
rect 7699 16065 7708 16099
rect 7656 16056 7708 16065
rect 8484 16099 8536 16108
rect 8484 16065 8493 16099
rect 8493 16065 8527 16099
rect 8527 16065 8536 16099
rect 8484 16056 8536 16065
rect 6276 15920 6328 15972
rect 7932 15988 7984 16040
rect 9496 16056 9548 16108
rect 11060 16124 11112 16176
rect 11152 16124 11204 16176
rect 16672 16124 16724 16176
rect 10324 16099 10376 16108
rect 10324 16065 10333 16099
rect 10333 16065 10367 16099
rect 10367 16065 10376 16099
rect 10324 16056 10376 16065
rect 10416 16056 10468 16108
rect 10600 15988 10652 16040
rect 20168 16192 20220 16244
rect 22560 16192 22612 16244
rect 26148 16192 26200 16244
rect 17960 16124 18012 16176
rect 20720 16124 20772 16176
rect 23572 16124 23624 16176
rect 27620 16192 27672 16244
rect 29736 16192 29788 16244
rect 27252 16124 27304 16176
rect 19984 16056 20036 16108
rect 21548 16056 21600 16108
rect 25412 16056 25464 16108
rect 25780 16099 25832 16108
rect 25780 16065 25789 16099
rect 25789 16065 25823 16099
rect 25823 16065 25832 16099
rect 25780 16056 25832 16065
rect 29000 16099 29052 16108
rect 29000 16065 29009 16099
rect 29009 16065 29043 16099
rect 29043 16065 29052 16099
rect 29000 16056 29052 16065
rect 18420 15988 18472 16040
rect 20996 15988 21048 16040
rect 26332 15988 26384 16040
rect 27896 16031 27948 16040
rect 27896 15997 27905 16031
rect 27905 15997 27939 16031
rect 27939 15997 27948 16031
rect 27896 15988 27948 15997
rect 36912 16056 36964 16108
rect 37740 15988 37792 16040
rect 1768 15895 1820 15904
rect 1768 15861 1777 15895
rect 1777 15861 1811 15895
rect 1811 15861 1820 15895
rect 1768 15852 1820 15861
rect 6644 15895 6696 15904
rect 6644 15861 6653 15895
rect 6653 15861 6687 15895
rect 6687 15861 6696 15895
rect 6644 15852 6696 15861
rect 9496 15920 9548 15972
rect 22836 15920 22888 15972
rect 24676 15920 24728 15972
rect 28172 15920 28224 15972
rect 10232 15852 10284 15904
rect 20352 15852 20404 15904
rect 20720 15895 20772 15904
rect 20720 15861 20729 15895
rect 20729 15861 20763 15895
rect 20763 15861 20772 15895
rect 20720 15852 20772 15861
rect 38016 15852 38068 15904
rect 38200 15895 38252 15904
rect 38200 15861 38209 15895
rect 38209 15861 38243 15895
rect 38243 15861 38252 15895
rect 38200 15852 38252 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 1860 15648 1912 15700
rect 3332 15691 3384 15700
rect 2780 15580 2832 15632
rect 3332 15657 3341 15691
rect 3341 15657 3375 15691
rect 3375 15657 3384 15691
rect 3332 15648 3384 15657
rect 4068 15691 4120 15700
rect 4068 15657 4077 15691
rect 4077 15657 4111 15691
rect 4111 15657 4120 15691
rect 4068 15648 4120 15657
rect 5816 15648 5868 15700
rect 6736 15691 6788 15700
rect 6736 15657 6745 15691
rect 6745 15657 6779 15691
rect 6779 15657 6788 15691
rect 6736 15648 6788 15657
rect 8668 15648 8720 15700
rect 9036 15648 9088 15700
rect 10600 15691 10652 15700
rect 10600 15657 10609 15691
rect 10609 15657 10643 15691
rect 10643 15657 10652 15691
rect 10600 15648 10652 15657
rect 12440 15648 12492 15700
rect 14556 15691 14608 15700
rect 5264 15580 5316 15632
rect 6920 15580 6972 15632
rect 8300 15580 8352 15632
rect 8760 15580 8812 15632
rect 9312 15580 9364 15632
rect 10232 15580 10284 15632
rect 14556 15657 14565 15691
rect 14565 15657 14599 15691
rect 14599 15657 14608 15691
rect 14556 15648 14608 15657
rect 15476 15691 15528 15700
rect 15476 15657 15485 15691
rect 15485 15657 15519 15691
rect 15519 15657 15528 15691
rect 15476 15648 15528 15657
rect 15844 15648 15896 15700
rect 16304 15648 16356 15700
rect 16764 15691 16816 15700
rect 16764 15657 16773 15691
rect 16773 15657 16807 15691
rect 16807 15657 16816 15691
rect 16764 15648 16816 15657
rect 17960 15648 18012 15700
rect 18144 15648 18196 15700
rect 22008 15648 22060 15700
rect 23848 15648 23900 15700
rect 18788 15580 18840 15632
rect 2320 15512 2372 15564
rect 8852 15512 8904 15564
rect 3976 15487 4028 15496
rect 3976 15453 3985 15487
rect 3985 15453 4019 15487
rect 4019 15453 4028 15487
rect 3976 15444 4028 15453
rect 5632 15444 5684 15496
rect 5908 15444 5960 15496
rect 6184 15444 6236 15496
rect 6828 15444 6880 15496
rect 6920 15444 6972 15496
rect 8300 15444 8352 15496
rect 9404 15512 9456 15564
rect 9588 15512 9640 15564
rect 12808 15512 12860 15564
rect 9128 15487 9180 15496
rect 1860 15308 1912 15360
rect 7656 15376 7708 15428
rect 9128 15453 9137 15487
rect 9137 15453 9171 15487
rect 9171 15453 9180 15487
rect 9128 15444 9180 15453
rect 10416 15444 10468 15496
rect 11612 15444 11664 15496
rect 15476 15444 15528 15496
rect 17040 15444 17092 15496
rect 17868 15444 17920 15496
rect 18052 15444 18104 15496
rect 5448 15308 5500 15360
rect 6000 15308 6052 15360
rect 11980 15308 12032 15360
rect 13636 15376 13688 15428
rect 15844 15376 15896 15428
rect 16304 15376 16356 15428
rect 19892 15444 19944 15496
rect 19984 15376 20036 15428
rect 24676 15512 24728 15564
rect 26884 15512 26936 15564
rect 22928 15444 22980 15496
rect 23388 15444 23440 15496
rect 21180 15419 21232 15428
rect 21180 15385 21189 15419
rect 21189 15385 21223 15419
rect 21223 15385 21232 15419
rect 21180 15376 21232 15385
rect 13084 15308 13136 15360
rect 15936 15308 15988 15360
rect 18144 15308 18196 15360
rect 26516 15376 26568 15428
rect 27436 15419 27488 15428
rect 27436 15385 27445 15419
rect 27445 15385 27479 15419
rect 27479 15385 27488 15419
rect 27436 15376 27488 15385
rect 37280 15308 37332 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 4620 15104 4672 15156
rect 4896 15104 4948 15156
rect 7196 15104 7248 15156
rect 6644 15036 6696 15088
rect 6828 15036 6880 15088
rect 14740 15104 14792 15156
rect 15384 15104 15436 15156
rect 16120 15104 16172 15156
rect 16488 15104 16540 15156
rect 18696 15104 18748 15156
rect 19340 15104 19392 15156
rect 4068 15011 4120 15020
rect 4068 14977 4077 15011
rect 4077 14977 4111 15011
rect 4111 14977 4120 15011
rect 4068 14968 4120 14977
rect 2964 14943 3016 14952
rect 2504 14832 2556 14884
rect 2964 14909 2973 14943
rect 2973 14909 3007 14943
rect 3007 14909 3016 14943
rect 2964 14900 3016 14909
rect 3148 14943 3200 14952
rect 3148 14909 3157 14943
rect 3157 14909 3191 14943
rect 3191 14909 3200 14943
rect 3148 14900 3200 14909
rect 5172 14968 5224 15020
rect 5448 14968 5500 15020
rect 8024 15036 8076 15088
rect 9680 15036 9732 15088
rect 20720 15104 20772 15156
rect 24860 15147 24912 15156
rect 20904 15079 20956 15088
rect 20904 15045 20913 15079
rect 20913 15045 20947 15079
rect 20947 15045 20956 15079
rect 20904 15036 20956 15045
rect 8392 14968 8444 15020
rect 8760 15011 8812 15020
rect 8760 14977 8769 15011
rect 8769 14977 8803 15011
rect 8803 14977 8812 15011
rect 8760 14968 8812 14977
rect 9772 15011 9824 15020
rect 9772 14977 9781 15011
rect 9781 14977 9815 15011
rect 9815 14977 9824 15011
rect 9772 14968 9824 14977
rect 5908 14900 5960 14952
rect 6276 14900 6328 14952
rect 6736 14900 6788 14952
rect 11704 14900 11756 14952
rect 11888 14943 11940 14952
rect 11888 14909 11897 14943
rect 11897 14909 11931 14943
rect 11931 14909 11940 14943
rect 11888 14900 11940 14909
rect 12072 14900 12124 14952
rect 12900 14943 12952 14952
rect 12900 14909 12909 14943
rect 12909 14909 12943 14943
rect 12943 14909 12952 14943
rect 16028 14968 16080 15020
rect 17040 15011 17092 15020
rect 17040 14977 17049 15011
rect 17049 14977 17083 15011
rect 17083 14977 17092 15011
rect 17040 14968 17092 14977
rect 18788 15011 18840 15020
rect 18788 14977 18797 15011
rect 18797 14977 18831 15011
rect 18831 14977 18840 15011
rect 18788 14968 18840 14977
rect 24860 15113 24869 15147
rect 24869 15113 24903 15147
rect 24903 15113 24912 15147
rect 24860 15104 24912 15113
rect 24952 15104 25004 15156
rect 26056 15104 26108 15156
rect 26516 15147 26568 15156
rect 26516 15113 26525 15147
rect 26525 15113 26559 15147
rect 26559 15113 26568 15147
rect 26516 15104 26568 15113
rect 27712 15147 27764 15156
rect 27712 15113 27721 15147
rect 27721 15113 27755 15147
rect 27755 15113 27764 15147
rect 27712 15104 27764 15113
rect 36912 15104 36964 15156
rect 23480 15079 23532 15088
rect 23480 15045 23489 15079
rect 23489 15045 23523 15079
rect 23523 15045 23532 15079
rect 23480 15036 23532 15045
rect 27896 15036 27948 15088
rect 12900 14900 12952 14909
rect 13636 14900 13688 14952
rect 14648 14943 14700 14952
rect 14648 14909 14657 14943
rect 14657 14909 14691 14943
rect 14691 14909 14700 14943
rect 14648 14900 14700 14909
rect 16120 14900 16172 14952
rect 19064 14900 19116 14952
rect 9404 14832 9456 14884
rect 3608 14807 3660 14816
rect 3608 14773 3617 14807
rect 3617 14773 3651 14807
rect 3651 14773 3660 14807
rect 3608 14764 3660 14773
rect 9956 14832 10008 14884
rect 10232 14832 10284 14884
rect 15844 14832 15896 14884
rect 27436 15011 27488 15020
rect 19340 14900 19392 14952
rect 10048 14764 10100 14816
rect 11520 14764 11572 14816
rect 16028 14764 16080 14816
rect 18696 14764 18748 14816
rect 19616 14832 19668 14884
rect 21088 14900 21140 14952
rect 22744 14764 22796 14816
rect 22928 14900 22980 14952
rect 25320 14900 25372 14952
rect 27436 14977 27445 15011
rect 27445 14977 27479 15011
rect 27479 14977 27488 15011
rect 27436 14968 27488 14977
rect 29368 15011 29420 15020
rect 29368 14977 29377 15011
rect 29377 14977 29411 15011
rect 29411 14977 29420 15011
rect 29368 14968 29420 14977
rect 27528 14900 27580 14952
rect 34520 14968 34572 15020
rect 37740 14968 37792 15020
rect 37096 14900 37148 14952
rect 35440 14832 35492 14884
rect 23572 14764 23624 14816
rect 29000 14764 29052 14816
rect 37924 14764 37976 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 3608 14560 3660 14612
rect 11888 14560 11940 14612
rect 12072 14560 12124 14612
rect 5724 14492 5776 14544
rect 12440 14492 12492 14544
rect 14372 14492 14424 14544
rect 2504 14467 2556 14476
rect 2504 14433 2513 14467
rect 2513 14433 2547 14467
rect 2547 14433 2556 14467
rect 2504 14424 2556 14433
rect 7012 14424 7064 14476
rect 8576 14424 8628 14476
rect 2872 14356 2924 14408
rect 2136 14331 2188 14340
rect 2136 14297 2145 14331
rect 2145 14297 2179 14331
rect 2179 14297 2188 14331
rect 2136 14288 2188 14297
rect 2228 14331 2280 14340
rect 2228 14297 2237 14331
rect 2237 14297 2271 14331
rect 2271 14297 2280 14331
rect 2228 14288 2280 14297
rect 4068 14288 4120 14340
rect 5632 14356 5684 14408
rect 7564 14356 7616 14408
rect 5908 14288 5960 14340
rect 6184 14331 6236 14340
rect 6184 14297 6193 14331
rect 6193 14297 6227 14331
rect 6227 14297 6236 14331
rect 10232 14424 10284 14476
rect 11152 14424 11204 14476
rect 12072 14424 12124 14476
rect 20168 14560 20220 14612
rect 21180 14560 21232 14612
rect 21364 14560 21416 14612
rect 21916 14560 21968 14612
rect 26056 14560 26108 14612
rect 15844 14492 15896 14544
rect 8944 14356 8996 14408
rect 15016 14424 15068 14476
rect 6184 14288 6236 14297
rect 5172 14220 5224 14272
rect 5448 14220 5500 14272
rect 10048 14331 10100 14340
rect 10048 14297 10057 14331
rect 10057 14297 10091 14331
rect 10091 14297 10100 14331
rect 10048 14288 10100 14297
rect 11060 14288 11112 14340
rect 11980 14331 12032 14340
rect 11980 14297 11989 14331
rect 11989 14297 12023 14331
rect 12023 14297 12032 14331
rect 13084 14356 13136 14408
rect 12900 14331 12952 14340
rect 11980 14288 12032 14297
rect 7656 14220 7708 14272
rect 7840 14220 7892 14272
rect 12900 14297 12909 14331
rect 12909 14297 12943 14331
rect 12943 14297 12952 14331
rect 12900 14288 12952 14297
rect 12440 14220 12492 14272
rect 15200 14331 15252 14340
rect 15200 14297 15209 14331
rect 15209 14297 15243 14331
rect 15243 14297 15252 14331
rect 15200 14288 15252 14297
rect 13268 14220 13320 14272
rect 14372 14220 14424 14272
rect 16028 14424 16080 14476
rect 16304 14467 16356 14476
rect 16304 14433 16313 14467
rect 16313 14433 16347 14467
rect 16347 14433 16356 14467
rect 16304 14424 16356 14433
rect 16672 14424 16724 14476
rect 19248 14424 19300 14476
rect 21088 14424 21140 14476
rect 20168 14399 20220 14408
rect 20168 14365 20177 14399
rect 20177 14365 20211 14399
rect 20211 14365 20220 14399
rect 20168 14356 20220 14365
rect 16396 14288 16448 14340
rect 19616 14331 19668 14340
rect 19616 14297 19625 14331
rect 19625 14297 19659 14331
rect 19659 14297 19668 14331
rect 23572 14424 23624 14476
rect 26148 14492 26200 14544
rect 29184 14424 29236 14476
rect 29000 14399 29052 14408
rect 29000 14365 29009 14399
rect 29009 14365 29043 14399
rect 29043 14365 29052 14399
rect 29000 14356 29052 14365
rect 31944 14399 31996 14408
rect 31944 14365 31953 14399
rect 31953 14365 31987 14399
rect 31987 14365 31996 14399
rect 31944 14356 31996 14365
rect 19616 14288 19668 14297
rect 22928 14288 22980 14340
rect 23664 14288 23716 14340
rect 21272 14220 21324 14272
rect 23296 14220 23348 14272
rect 25596 14288 25648 14340
rect 30288 14331 30340 14340
rect 30288 14297 30297 14331
rect 30297 14297 30331 14331
rect 30331 14297 30340 14331
rect 30288 14288 30340 14297
rect 30380 14331 30432 14340
rect 30380 14297 30389 14331
rect 30389 14297 30423 14331
rect 30423 14297 30432 14331
rect 30380 14288 30432 14297
rect 28448 14220 28500 14272
rect 38200 14263 38252 14272
rect 38200 14229 38209 14263
rect 38209 14229 38243 14263
rect 38243 14229 38252 14263
rect 38200 14220 38252 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 2136 14016 2188 14068
rect 3424 14016 3476 14068
rect 4988 14016 5040 14068
rect 9496 14016 9548 14068
rect 3700 13991 3752 14000
rect 3700 13957 3709 13991
rect 3709 13957 3743 13991
rect 3743 13957 3752 13991
rect 3700 13948 3752 13957
rect 5448 13948 5500 14000
rect 7656 13991 7708 14000
rect 7656 13957 7665 13991
rect 7665 13957 7699 13991
rect 7699 13957 7708 13991
rect 7656 13948 7708 13957
rect 9220 13991 9272 14000
rect 9220 13957 9229 13991
rect 9229 13957 9263 13991
rect 9263 13957 9272 13991
rect 9220 13948 9272 13957
rect 9404 13948 9456 14000
rect 9772 13948 9824 14000
rect 10600 13991 10652 14000
rect 10600 13957 10609 13991
rect 10609 13957 10643 13991
rect 10643 13957 10652 13991
rect 10600 13948 10652 13957
rect 11888 13991 11940 14000
rect 11888 13957 11897 13991
rect 11897 13957 11931 13991
rect 11931 13957 11940 13991
rect 11888 13948 11940 13957
rect 1400 13880 1452 13932
rect 2872 13923 2924 13932
rect 2872 13889 2881 13923
rect 2881 13889 2915 13923
rect 2915 13889 2924 13923
rect 2872 13880 2924 13889
rect 2964 13812 3016 13864
rect 3332 13812 3384 13864
rect 6368 13880 6420 13932
rect 3424 13744 3476 13796
rect 6736 13812 6788 13864
rect 7840 13812 7892 13864
rect 9128 13855 9180 13864
rect 9128 13821 9137 13855
rect 9137 13821 9171 13855
rect 9171 13821 9180 13855
rect 9128 13812 9180 13821
rect 9404 13855 9456 13864
rect 9404 13821 9413 13855
rect 9413 13821 9447 13855
rect 9447 13821 9456 13855
rect 9404 13812 9456 13821
rect 10508 13855 10560 13864
rect 10508 13821 10517 13855
rect 10517 13821 10551 13855
rect 10551 13821 10560 13855
rect 10508 13812 10560 13821
rect 11244 13812 11296 13864
rect 11520 13812 11572 13864
rect 12072 13855 12124 13864
rect 12072 13821 12081 13855
rect 12081 13821 12115 13855
rect 12115 13821 12124 13855
rect 12072 13812 12124 13821
rect 16304 14016 16356 14068
rect 20996 14059 21048 14068
rect 14096 13948 14148 14000
rect 15752 13948 15804 14000
rect 19064 13948 19116 14000
rect 16672 13880 16724 13932
rect 17316 13880 17368 13932
rect 17500 13923 17552 13932
rect 17500 13889 17509 13923
rect 17509 13889 17543 13923
rect 17543 13889 17552 13923
rect 17500 13880 17552 13889
rect 19892 13991 19944 14000
rect 19892 13957 19901 13991
rect 19901 13957 19935 13991
rect 19935 13957 19944 13991
rect 19892 13948 19944 13957
rect 20996 14025 21005 14059
rect 21005 14025 21039 14059
rect 21039 14025 21048 14059
rect 20996 14016 21048 14025
rect 21088 14016 21140 14068
rect 30288 14016 30340 14068
rect 25964 13991 26016 14000
rect 25964 13957 25973 13991
rect 25973 13957 26007 13991
rect 26007 13957 26016 13991
rect 25964 13948 26016 13957
rect 26056 13948 26108 14000
rect 30472 13948 30524 14000
rect 21548 13880 21600 13932
rect 21824 13880 21876 13932
rect 22008 13923 22060 13932
rect 22008 13889 22017 13923
rect 22017 13889 22051 13923
rect 22051 13889 22060 13923
rect 22008 13880 22060 13889
rect 25228 13880 25280 13932
rect 28448 13923 28500 13932
rect 28448 13889 28457 13923
rect 28457 13889 28491 13923
rect 28491 13889 28500 13923
rect 28448 13880 28500 13889
rect 36912 13880 36964 13932
rect 13636 13812 13688 13864
rect 13912 13812 13964 13864
rect 14096 13812 14148 13864
rect 17132 13812 17184 13864
rect 19340 13812 19392 13864
rect 3976 13676 4028 13728
rect 17500 13744 17552 13796
rect 22192 13812 22244 13864
rect 26516 13812 26568 13864
rect 27528 13812 27580 13864
rect 19892 13744 19944 13796
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 2596 13515 2648 13524
rect 2596 13481 2605 13515
rect 2605 13481 2639 13515
rect 2639 13481 2648 13515
rect 2596 13472 2648 13481
rect 3332 13515 3384 13524
rect 3332 13481 3341 13515
rect 3341 13481 3375 13515
rect 3375 13481 3384 13515
rect 3332 13472 3384 13481
rect 3700 13472 3752 13524
rect 4712 13515 4764 13524
rect 4712 13481 4721 13515
rect 4721 13481 4755 13515
rect 4755 13481 4764 13515
rect 4712 13472 4764 13481
rect 6184 13472 6236 13524
rect 9220 13472 9272 13524
rect 11888 13472 11940 13524
rect 8300 13404 8352 13456
rect 9128 13404 9180 13456
rect 12348 13404 12400 13456
rect 16396 13404 16448 13456
rect 16672 13472 16724 13524
rect 21456 13472 21508 13524
rect 22376 13472 22428 13524
rect 25964 13515 26016 13524
rect 25964 13481 25973 13515
rect 25973 13481 26007 13515
rect 26007 13481 26016 13515
rect 25964 13472 26016 13481
rect 31944 13404 31996 13456
rect 1676 13311 1728 13320
rect 1676 13277 1685 13311
rect 1685 13277 1719 13311
rect 1719 13277 1728 13311
rect 1676 13268 1728 13277
rect 2964 13268 3016 13320
rect 3240 13311 3292 13320
rect 3240 13277 3249 13311
rect 3249 13277 3283 13311
rect 3283 13277 3292 13311
rect 3240 13268 3292 13277
rect 4160 13268 4212 13320
rect 5356 13268 5408 13320
rect 5448 13268 5500 13320
rect 8116 13311 8168 13320
rect 8116 13277 8125 13311
rect 8125 13277 8159 13311
rect 8159 13277 8168 13311
rect 8116 13268 8168 13277
rect 9496 13311 9548 13320
rect 9496 13277 9505 13311
rect 9505 13277 9539 13311
rect 9539 13277 9548 13311
rect 9496 13268 9548 13277
rect 10140 13268 10192 13320
rect 5080 13200 5132 13252
rect 4160 13132 4212 13184
rect 5540 13200 5592 13252
rect 12716 13268 12768 13320
rect 14280 13268 14332 13320
rect 9312 13175 9364 13184
rect 9312 13141 9321 13175
rect 9321 13141 9355 13175
rect 9355 13141 9364 13175
rect 9312 13132 9364 13141
rect 13728 13132 13780 13184
rect 15568 13200 15620 13252
rect 15752 13243 15804 13252
rect 15752 13209 15761 13243
rect 15761 13209 15795 13243
rect 15795 13209 15804 13243
rect 15752 13200 15804 13209
rect 16304 13243 16356 13252
rect 16304 13209 16313 13243
rect 16313 13209 16347 13243
rect 16347 13209 16356 13243
rect 16304 13200 16356 13209
rect 17224 13200 17276 13252
rect 17684 13268 17736 13320
rect 23296 13336 23348 13388
rect 21916 13268 21968 13320
rect 23388 13311 23440 13320
rect 17500 13200 17552 13252
rect 16672 13132 16724 13184
rect 16856 13132 16908 13184
rect 22652 13200 22704 13252
rect 23388 13277 23397 13311
rect 23397 13277 23431 13311
rect 23431 13277 23440 13311
rect 23388 13268 23440 13277
rect 25688 13268 25740 13320
rect 25964 13268 26016 13320
rect 27896 13268 27948 13320
rect 32312 13268 32364 13320
rect 23940 13200 23992 13252
rect 25228 13243 25280 13252
rect 25228 13209 25237 13243
rect 25237 13209 25271 13243
rect 25271 13209 25280 13243
rect 25228 13200 25280 13209
rect 37740 13200 37792 13252
rect 23756 13132 23808 13184
rect 25320 13175 25372 13184
rect 25320 13141 25329 13175
rect 25329 13141 25363 13175
rect 25363 13141 25372 13175
rect 25320 13132 25372 13141
rect 26056 13132 26108 13184
rect 32496 13132 32548 13184
rect 38200 13175 38252 13184
rect 38200 13141 38209 13175
rect 38209 13141 38243 13175
rect 38243 13141 38252 13175
rect 38200 13132 38252 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 3056 12928 3108 12980
rect 3792 12928 3844 12980
rect 4620 12928 4672 12980
rect 2136 12860 2188 12912
rect 7196 12903 7248 12912
rect 7196 12869 7205 12903
rect 7205 12869 7239 12903
rect 7239 12869 7248 12903
rect 7196 12860 7248 12869
rect 2872 12792 2924 12844
rect 3424 12835 3476 12844
rect 3424 12801 3433 12835
rect 3433 12801 3467 12835
rect 3467 12801 3476 12835
rect 3424 12792 3476 12801
rect 3884 12792 3936 12844
rect 4988 12835 5040 12844
rect 4988 12801 4997 12835
rect 4997 12801 5031 12835
rect 5031 12801 5040 12835
rect 4988 12792 5040 12801
rect 1676 12767 1728 12776
rect 1676 12733 1685 12767
rect 1685 12733 1719 12767
rect 1719 12733 1728 12767
rect 1676 12724 1728 12733
rect 8300 12724 8352 12776
rect 2320 12656 2372 12708
rect 11060 12860 11112 12912
rect 14648 12928 14700 12980
rect 15568 12971 15620 12980
rect 15568 12937 15577 12971
rect 15577 12937 15611 12971
rect 15611 12937 15620 12971
rect 15568 12928 15620 12937
rect 16856 12971 16908 12980
rect 16856 12937 16865 12971
rect 16865 12937 16899 12971
rect 16899 12937 16908 12971
rect 16856 12928 16908 12937
rect 17224 12928 17276 12980
rect 18972 12928 19024 12980
rect 25320 12928 25372 12980
rect 29184 12971 29236 12980
rect 29184 12937 29193 12971
rect 29193 12937 29227 12971
rect 29227 12937 29236 12971
rect 29184 12928 29236 12937
rect 32312 12971 32364 12980
rect 32312 12937 32321 12971
rect 32321 12937 32355 12971
rect 32355 12937 32364 12971
rect 32312 12928 32364 12937
rect 15384 12792 15436 12844
rect 17040 12835 17092 12844
rect 13820 12724 13872 12776
rect 17040 12801 17049 12835
rect 17049 12801 17083 12835
rect 17083 12801 17092 12835
rect 17040 12792 17092 12801
rect 17868 12860 17920 12912
rect 17500 12792 17552 12844
rect 22836 12860 22888 12912
rect 23756 12903 23808 12912
rect 23756 12869 23765 12903
rect 23765 12869 23799 12903
rect 23799 12869 23808 12903
rect 23756 12860 23808 12869
rect 17868 12724 17920 12776
rect 22468 12792 22520 12844
rect 32496 12835 32548 12844
rect 16396 12656 16448 12708
rect 23480 12724 23532 12776
rect 15200 12588 15252 12640
rect 21640 12656 21692 12708
rect 23572 12656 23624 12708
rect 32496 12801 32505 12835
rect 32505 12801 32539 12835
rect 32539 12801 32548 12835
rect 32496 12792 32548 12801
rect 38292 12835 38344 12844
rect 38292 12801 38301 12835
rect 38301 12801 38335 12835
rect 38335 12801 38344 12835
rect 38292 12792 38344 12801
rect 20076 12588 20128 12640
rect 20812 12588 20864 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 2412 12427 2464 12436
rect 2412 12393 2421 12427
rect 2421 12393 2455 12427
rect 2455 12393 2464 12427
rect 2412 12384 2464 12393
rect 2780 12384 2832 12436
rect 7196 12384 7248 12436
rect 8576 12384 8628 12436
rect 1768 12359 1820 12368
rect 1768 12325 1777 12359
rect 1777 12325 1811 12359
rect 1811 12325 1820 12359
rect 1768 12316 1820 12325
rect 10600 12316 10652 12368
rect 2412 12248 2464 12300
rect 3424 12248 3476 12300
rect 11520 12248 11572 12300
rect 2964 12223 3016 12232
rect 2964 12189 2973 12223
rect 2973 12189 3007 12223
rect 3007 12189 3016 12223
rect 2964 12180 3016 12189
rect 5540 12223 5592 12232
rect 5540 12189 5549 12223
rect 5549 12189 5583 12223
rect 5583 12189 5592 12223
rect 5540 12180 5592 12189
rect 6460 12180 6512 12232
rect 13452 12316 13504 12368
rect 15384 12384 15436 12436
rect 18604 12384 18656 12436
rect 23756 12384 23808 12436
rect 18420 12316 18472 12368
rect 19248 12316 19300 12368
rect 13820 12248 13872 12300
rect 14372 12291 14424 12300
rect 14372 12257 14381 12291
rect 14381 12257 14415 12291
rect 14415 12257 14424 12291
rect 14372 12248 14424 12257
rect 16304 12248 16356 12300
rect 20536 12248 20588 12300
rect 24860 12316 24912 12368
rect 22652 12291 22704 12300
rect 22652 12257 22661 12291
rect 22661 12257 22695 12291
rect 22695 12257 22704 12291
rect 22652 12248 22704 12257
rect 23572 12248 23624 12300
rect 30840 12248 30892 12300
rect 11704 12180 11756 12232
rect 16120 12223 16172 12232
rect 3792 12112 3844 12164
rect 4620 12112 4672 12164
rect 10324 12112 10376 12164
rect 7932 12044 7984 12096
rect 11336 12044 11388 12096
rect 16120 12189 16129 12223
rect 16129 12189 16163 12223
rect 16163 12189 16172 12223
rect 16120 12180 16172 12189
rect 23756 12223 23808 12232
rect 23756 12189 23765 12223
rect 23765 12189 23799 12223
rect 23799 12189 23808 12223
rect 23756 12180 23808 12189
rect 14740 12112 14792 12164
rect 20076 12155 20128 12164
rect 20076 12121 20085 12155
rect 20085 12121 20119 12155
rect 20119 12121 20128 12155
rect 20076 12112 20128 12121
rect 17316 12044 17368 12096
rect 24308 12112 24360 12164
rect 24768 12155 24820 12164
rect 24768 12121 24777 12155
rect 24777 12121 24811 12155
rect 24811 12121 24820 12155
rect 26516 12155 26568 12164
rect 24768 12112 24820 12121
rect 26516 12121 26525 12155
rect 26525 12121 26559 12155
rect 26559 12121 26568 12155
rect 26516 12112 26568 12121
rect 26976 12112 27028 12164
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 2964 11840 3016 11892
rect 5632 11883 5684 11892
rect 5632 11849 5641 11883
rect 5641 11849 5675 11883
rect 5675 11849 5684 11883
rect 5632 11840 5684 11849
rect 7932 11883 7984 11892
rect 7932 11849 7941 11883
rect 7941 11849 7975 11883
rect 7975 11849 7984 11883
rect 7932 11840 7984 11849
rect 2320 11772 2372 11824
rect 2872 11772 2924 11824
rect 6736 11815 6788 11824
rect 6736 11781 6745 11815
rect 6745 11781 6779 11815
rect 6779 11781 6788 11815
rect 6736 11772 6788 11781
rect 7840 11772 7892 11824
rect 2412 11704 2464 11756
rect 3608 11704 3660 11756
rect 6460 11704 6512 11756
rect 2504 11568 2556 11620
rect 6828 11636 6880 11688
rect 9772 11772 9824 11824
rect 11980 11772 12032 11824
rect 14372 11840 14424 11892
rect 14740 11883 14792 11892
rect 14740 11849 14749 11883
rect 14749 11849 14783 11883
rect 14783 11849 14792 11883
rect 14740 11840 14792 11849
rect 17040 11840 17092 11892
rect 19340 11840 19392 11892
rect 19524 11840 19576 11892
rect 23296 11840 23348 11892
rect 21916 11772 21968 11824
rect 13728 11704 13780 11756
rect 10508 11636 10560 11688
rect 10692 11679 10744 11688
rect 10692 11645 10701 11679
rect 10701 11645 10735 11679
rect 10735 11645 10744 11679
rect 10692 11636 10744 11645
rect 14188 11704 14240 11756
rect 14556 11704 14608 11756
rect 17224 11704 17276 11756
rect 20720 11704 20772 11756
rect 34520 11704 34572 11756
rect 7932 11568 7984 11620
rect 5724 11500 5776 11552
rect 9772 11500 9824 11552
rect 10416 11500 10468 11552
rect 15660 11636 15712 11688
rect 25780 11636 25832 11688
rect 28172 11679 28224 11688
rect 28172 11645 28181 11679
rect 28181 11645 28215 11679
rect 28215 11645 28224 11679
rect 28172 11636 28224 11645
rect 28356 11679 28408 11688
rect 28356 11645 28365 11679
rect 28365 11645 28399 11679
rect 28399 11645 28408 11679
rect 28356 11636 28408 11645
rect 11152 11568 11204 11620
rect 11612 11568 11664 11620
rect 10876 11500 10928 11552
rect 16028 11568 16080 11620
rect 28540 11611 28592 11620
rect 28540 11577 28549 11611
rect 28549 11577 28583 11611
rect 28583 11577 28592 11611
rect 28540 11568 28592 11577
rect 14188 11500 14240 11552
rect 18236 11500 18288 11552
rect 22192 11500 22244 11552
rect 24216 11500 24268 11552
rect 27344 11500 27396 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1860 11296 1912 11348
rect 3976 11160 4028 11212
rect 6828 11296 6880 11348
rect 10508 11296 10560 11348
rect 11980 11296 12032 11348
rect 14188 11296 14240 11348
rect 17040 11296 17092 11348
rect 22100 11296 22152 11348
rect 26516 11296 26568 11348
rect 27344 11296 27396 11348
rect 37096 11296 37148 11348
rect 5172 11203 5224 11212
rect 5172 11169 5181 11203
rect 5181 11169 5215 11203
rect 5215 11169 5224 11203
rect 5172 11160 5224 11169
rect 8208 11160 8260 11212
rect 10692 11203 10744 11212
rect 1308 11092 1360 11144
rect 6092 11092 6144 11144
rect 7104 11092 7156 11144
rect 8576 11135 8628 11144
rect 8576 11101 8585 11135
rect 8585 11101 8619 11135
rect 8619 11101 8628 11135
rect 10692 11169 10701 11203
rect 10701 11169 10735 11203
rect 10735 11169 10744 11203
rect 10692 11160 10744 11169
rect 11152 11203 11204 11212
rect 11152 11169 11161 11203
rect 11161 11169 11195 11203
rect 11195 11169 11204 11203
rect 11152 11160 11204 11169
rect 8576 11092 8628 11101
rect 9864 11092 9916 11144
rect 10508 11092 10560 11144
rect 2320 11067 2372 11076
rect 2320 11033 2329 11067
rect 2329 11033 2363 11067
rect 2363 11033 2372 11067
rect 2320 11024 2372 11033
rect 2412 11067 2464 11076
rect 2412 11033 2421 11067
rect 2421 11033 2455 11067
rect 2455 11033 2464 11067
rect 2412 11024 2464 11033
rect 4896 11067 4948 11076
rect 4896 11033 4905 11067
rect 4905 11033 4939 11067
rect 4939 11033 4948 11067
rect 4896 11024 4948 11033
rect 7932 11067 7984 11076
rect 7932 11033 7941 11067
rect 7941 11033 7975 11067
rect 7975 11033 7984 11067
rect 7932 11024 7984 11033
rect 11612 11160 11664 11212
rect 14648 11228 14700 11280
rect 37832 11228 37884 11280
rect 17684 11160 17736 11212
rect 22192 11203 22244 11212
rect 22192 11169 22201 11203
rect 22201 11169 22235 11203
rect 22235 11169 22244 11203
rect 22192 11160 22244 11169
rect 25780 11203 25832 11212
rect 12992 11092 13044 11144
rect 15660 11092 15712 11144
rect 17040 11024 17092 11076
rect 17316 11067 17368 11076
rect 17316 11033 17325 11067
rect 17325 11033 17359 11067
rect 17359 11033 17368 11067
rect 18236 11067 18288 11076
rect 17316 11024 17368 11033
rect 18236 11033 18245 11067
rect 18245 11033 18279 11067
rect 18279 11033 18288 11067
rect 20536 11067 20588 11076
rect 18236 11024 18288 11033
rect 20536 11033 20545 11067
rect 20545 11033 20579 11067
rect 20579 11033 20588 11067
rect 20536 11024 20588 11033
rect 20812 11024 20864 11076
rect 23204 11092 23256 11144
rect 22100 11024 22152 11076
rect 23112 11024 23164 11076
rect 24768 11067 24820 11076
rect 24768 11033 24777 11067
rect 24777 11033 24811 11067
rect 24811 11033 24820 11067
rect 24768 11024 24820 11033
rect 25320 11067 25372 11076
rect 25320 11033 25329 11067
rect 25329 11033 25363 11067
rect 25363 11033 25372 11067
rect 25320 11024 25372 11033
rect 25780 11169 25789 11203
rect 25789 11169 25823 11203
rect 25823 11169 25832 11203
rect 25780 11160 25832 11169
rect 28172 11203 28224 11212
rect 28172 11169 28181 11203
rect 28181 11169 28215 11203
rect 28215 11169 28224 11203
rect 28172 11160 28224 11169
rect 25504 11092 25556 11144
rect 27252 11092 27304 11144
rect 38292 11135 38344 11144
rect 38292 11101 38301 11135
rect 38301 11101 38335 11135
rect 38335 11101 38344 11135
rect 38292 11092 38344 11101
rect 28540 11024 28592 11076
rect 23756 10956 23808 11008
rect 25412 10956 25464 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 2320 10752 2372 10804
rect 4896 10752 4948 10804
rect 6736 10752 6788 10804
rect 13912 10752 13964 10804
rect 17684 10795 17736 10804
rect 17684 10761 17693 10795
rect 17693 10761 17727 10795
rect 17727 10761 17736 10795
rect 17684 10752 17736 10761
rect 1860 10727 1912 10736
rect 1860 10693 1869 10727
rect 1869 10693 1903 10727
rect 1903 10693 1912 10727
rect 1860 10684 1912 10693
rect 2412 10684 2464 10736
rect 3516 10659 3568 10668
rect 3516 10625 3525 10659
rect 3525 10625 3559 10659
rect 3559 10625 3568 10659
rect 3516 10616 3568 10625
rect 4804 10684 4856 10736
rect 6828 10684 6880 10736
rect 12992 10684 13044 10736
rect 4712 10616 4764 10668
rect 5632 10659 5684 10668
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 6552 10659 6604 10668
rect 6552 10625 6561 10659
rect 6561 10625 6595 10659
rect 6595 10625 6604 10659
rect 6552 10616 6604 10625
rect 13544 10616 13596 10668
rect 14556 10659 14608 10668
rect 14556 10625 14565 10659
rect 14565 10625 14599 10659
rect 14599 10625 14608 10659
rect 14556 10616 14608 10625
rect 24768 10752 24820 10804
rect 25872 10752 25924 10804
rect 2504 10548 2556 10600
rect 5356 10548 5408 10600
rect 3608 10480 3660 10532
rect 3240 10412 3292 10464
rect 11888 10412 11940 10464
rect 17776 10412 17828 10464
rect 18696 10616 18748 10668
rect 20720 10659 20772 10668
rect 20720 10625 20729 10659
rect 20729 10625 20763 10659
rect 20763 10625 20772 10659
rect 20720 10616 20772 10625
rect 22008 10659 22060 10668
rect 22008 10625 22017 10659
rect 22017 10625 22051 10659
rect 22051 10625 22060 10659
rect 22008 10616 22060 10625
rect 23480 10659 23532 10668
rect 19064 10591 19116 10600
rect 19064 10557 19073 10591
rect 19073 10557 19107 10591
rect 19107 10557 19116 10591
rect 19064 10548 19116 10557
rect 19432 10591 19484 10600
rect 19432 10557 19441 10591
rect 19441 10557 19475 10591
rect 19475 10557 19484 10591
rect 19432 10548 19484 10557
rect 23480 10625 23489 10659
rect 23489 10625 23523 10659
rect 23523 10625 23532 10659
rect 23480 10616 23532 10625
rect 25228 10684 25280 10736
rect 28356 10752 28408 10804
rect 24768 10659 24820 10668
rect 24768 10625 24777 10659
rect 24777 10625 24811 10659
rect 24811 10625 24820 10659
rect 24768 10616 24820 10625
rect 25412 10659 25464 10668
rect 25412 10625 25421 10659
rect 25421 10625 25455 10659
rect 25455 10625 25464 10659
rect 25412 10616 25464 10625
rect 27344 10616 27396 10668
rect 24308 10548 24360 10600
rect 20720 10480 20772 10532
rect 23848 10480 23900 10532
rect 25504 10480 25556 10532
rect 26332 10548 26384 10600
rect 29920 10548 29972 10600
rect 20076 10412 20128 10464
rect 20812 10455 20864 10464
rect 20812 10421 20821 10455
rect 20821 10421 20855 10455
rect 20855 10421 20864 10455
rect 20812 10412 20864 10421
rect 20904 10412 20956 10464
rect 22560 10412 22612 10464
rect 25412 10412 25464 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2228 10208 2280 10260
rect 3148 10208 3200 10260
rect 23572 10208 23624 10260
rect 24768 10208 24820 10260
rect 25228 10251 25280 10260
rect 25228 10217 25237 10251
rect 25237 10217 25271 10251
rect 25271 10217 25280 10251
rect 25228 10208 25280 10217
rect 13176 10140 13228 10192
rect 2044 10047 2096 10056
rect 2044 10013 2053 10047
rect 2053 10013 2087 10047
rect 2087 10013 2096 10047
rect 2044 10004 2096 10013
rect 2320 10004 2372 10056
rect 3700 10072 3752 10124
rect 17776 10115 17828 10124
rect 17776 10081 17785 10115
rect 17785 10081 17819 10115
rect 17819 10081 17828 10115
rect 17776 10072 17828 10081
rect 17868 10072 17920 10124
rect 20812 10072 20864 10124
rect 3424 10004 3476 10056
rect 7288 10004 7340 10056
rect 13820 9936 13872 9988
rect 15752 9979 15804 9988
rect 15752 9945 15761 9979
rect 15761 9945 15795 9979
rect 15795 9945 15804 9979
rect 15752 9936 15804 9945
rect 3700 9868 3752 9920
rect 5908 9911 5960 9920
rect 5908 9877 5917 9911
rect 5917 9877 5951 9911
rect 5951 9877 5960 9911
rect 17408 9936 17460 9988
rect 20720 10004 20772 10056
rect 23480 10140 23532 10192
rect 24308 10072 24360 10124
rect 28632 10072 28684 10124
rect 23848 10047 23900 10056
rect 23848 10013 23857 10047
rect 23857 10013 23891 10047
rect 23891 10013 23900 10047
rect 23848 10004 23900 10013
rect 25412 10047 25464 10056
rect 25412 10013 25421 10047
rect 25421 10013 25455 10047
rect 25455 10013 25464 10047
rect 25412 10004 25464 10013
rect 37188 10004 37240 10056
rect 19248 9936 19300 9988
rect 18696 9911 18748 9920
rect 5908 9868 5960 9877
rect 18696 9877 18705 9911
rect 18705 9877 18739 9911
rect 18739 9877 18748 9911
rect 18696 9868 18748 9877
rect 20720 9868 20772 9920
rect 22560 9979 22612 9988
rect 22560 9945 22569 9979
rect 22569 9945 22603 9979
rect 22603 9945 22612 9979
rect 22560 9936 22612 9945
rect 25688 9868 25740 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 1860 9664 1912 9716
rect 19064 9664 19116 9716
rect 2136 9596 2188 9648
rect 2872 9596 2924 9648
rect 3792 9639 3844 9648
rect 3792 9605 3801 9639
rect 3801 9605 3835 9639
rect 3835 9605 3844 9639
rect 3792 9596 3844 9605
rect 14740 9596 14792 9648
rect 17132 9639 17184 9648
rect 17132 9605 17141 9639
rect 17141 9605 17175 9639
rect 17175 9605 17184 9639
rect 17132 9596 17184 9605
rect 19432 9596 19484 9648
rect 20904 9664 20956 9716
rect 20720 9639 20772 9648
rect 20720 9605 20729 9639
rect 20729 9605 20763 9639
rect 20763 9605 20772 9639
rect 20720 9596 20772 9605
rect 24308 9596 24360 9648
rect 1124 9528 1176 9580
rect 2320 9571 2372 9580
rect 2320 9537 2329 9571
rect 2329 9537 2363 9571
rect 2363 9537 2372 9571
rect 2320 9528 2372 9537
rect 3056 9571 3108 9580
rect 3056 9537 3065 9571
rect 3065 9537 3099 9571
rect 3099 9537 3108 9571
rect 3056 9528 3108 9537
rect 3700 9571 3752 9580
rect 3700 9537 3709 9571
rect 3709 9537 3743 9571
rect 3743 9537 3752 9571
rect 3700 9528 3752 9537
rect 5632 9528 5684 9580
rect 14004 9528 14056 9580
rect 14464 9528 14516 9580
rect 18604 9571 18656 9580
rect 7932 9460 7984 9512
rect 15384 9460 15436 9512
rect 18604 9537 18613 9571
rect 18613 9537 18647 9571
rect 18647 9537 18656 9571
rect 18604 9528 18656 9537
rect 17684 9460 17736 9512
rect 20168 9528 20220 9580
rect 25228 9571 25280 9580
rect 25228 9537 25237 9571
rect 25237 9537 25271 9571
rect 25271 9537 25280 9571
rect 25228 9528 25280 9537
rect 25688 9571 25740 9580
rect 25688 9537 25697 9571
rect 25697 9537 25731 9571
rect 25731 9537 25740 9571
rect 25688 9528 25740 9537
rect 26332 9571 26384 9580
rect 26332 9537 26341 9571
rect 26341 9537 26375 9571
rect 26375 9537 26384 9571
rect 26332 9528 26384 9537
rect 27712 9528 27764 9580
rect 19432 9503 19484 9512
rect 19432 9469 19441 9503
rect 19441 9469 19475 9503
rect 19475 9469 19484 9503
rect 19432 9460 19484 9469
rect 19708 9392 19760 9444
rect 25320 9460 25372 9512
rect 26516 9460 26568 9512
rect 25964 9392 26016 9444
rect 37188 9460 37240 9512
rect 14464 9324 14516 9376
rect 19800 9324 19852 9376
rect 26240 9324 26292 9376
rect 26332 9324 26384 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 4620 9120 4672 9172
rect 17868 9163 17920 9172
rect 17868 9129 17877 9163
rect 17877 9129 17911 9163
rect 17911 9129 17920 9163
rect 17868 9120 17920 9129
rect 19800 9163 19852 9172
rect 19800 9129 19809 9163
rect 19809 9129 19843 9163
rect 19843 9129 19852 9163
rect 19800 9120 19852 9129
rect 25964 9163 26016 9172
rect 25964 9129 25973 9163
rect 25973 9129 26007 9163
rect 26007 9129 26016 9163
rect 25964 9120 26016 9129
rect 26516 9163 26568 9172
rect 26516 9129 26525 9163
rect 26525 9129 26559 9163
rect 26559 9129 26568 9163
rect 26516 9120 26568 9129
rect 2044 9095 2096 9104
rect 2044 9061 2053 9095
rect 2053 9061 2087 9095
rect 2087 9061 2096 9095
rect 2044 9052 2096 9061
rect 3056 9052 3108 9104
rect 9588 9052 9640 9104
rect 13544 9052 13596 9104
rect 4804 8984 4856 9036
rect 10968 8984 11020 9036
rect 3148 8959 3200 8968
rect 3148 8925 3157 8959
rect 3157 8925 3191 8959
rect 3191 8925 3200 8959
rect 3148 8916 3200 8925
rect 1584 8848 1636 8900
rect 4988 8848 5040 8900
rect 11244 8891 11296 8900
rect 11244 8857 11253 8891
rect 11253 8857 11287 8891
rect 11287 8857 11296 8891
rect 11244 8848 11296 8857
rect 11336 8891 11388 8900
rect 11336 8857 11345 8891
rect 11345 8857 11379 8891
rect 11379 8857 11388 8891
rect 15936 9027 15988 9036
rect 14464 8959 14516 8968
rect 14464 8925 14473 8959
rect 14473 8925 14507 8959
rect 14507 8925 14516 8959
rect 14464 8916 14516 8925
rect 15936 8993 15945 9027
rect 15945 8993 15979 9027
rect 15979 8993 15988 9027
rect 15936 8984 15988 8993
rect 16212 8984 16264 9036
rect 17776 8959 17828 8968
rect 11336 8848 11388 8857
rect 15476 8848 15528 8900
rect 16856 8780 16908 8832
rect 17776 8925 17785 8959
rect 17785 8925 17819 8959
rect 17819 8925 17828 8959
rect 17776 8916 17828 8925
rect 23296 8984 23348 9036
rect 23480 9027 23532 9036
rect 23480 8993 23489 9027
rect 23489 8993 23523 9027
rect 23523 8993 23532 9027
rect 23480 8984 23532 8993
rect 19064 8916 19116 8968
rect 22376 8959 22428 8968
rect 17684 8848 17736 8900
rect 22376 8925 22385 8959
rect 22385 8925 22419 8959
rect 22419 8925 22428 8959
rect 22376 8916 22428 8925
rect 25228 8916 25280 8968
rect 26240 8916 26292 8968
rect 35992 8959 36044 8968
rect 35992 8925 36001 8959
rect 36001 8925 36035 8959
rect 36035 8925 36044 8959
rect 35992 8916 36044 8925
rect 20260 8780 20312 8832
rect 27344 8848 27396 8900
rect 36452 8780 36504 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 1768 8619 1820 8628
rect 1768 8585 1777 8619
rect 1777 8585 1811 8619
rect 1811 8585 1820 8619
rect 1768 8576 1820 8585
rect 15384 8619 15436 8628
rect 15384 8585 15393 8619
rect 15393 8585 15427 8619
rect 15427 8585 15436 8619
rect 15384 8576 15436 8585
rect 15476 8576 15528 8628
rect 19156 8576 19208 8628
rect 27528 8576 27580 8628
rect 36912 8576 36964 8628
rect 1676 8508 1728 8560
rect 1492 8440 1544 8492
rect 1216 8372 1268 8424
rect 12164 8440 12216 8492
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 16212 8483 16264 8492
rect 2964 8372 3016 8424
rect 11152 8372 11204 8424
rect 15660 8304 15712 8356
rect 16212 8449 16221 8483
rect 16221 8449 16255 8483
rect 16255 8449 16264 8483
rect 16212 8440 16264 8449
rect 17224 8508 17276 8560
rect 25228 8508 25280 8560
rect 20076 8440 20128 8492
rect 26240 8440 26292 8492
rect 36452 8483 36504 8492
rect 36452 8449 36461 8483
rect 36461 8449 36495 8483
rect 36495 8449 36504 8483
rect 36452 8440 36504 8449
rect 38292 8483 38344 8492
rect 38292 8449 38301 8483
rect 38301 8449 38335 8483
rect 38335 8449 38344 8483
rect 38292 8440 38344 8449
rect 23480 8372 23532 8424
rect 23388 8304 23440 8356
rect 38016 8304 38068 8356
rect 12440 8279 12492 8288
rect 12440 8245 12449 8279
rect 12449 8245 12483 8279
rect 12483 8245 12492 8279
rect 12440 8236 12492 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 20536 8032 20588 8084
rect 11244 7964 11296 8016
rect 12164 7964 12216 8016
rect 3056 7896 3108 7948
rect 3608 7896 3660 7948
rect 5540 7828 5592 7880
rect 12440 7896 12492 7948
rect 14740 7939 14792 7948
rect 14740 7905 14749 7939
rect 14749 7905 14783 7939
rect 14783 7905 14792 7939
rect 14740 7896 14792 7905
rect 12072 7871 12124 7880
rect 12072 7837 12081 7871
rect 12081 7837 12115 7871
rect 12115 7837 12124 7871
rect 12072 7828 12124 7837
rect 13544 7760 13596 7812
rect 14832 7803 14884 7812
rect 14832 7769 14841 7803
rect 14841 7769 14875 7803
rect 14875 7769 14884 7803
rect 15660 7828 15712 7880
rect 17500 7828 17552 7880
rect 25596 7828 25648 7880
rect 27344 7871 27396 7880
rect 27344 7837 27353 7871
rect 27353 7837 27387 7871
rect 27387 7837 27396 7871
rect 27344 7828 27396 7837
rect 38292 7871 38344 7880
rect 38292 7837 38301 7871
rect 38301 7837 38335 7871
rect 38335 7837 38344 7871
rect 38292 7828 38344 7837
rect 14832 7760 14884 7769
rect 20076 7760 20128 7812
rect 21548 7803 21600 7812
rect 21548 7769 21557 7803
rect 21557 7769 21591 7803
rect 21591 7769 21600 7803
rect 21548 7760 21600 7769
rect 21640 7803 21692 7812
rect 21640 7769 21649 7803
rect 21649 7769 21683 7803
rect 21683 7769 21692 7803
rect 21640 7760 21692 7769
rect 22100 7760 22152 7812
rect 10324 7735 10376 7744
rect 10324 7701 10333 7735
rect 10333 7701 10367 7735
rect 10367 7701 10376 7735
rect 10324 7692 10376 7701
rect 12900 7692 12952 7744
rect 17868 7692 17920 7744
rect 19432 7692 19484 7744
rect 19984 7692 20036 7744
rect 26056 7760 26108 7812
rect 36360 7692 36412 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 1584 7531 1636 7540
rect 1584 7497 1593 7531
rect 1593 7497 1627 7531
rect 1627 7497 1636 7531
rect 1584 7488 1636 7497
rect 13544 7531 13596 7540
rect 13544 7497 13553 7531
rect 13553 7497 13587 7531
rect 13587 7497 13596 7531
rect 13544 7488 13596 7497
rect 14832 7488 14884 7540
rect 21548 7488 21600 7540
rect 2964 7463 3016 7472
rect 2964 7429 2973 7463
rect 2973 7429 3007 7463
rect 3007 7429 3016 7463
rect 2964 7420 3016 7429
rect 3240 7420 3292 7472
rect 5724 7420 5776 7472
rect 11888 7463 11940 7472
rect 11888 7429 11897 7463
rect 11897 7429 11931 7463
rect 11931 7429 11940 7463
rect 11888 7420 11940 7429
rect 18328 7463 18380 7472
rect 18328 7429 18337 7463
rect 18337 7429 18371 7463
rect 18371 7429 18380 7463
rect 18328 7420 18380 7429
rect 19156 7420 19208 7472
rect 19432 7420 19484 7472
rect 23480 7420 23532 7472
rect 1768 7395 1820 7404
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 1952 7352 2004 7404
rect 10968 7352 11020 7404
rect 11152 7395 11204 7404
rect 11152 7361 11161 7395
rect 11161 7361 11195 7395
rect 11195 7361 11204 7395
rect 11152 7352 11204 7361
rect 12900 7395 12952 7404
rect 12900 7361 12909 7395
rect 12909 7361 12943 7395
rect 12943 7361 12952 7395
rect 12900 7352 12952 7361
rect 14280 7352 14332 7404
rect 15568 7352 15620 7404
rect 22008 7395 22060 7404
rect 22008 7361 22017 7395
rect 22017 7361 22051 7395
rect 22051 7361 22060 7395
rect 22008 7352 22060 7361
rect 11796 7327 11848 7336
rect 11796 7293 11805 7327
rect 11805 7293 11839 7327
rect 11839 7293 11848 7327
rect 11796 7284 11848 7293
rect 12164 7327 12216 7336
rect 12164 7293 12173 7327
rect 12173 7293 12207 7327
rect 12207 7293 12216 7327
rect 12164 7284 12216 7293
rect 13084 7327 13136 7336
rect 13084 7293 13093 7327
rect 13093 7293 13127 7327
rect 13127 7293 13136 7327
rect 13084 7284 13136 7293
rect 17408 7327 17460 7336
rect 17408 7293 17417 7327
rect 17417 7293 17451 7327
rect 17451 7293 17460 7327
rect 17408 7284 17460 7293
rect 18236 7327 18288 7336
rect 18236 7293 18245 7327
rect 18245 7293 18279 7327
rect 18279 7293 18288 7327
rect 18236 7284 18288 7293
rect 19892 7284 19944 7336
rect 20076 7327 20128 7336
rect 20076 7293 20085 7327
rect 20085 7293 20119 7327
rect 20119 7293 20128 7327
rect 20076 7284 20128 7293
rect 24584 7284 24636 7336
rect 23572 7259 23624 7268
rect 23572 7225 23581 7259
rect 23581 7225 23615 7259
rect 23615 7225 23624 7259
rect 23572 7216 23624 7225
rect 3240 7148 3292 7200
rect 6736 7148 6788 7200
rect 11704 7148 11756 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 12072 6944 12124 6996
rect 23480 6987 23532 6996
rect 23480 6953 23489 6987
rect 23489 6953 23523 6987
rect 23523 6953 23532 6987
rect 23480 6944 23532 6953
rect 14740 6808 14792 6860
rect 17408 6808 17460 6860
rect 1768 6783 1820 6792
rect 1768 6749 1777 6783
rect 1777 6749 1811 6783
rect 1811 6749 1820 6783
rect 1768 6740 1820 6749
rect 3240 6783 3292 6792
rect 3240 6749 3249 6783
rect 3249 6749 3283 6783
rect 3283 6749 3292 6783
rect 3240 6740 3292 6749
rect 10324 6740 10376 6792
rect 11704 6783 11756 6792
rect 11704 6749 11713 6783
rect 11713 6749 11747 6783
rect 11747 6749 11756 6783
rect 11704 6740 11756 6749
rect 12348 6783 12400 6792
rect 12348 6749 12357 6783
rect 12357 6749 12391 6783
rect 12391 6749 12400 6783
rect 12348 6740 12400 6749
rect 14372 6740 14424 6792
rect 15660 6740 15712 6792
rect 17592 6740 17644 6792
rect 18236 6808 18288 6860
rect 20720 6740 20772 6792
rect 22376 6740 22428 6792
rect 1400 6604 1452 6656
rect 3056 6647 3108 6656
rect 3056 6613 3065 6647
rect 3065 6613 3099 6647
rect 3099 6613 3108 6647
rect 3056 6604 3108 6613
rect 6644 6647 6696 6656
rect 6644 6613 6653 6647
rect 6653 6613 6687 6647
rect 6687 6613 6696 6647
rect 6644 6604 6696 6613
rect 15016 6604 15068 6656
rect 19340 6604 19392 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 1952 6443 2004 6452
rect 1952 6409 1961 6443
rect 1961 6409 1995 6443
rect 1995 6409 2004 6443
rect 1952 6400 2004 6409
rect 11796 6400 11848 6452
rect 13084 6400 13136 6452
rect 15660 6443 15712 6452
rect 2872 6332 2924 6384
rect 6736 6307 6788 6316
rect 6736 6273 6745 6307
rect 6745 6273 6779 6307
rect 6779 6273 6788 6307
rect 6736 6264 6788 6273
rect 12992 6264 13044 6316
rect 15660 6409 15669 6443
rect 15669 6409 15703 6443
rect 15703 6409 15712 6443
rect 15660 6400 15712 6409
rect 17592 6443 17644 6452
rect 17592 6409 17601 6443
rect 17601 6409 17635 6443
rect 17635 6409 17644 6443
rect 17592 6400 17644 6409
rect 19432 6400 19484 6452
rect 24584 6400 24636 6452
rect 14004 6307 14056 6316
rect 14004 6273 14013 6307
rect 14013 6273 14047 6307
rect 14047 6273 14056 6307
rect 14004 6264 14056 6273
rect 15568 6307 15620 6316
rect 15568 6273 15577 6307
rect 15577 6273 15611 6307
rect 15611 6273 15620 6307
rect 15568 6264 15620 6273
rect 16580 6264 16632 6316
rect 25320 6264 25372 6316
rect 27528 6264 27580 6316
rect 38292 6307 38344 6316
rect 38292 6273 38301 6307
rect 38301 6273 38335 6307
rect 38335 6273 38344 6307
rect 38292 6264 38344 6273
rect 4068 6060 4120 6112
rect 25688 6060 25740 6112
rect 27436 6060 27488 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 14372 5899 14424 5908
rect 14372 5865 14381 5899
rect 14381 5865 14415 5899
rect 14415 5865 14424 5899
rect 14372 5856 14424 5865
rect 27712 5899 27764 5908
rect 27712 5865 27721 5899
rect 27721 5865 27755 5899
rect 27755 5865 27764 5899
rect 27712 5856 27764 5865
rect 2044 5831 2096 5840
rect 2044 5797 2053 5831
rect 2053 5797 2087 5831
rect 2087 5797 2096 5831
rect 2044 5788 2096 5797
rect 2504 5695 2556 5704
rect 2504 5661 2513 5695
rect 2513 5661 2547 5695
rect 2547 5661 2556 5695
rect 2504 5652 2556 5661
rect 12532 5652 12584 5704
rect 25688 5695 25740 5704
rect 25688 5661 25697 5695
rect 25697 5661 25731 5695
rect 25731 5661 25740 5695
rect 25688 5652 25740 5661
rect 30288 5652 30340 5704
rect 25228 5516 25280 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 6552 5312 6604 5364
rect 15752 5312 15804 5364
rect 16028 5244 16080 5296
rect 1768 5219 1820 5228
rect 1768 5185 1777 5219
rect 1777 5185 1811 5219
rect 1811 5185 1820 5219
rect 1768 5176 1820 5185
rect 18512 5108 18564 5160
rect 29920 5219 29972 5228
rect 29920 5185 29929 5219
rect 29929 5185 29963 5219
rect 29963 5185 29972 5219
rect 29920 5176 29972 5185
rect 38016 5219 38068 5228
rect 38016 5185 38025 5219
rect 38025 5185 38059 5219
rect 38059 5185 38068 5219
rect 38016 5176 38068 5185
rect 20536 5108 20588 5160
rect 31668 4972 31720 5024
rect 38200 5015 38252 5024
rect 38200 4981 38209 5015
rect 38209 4981 38243 5015
rect 38243 4981 38252 5015
rect 38200 4972 38252 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 37188 4768 37240 4820
rect 6644 4564 6696 4616
rect 38292 4607 38344 4616
rect 38292 4573 38301 4607
rect 38301 4573 38335 4607
rect 38335 4573 38344 4607
rect 38292 4564 38344 4573
rect 1768 4471 1820 4480
rect 1768 4437 1777 4471
rect 1777 4437 1811 4471
rect 1811 4437 1820 4471
rect 1768 4428 1820 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 37188 4156 37240 4208
rect 1400 4088 1452 4140
rect 5724 4088 5776 4140
rect 19432 4088 19484 4140
rect 20536 4131 20588 4140
rect 20536 4097 20545 4131
rect 20545 4097 20579 4131
rect 20579 4097 20588 4131
rect 20536 4088 20588 4097
rect 36360 4131 36412 4140
rect 36360 4097 36369 4131
rect 36369 4097 36403 4131
rect 36403 4097 36412 4131
rect 36360 4088 36412 4097
rect 18512 4020 18564 4072
rect 5632 3952 5684 4004
rect 21732 3952 21784 4004
rect 6736 3884 6788 3936
rect 21916 3884 21968 3936
rect 34796 3884 34848 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 21916 3519 21968 3528
rect 21916 3485 21925 3519
rect 21925 3485 21959 3519
rect 21959 3485 21968 3519
rect 21916 3476 21968 3485
rect 31668 3476 31720 3528
rect 37924 3476 37976 3528
rect 30564 3408 30616 3460
rect 1676 3383 1728 3392
rect 1676 3349 1685 3383
rect 1685 3349 1719 3383
rect 1719 3349 1728 3383
rect 1676 3340 1728 3349
rect 22652 3340 22704 3392
rect 33784 3340 33836 3392
rect 37464 3383 37516 3392
rect 37464 3349 37473 3383
rect 37473 3349 37507 3383
rect 37507 3349 37516 3383
rect 37464 3340 37516 3349
rect 38016 3340 38068 3392
rect 38200 3383 38252 3392
rect 38200 3349 38209 3383
rect 38209 3349 38243 3383
rect 38243 3349 38252 3383
rect 38200 3340 38252 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 3148 3136 3200 3188
rect 4068 3068 4120 3120
rect 35440 3136 35492 3188
rect 3056 3000 3108 3052
rect 6736 3043 6788 3052
rect 2780 2932 2832 2984
rect 6736 3009 6745 3043
rect 6745 3009 6779 3043
rect 6779 3009 6788 3043
rect 6736 3000 6788 3009
rect 9680 3000 9732 3052
rect 14188 3000 14240 3052
rect 17776 3000 17828 3052
rect 37464 3068 37516 3120
rect 37280 3000 37332 3052
rect 39304 3000 39356 3052
rect 20 2864 72 2916
rect 24492 2864 24544 2916
rect 27252 2864 27304 2916
rect 664 2796 716 2848
rect 6552 2839 6604 2848
rect 6552 2805 6561 2839
rect 6561 2805 6595 2839
rect 6595 2805 6604 2839
rect 6552 2796 6604 2805
rect 14924 2796 14976 2848
rect 17040 2839 17092 2848
rect 17040 2805 17049 2839
rect 17049 2805 17083 2839
rect 17083 2805 17092 2839
rect 17040 2796 17092 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 7288 2635 7340 2644
rect 7288 2601 7297 2635
rect 7297 2601 7331 2635
rect 7331 2601 7340 2635
rect 7288 2592 7340 2601
rect 12532 2592 12584 2644
rect 12992 2635 13044 2644
rect 12992 2601 13001 2635
rect 13001 2601 13035 2635
rect 13035 2601 13044 2635
rect 12992 2592 13044 2601
rect 16856 2635 16908 2644
rect 16856 2601 16865 2635
rect 16865 2601 16899 2635
rect 16899 2601 16908 2635
rect 16856 2592 16908 2601
rect 17500 2635 17552 2644
rect 17500 2601 17509 2635
rect 17509 2601 17543 2635
rect 17543 2601 17552 2635
rect 17500 2592 17552 2601
rect 19432 2635 19484 2644
rect 19432 2601 19441 2635
rect 19441 2601 19475 2635
rect 19475 2601 19484 2635
rect 19432 2592 19484 2601
rect 20720 2635 20772 2644
rect 20720 2601 20729 2635
rect 20729 2601 20763 2635
rect 20763 2601 20772 2635
rect 20720 2592 20772 2601
rect 22008 2635 22060 2644
rect 22008 2601 22017 2635
rect 22017 2601 22051 2635
rect 22051 2601 22060 2635
rect 22008 2592 22060 2601
rect 26240 2592 26292 2644
rect 27344 2592 27396 2644
rect 10416 2524 10468 2576
rect 12348 2524 12400 2576
rect 13268 2524 13320 2576
rect 3884 2388 3936 2440
rect 9312 2456 9364 2508
rect 18604 2456 18656 2508
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 6552 2431 6604 2440
rect 6552 2397 6561 2431
rect 6561 2397 6595 2431
rect 6595 2397 6604 2431
rect 6552 2388 6604 2397
rect 7104 2388 7156 2440
rect 8392 2388 8444 2440
rect 10968 2388 11020 2440
rect 11612 2388 11664 2440
rect 12900 2388 12952 2440
rect 14924 2431 14976 2440
rect 14924 2397 14933 2431
rect 14933 2397 14967 2431
rect 14967 2397 14976 2431
rect 14924 2388 14976 2397
rect 16120 2388 16172 2440
rect 17408 2388 17460 2440
rect 17868 2388 17920 2440
rect 19340 2388 19392 2440
rect 20628 2388 20680 2440
rect 21916 2388 21968 2440
rect 22652 2431 22704 2440
rect 22652 2397 22661 2431
rect 22661 2397 22695 2431
rect 22695 2397 22704 2431
rect 22652 2388 22704 2397
rect 25596 2524 25648 2576
rect 30288 2592 30340 2644
rect 27528 2524 27580 2576
rect 34520 2524 34572 2576
rect 23388 2456 23440 2508
rect 23848 2388 23900 2440
rect 25228 2431 25280 2440
rect 25228 2397 25237 2431
rect 25237 2397 25271 2431
rect 25271 2397 25280 2431
rect 25228 2388 25280 2397
rect 27068 2388 27120 2440
rect 28356 2388 28408 2440
rect 30288 2388 30340 2440
rect 31576 2388 31628 2440
rect 34796 2456 34848 2508
rect 37740 2499 37792 2508
rect 37740 2465 37749 2499
rect 37749 2465 37783 2499
rect 37783 2465 37792 2499
rect 37740 2456 37792 2465
rect 33784 2388 33836 2440
rect 1952 2252 2004 2304
rect 3240 2295 3292 2304
rect 3240 2261 3249 2295
rect 3249 2261 3283 2295
rect 3283 2261 3292 2295
rect 3240 2252 3292 2261
rect 5172 2252 5224 2304
rect 6460 2252 6512 2304
rect 14832 2252 14884 2304
rect 18052 2252 18104 2304
rect 22560 2252 22612 2304
rect 29828 2320 29880 2372
rect 25044 2252 25096 2304
rect 25136 2252 25188 2304
rect 25780 2252 25832 2304
rect 29644 2252 29696 2304
rect 32864 2320 32916 2372
rect 36728 2388 36780 2440
rect 33508 2252 33560 2304
rect 34796 2252 34848 2304
rect 36084 2252 36136 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 5264 2048 5316 2100
rect 17040 2048 17092 2100
rect 24400 2048 24452 2100
rect 29828 2048 29880 2100
<< metal2 >>
rect 18 39200 74 39800
rect 1306 39200 1362 39800
rect 2594 39200 2650 39800
rect 3238 39200 3294 39800
rect 4526 39200 4582 39800
rect 5814 39200 5870 39800
rect 6458 39200 6514 39800
rect 7746 39200 7802 39800
rect 9034 39200 9090 39800
rect 9678 39200 9734 39800
rect 10966 39200 11022 39800
rect 12254 39200 12310 39800
rect 13542 39200 13598 39800
rect 14186 39200 14242 39800
rect 15474 39200 15530 39800
rect 16762 39200 16818 39800
rect 17406 39200 17462 39800
rect 18694 39200 18750 39800
rect 19982 39200 20038 39800
rect 21270 39200 21326 39800
rect 21914 39200 21970 39800
rect 23202 39200 23258 39800
rect 24490 39200 24546 39800
rect 25134 39200 25190 39800
rect 26422 39200 26478 39800
rect 27710 39200 27766 39800
rect 28354 39200 28410 39800
rect 29642 39200 29698 39800
rect 30930 39200 30986 39800
rect 32218 39200 32274 39800
rect 32862 39200 32918 39800
rect 34150 39200 34206 39800
rect 35438 39200 35494 39800
rect 35544 39222 35848 39250
rect 32 36854 60 39200
rect 20 36848 72 36854
rect 20 36790 72 36796
rect 1320 36174 1348 39200
rect 1582 38856 1638 38865
rect 1582 38791 1638 38800
rect 1596 37330 1624 38791
rect 1766 38176 1822 38185
rect 1766 38111 1822 38120
rect 1584 37324 1636 37330
rect 1584 37266 1636 37272
rect 1780 36922 1808 38111
rect 2608 37210 2636 39200
rect 3252 37262 3280 39200
rect 4540 37754 4568 39200
rect 4540 37726 4660 37754
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4632 37262 4660 37726
rect 5828 37262 5856 39200
rect 5908 37460 5960 37466
rect 5908 37402 5960 37408
rect 2872 37256 2924 37262
rect 2608 37182 2820 37210
rect 2872 37198 2924 37204
rect 3240 37256 3292 37262
rect 3240 37198 3292 37204
rect 4620 37256 4672 37262
rect 4620 37198 4672 37204
rect 5816 37256 5868 37262
rect 5816 37198 5868 37204
rect 2792 37126 2820 37182
rect 2780 37120 2832 37126
rect 2780 37062 2832 37068
rect 1768 36916 1820 36922
rect 1768 36858 1820 36864
rect 1584 36780 1636 36786
rect 1584 36722 1636 36728
rect 1596 36417 1624 36722
rect 1582 36408 1638 36417
rect 1582 36343 1638 36352
rect 1308 36168 1360 36174
rect 1308 36110 1360 36116
rect 2688 36032 2740 36038
rect 2688 35974 2740 35980
rect 1584 35624 1636 35630
rect 1584 35566 1636 35572
rect 1596 34542 1624 35566
rect 1766 35456 1822 35465
rect 1766 35391 1822 35400
rect 1780 35290 1808 35391
rect 1768 35284 1820 35290
rect 1768 35226 1820 35232
rect 2700 35086 2728 35974
rect 2688 35080 2740 35086
rect 2688 35022 2740 35028
rect 1766 34776 1822 34785
rect 1766 34711 1822 34720
rect 1780 34610 1808 34711
rect 1768 34604 1820 34610
rect 1768 34546 1820 34552
rect 1584 34536 1636 34542
rect 1584 34478 1636 34484
rect 1596 33522 1624 34478
rect 2410 34096 2466 34105
rect 2410 34031 2466 34040
rect 2424 33998 2452 34031
rect 2412 33992 2464 33998
rect 2412 33934 2464 33940
rect 2504 33992 2556 33998
rect 2504 33934 2556 33940
rect 1768 33856 1820 33862
rect 1768 33798 1820 33804
rect 1860 33856 1912 33862
rect 1860 33798 1912 33804
rect 1584 33516 1636 33522
rect 1584 33458 1636 33464
rect 1780 33425 1808 33798
rect 1766 33416 1822 33425
rect 1766 33351 1822 33360
rect 1676 32428 1728 32434
rect 1676 32370 1728 32376
rect 1688 32065 1716 32370
rect 1674 32056 1730 32065
rect 1674 31991 1730 32000
rect 1872 31822 1900 33798
rect 2516 33114 2544 33934
rect 2504 33108 2556 33114
rect 2504 33050 2556 33056
rect 2228 32292 2280 32298
rect 2228 32234 2280 32240
rect 1860 31816 1912 31822
rect 1860 31758 1912 31764
rect 1768 31680 1820 31686
rect 1768 31622 1820 31628
rect 1780 31385 1808 31622
rect 1766 31376 1822 31385
rect 1766 31311 1822 31320
rect 1584 30252 1636 30258
rect 1584 30194 1636 30200
rect 1596 29073 1624 30194
rect 1768 30048 1820 30054
rect 1766 30016 1768 30025
rect 1820 30016 1822 30025
rect 1766 29951 1822 29960
rect 1768 29164 1820 29170
rect 1768 29106 1820 29112
rect 1582 29064 1638 29073
rect 1582 28999 1638 29008
rect 1780 28665 1808 29106
rect 1860 28960 1912 28966
rect 1860 28902 1912 28908
rect 1766 28656 1822 28665
rect 1766 28591 1822 28600
rect 1872 28558 1900 28902
rect 1860 28552 1912 28558
rect 1860 28494 1912 28500
rect 2136 28416 2188 28422
rect 2136 28358 2188 28364
rect 1584 27464 1636 27470
rect 1584 27406 1636 27412
rect 1596 26353 1624 27406
rect 1768 27328 1820 27334
rect 1766 27296 1768 27305
rect 1820 27296 1822 27305
rect 1766 27231 1822 27240
rect 1768 26988 1820 26994
rect 1768 26930 1820 26936
rect 1780 26625 1808 26930
rect 1766 26616 1822 26625
rect 1766 26551 1822 26560
rect 2148 26450 2176 28358
rect 2136 26444 2188 26450
rect 2136 26386 2188 26392
rect 1582 26344 1638 26353
rect 1582 26279 1638 26288
rect 1952 25968 2004 25974
rect 1952 25910 2004 25916
rect 1676 25288 1728 25294
rect 1674 25256 1676 25265
rect 1728 25256 1730 25265
rect 1674 25191 1730 25200
rect 1768 24812 1820 24818
rect 1768 24754 1820 24760
rect 1216 24608 1268 24614
rect 1216 24550 1268 24556
rect 1124 24132 1176 24138
rect 1124 24074 1176 24080
rect 1136 9586 1164 24074
rect 1124 9580 1176 9586
rect 1124 9522 1176 9528
rect 1228 8430 1256 24550
rect 1780 23905 1808 24754
rect 1964 24138 1992 25910
rect 1952 24132 2004 24138
rect 1952 24074 2004 24080
rect 2044 24064 2096 24070
rect 2044 24006 2096 24012
rect 1766 23896 1822 23905
rect 1766 23831 1822 23840
rect 1492 23520 1544 23526
rect 1492 23462 1544 23468
rect 1400 22704 1452 22710
rect 1400 22646 1452 22652
rect 1412 19258 1440 22646
rect 1320 19230 1440 19258
rect 1320 18970 1348 19230
rect 1308 18964 1360 18970
rect 1308 18906 1360 18912
rect 1320 11150 1348 18906
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1308 11144 1360 11150
rect 1308 11086 1360 11092
rect 1216 8424 1268 8430
rect 1216 8366 1268 8372
rect 1412 6662 1440 13874
rect 1504 8498 1532 23462
rect 1584 23112 1636 23118
rect 1584 23054 1636 23060
rect 1596 22574 1624 23054
rect 2056 23050 2084 24006
rect 2044 23044 2096 23050
rect 2044 22986 2096 22992
rect 1584 22568 1636 22574
rect 1584 22510 1636 22516
rect 1596 20398 1624 22510
rect 1676 21956 1728 21962
rect 1676 21898 1728 21904
rect 1688 21865 1716 21898
rect 1674 21856 1730 21865
rect 1674 21791 1730 21800
rect 1676 20868 1728 20874
rect 1676 20810 1728 20816
rect 1688 20505 1716 20810
rect 1674 20496 1730 20505
rect 1674 20431 1730 20440
rect 1768 20460 1820 20466
rect 1768 20402 1820 20408
rect 1584 20392 1636 20398
rect 1584 20334 1636 20340
rect 1596 19854 1624 20334
rect 1584 19848 1636 19854
rect 1584 19790 1636 19796
rect 1596 19310 1624 19790
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1596 18766 1624 19246
rect 1780 19145 1808 20402
rect 1766 19136 1822 19145
rect 1766 19071 1822 19080
rect 1584 18760 1636 18766
rect 1584 18702 1636 18708
rect 1596 17746 1624 18702
rect 1674 18456 1730 18465
rect 1674 18391 1730 18400
rect 1688 18358 1716 18391
rect 1676 18352 1728 18358
rect 1676 18294 1728 18300
rect 1584 17740 1636 17746
rect 1584 17682 1636 17688
rect 1676 17196 1728 17202
rect 1676 17138 1728 17144
rect 1688 17105 1716 17138
rect 1674 17096 1730 17105
rect 1674 17031 1730 17040
rect 1860 17060 1912 17066
rect 1860 17002 1912 17008
rect 1952 17060 2004 17066
rect 1952 17002 2004 17008
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1780 15745 1808 15846
rect 1766 15736 1822 15745
rect 1872 15706 1900 17002
rect 1964 16658 1992 17002
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 1766 15671 1822 15680
rect 1860 15700 1912 15706
rect 1860 15642 1912 15648
rect 1860 15360 1912 15366
rect 1860 15302 1912 15308
rect 1674 13696 1730 13705
rect 1674 13631 1730 13640
rect 1688 13326 1716 13631
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1584 8900 1636 8906
rect 1584 8842 1636 8848
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 1596 7546 1624 8842
rect 1688 8566 1716 12718
rect 1768 12368 1820 12374
rect 1766 12336 1768 12345
rect 1820 12336 1822 12345
rect 1766 12271 1822 12280
rect 1872 11354 1900 15302
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1860 10736 1912 10742
rect 1860 10678 1912 10684
rect 1872 9722 1900 10678
rect 1860 9716 1912 9722
rect 1860 9658 1912 9664
rect 1766 8936 1822 8945
rect 1766 8871 1822 8880
rect 1780 8634 1808 8871
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1676 8560 1728 8566
rect 1676 8502 1728 8508
rect 1766 7576 1822 7585
rect 1584 7540 1636 7546
rect 1766 7511 1822 7520
rect 1584 7482 1636 7488
rect 1780 7410 1808 7511
rect 1964 7410 1992 16594
rect 2056 10062 2084 22986
rect 2136 20256 2188 20262
rect 2136 20198 2188 20204
rect 2148 16726 2176 20198
rect 2136 16720 2188 16726
rect 2136 16662 2188 16668
rect 2240 16017 2268 32234
rect 2320 31816 2372 31822
rect 2412 31816 2464 31822
rect 2320 31758 2372 31764
rect 2410 31784 2412 31793
rect 2464 31784 2466 31793
rect 2332 27130 2360 31758
rect 2410 31719 2466 31728
rect 2780 30728 2832 30734
rect 2780 30670 2832 30676
rect 2792 29238 2820 30670
rect 2780 29232 2832 29238
rect 2780 29174 2832 29180
rect 2792 28014 2820 29174
rect 2780 28008 2832 28014
rect 2780 27950 2832 27956
rect 2884 27674 2912 37198
rect 4712 37188 4764 37194
rect 4712 37130 4764 37136
rect 4620 37120 4672 37126
rect 4620 37062 4672 37068
rect 3330 36816 3386 36825
rect 2964 36780 3016 36786
rect 3330 36751 3386 36760
rect 3976 36780 4028 36786
rect 2964 36722 3016 36728
rect 2976 36378 3004 36722
rect 3056 36576 3108 36582
rect 3056 36518 3108 36524
rect 2964 36372 3016 36378
rect 2964 36314 3016 36320
rect 3068 36310 3096 36518
rect 3056 36304 3108 36310
rect 3056 36246 3108 36252
rect 3240 35760 3292 35766
rect 3240 35702 3292 35708
rect 3252 34202 3280 35702
rect 3240 34196 3292 34202
rect 3240 34138 3292 34144
rect 2872 27668 2924 27674
rect 2872 27610 2924 27616
rect 3344 27130 3372 36751
rect 3976 36722 4028 36728
rect 3988 36378 4016 36722
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4632 36378 4660 37062
rect 3976 36372 4028 36378
rect 3976 36314 4028 36320
rect 4620 36372 4672 36378
rect 4620 36314 4672 36320
rect 4160 36168 4212 36174
rect 4160 36110 4212 36116
rect 4172 35630 4200 36110
rect 4160 35624 4212 35630
rect 4160 35566 4212 35572
rect 4620 35624 4672 35630
rect 4620 35566 4672 35572
rect 4172 35494 4200 35566
rect 4160 35488 4212 35494
rect 4160 35430 4212 35436
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4632 35154 4660 35566
rect 4620 35148 4672 35154
rect 4620 35090 4672 35096
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4068 33584 4120 33590
rect 4066 33552 4068 33561
rect 4120 33552 4122 33561
rect 4066 33487 4122 33496
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4724 31754 4752 37130
rect 4804 36712 4856 36718
rect 4804 36654 4856 36660
rect 4816 36242 4844 36654
rect 4896 36576 4948 36582
rect 4896 36518 4948 36524
rect 4804 36236 4856 36242
rect 4804 36178 4856 36184
rect 4908 36106 4936 36518
rect 5920 36242 5948 37402
rect 6472 37262 6500 39200
rect 6920 37392 6972 37398
rect 6920 37334 6972 37340
rect 6460 37256 6512 37262
rect 6460 37198 6512 37204
rect 6552 37120 6604 37126
rect 6552 37062 6604 37068
rect 6564 36922 6592 37062
rect 6552 36916 6604 36922
rect 6552 36858 6604 36864
rect 6932 36582 6960 37334
rect 7760 37126 7788 39200
rect 8760 37392 8812 37398
rect 8760 37334 8812 37340
rect 8392 37256 8444 37262
rect 8392 37198 8444 37204
rect 7748 37120 7800 37126
rect 7748 37062 7800 37068
rect 7932 36848 7984 36854
rect 7932 36790 7984 36796
rect 6460 36576 6512 36582
rect 6460 36518 6512 36524
rect 6920 36576 6972 36582
rect 6920 36518 6972 36524
rect 5908 36236 5960 36242
rect 5908 36178 5960 36184
rect 5920 36122 5948 36178
rect 4896 36100 4948 36106
rect 4896 36042 4948 36048
rect 4988 36100 5040 36106
rect 4988 36042 5040 36048
rect 5828 36094 5948 36122
rect 6472 36106 6500 36518
rect 7944 36378 7972 36790
rect 8300 36780 8352 36786
rect 8300 36722 8352 36728
rect 7932 36372 7984 36378
rect 7932 36314 7984 36320
rect 8312 36106 8340 36722
rect 6460 36100 6512 36106
rect 4896 35012 4948 35018
rect 4896 34954 4948 34960
rect 4908 34921 4936 34954
rect 4894 34912 4950 34921
rect 4894 34847 4950 34856
rect 5000 34406 5028 36042
rect 5448 35624 5500 35630
rect 5448 35566 5500 35572
rect 4988 34400 5040 34406
rect 4988 34342 5040 34348
rect 5000 33318 5028 34342
rect 5460 34066 5488 35566
rect 5448 34060 5500 34066
rect 5448 34002 5500 34008
rect 5460 33658 5488 34002
rect 5448 33652 5500 33658
rect 5448 33594 5500 33600
rect 5264 33448 5316 33454
rect 5264 33390 5316 33396
rect 4988 33312 5040 33318
rect 4988 33254 5040 33260
rect 4724 31726 4844 31754
rect 3608 31680 3660 31686
rect 3608 31622 3660 31628
rect 3620 31414 3648 31622
rect 3608 31408 3660 31414
rect 3608 31350 3660 31356
rect 3424 28484 3476 28490
rect 3424 28426 3476 28432
rect 2320 27124 2372 27130
rect 2320 27066 2372 27072
rect 3332 27124 3384 27130
rect 3332 27066 3384 27072
rect 2964 26580 3016 26586
rect 2964 26522 3016 26528
rect 2976 25906 3004 26522
rect 3056 26308 3108 26314
rect 3056 26250 3108 26256
rect 3068 26042 3096 26250
rect 3056 26036 3108 26042
rect 3056 25978 3108 25984
rect 2964 25900 3016 25906
rect 2964 25842 3016 25848
rect 2688 25220 2740 25226
rect 2688 25162 2740 25168
rect 2700 24410 2728 25162
rect 2688 24404 2740 24410
rect 2688 24346 2740 24352
rect 2504 24132 2556 24138
rect 2504 24074 2556 24080
rect 2516 19666 2544 24074
rect 2780 23724 2832 23730
rect 2780 23666 2832 23672
rect 2688 23520 2740 23526
rect 2688 23462 2740 23468
rect 2424 19638 2544 19666
rect 2226 16008 2282 16017
rect 2226 15943 2282 15952
rect 2320 15564 2372 15570
rect 2320 15506 2372 15512
rect 2136 14340 2188 14346
rect 2136 14282 2188 14288
rect 2228 14340 2280 14346
rect 2228 14282 2280 14288
rect 2148 14074 2176 14282
rect 2136 14068 2188 14074
rect 2136 14010 2188 14016
rect 2136 12912 2188 12918
rect 2136 12854 2188 12860
rect 2044 10056 2096 10062
rect 2044 9998 2096 10004
rect 2148 9654 2176 12854
rect 2240 10266 2268 14282
rect 2332 12714 2360 15506
rect 2320 12708 2372 12714
rect 2320 12650 2372 12656
rect 2424 12442 2452 19638
rect 2596 18216 2648 18222
rect 2596 18158 2648 18164
rect 2608 17746 2636 18158
rect 2596 17740 2648 17746
rect 2596 17682 2648 17688
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 2516 15065 2544 17138
rect 2596 16516 2648 16522
rect 2596 16458 2648 16464
rect 2502 15056 2558 15065
rect 2502 14991 2558 15000
rect 2504 14884 2556 14890
rect 2504 14826 2556 14832
rect 2516 14482 2544 14826
rect 2504 14476 2556 14482
rect 2504 14418 2556 14424
rect 2412 12436 2464 12442
rect 2412 12378 2464 12384
rect 2412 12300 2464 12306
rect 2412 12242 2464 12248
rect 2318 11928 2374 11937
rect 2318 11863 2374 11872
rect 2332 11830 2360 11863
rect 2320 11824 2372 11830
rect 2320 11766 2372 11772
rect 2424 11762 2452 12242
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2516 11626 2544 14418
rect 2608 13530 2636 16458
rect 2700 13841 2728 23462
rect 2792 23225 2820 23666
rect 2872 23656 2924 23662
rect 2872 23598 2924 23604
rect 2778 23216 2834 23225
rect 2778 23151 2834 23160
rect 2884 18222 2912 23598
rect 3436 22982 3464 28426
rect 3516 28008 3568 28014
rect 3516 27950 3568 27956
rect 3528 26586 3556 27950
rect 3516 26580 3568 26586
rect 3516 26522 3568 26528
rect 3424 22976 3476 22982
rect 3424 22918 3476 22924
rect 3148 22704 3200 22710
rect 3148 22646 3200 22652
rect 3056 20392 3108 20398
rect 3056 20334 3108 20340
rect 3068 18834 3096 20334
rect 3056 18828 3108 18834
rect 3056 18770 3108 18776
rect 2872 18216 2924 18222
rect 2872 18158 2924 18164
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2792 16658 2820 16730
rect 2780 16652 2832 16658
rect 2780 16594 2832 16600
rect 2780 15632 2832 15638
rect 2780 15574 2832 15580
rect 2792 14385 2820 15574
rect 2884 15065 2912 18158
rect 2964 16448 3016 16454
rect 2964 16390 3016 16396
rect 2976 16046 3004 16390
rect 2964 16040 3016 16046
rect 2964 15982 3016 15988
rect 2870 15056 2926 15065
rect 3160 15042 3188 22646
rect 3332 21956 3384 21962
rect 3332 21898 3384 21904
rect 3344 20058 3372 21898
rect 3332 20052 3384 20058
rect 3332 19994 3384 20000
rect 3240 19508 3292 19514
rect 3240 19450 3292 19456
rect 3252 17542 3280 19450
rect 3436 19417 3464 22918
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3332 18352 3384 18358
rect 3332 18294 3384 18300
rect 3240 17536 3292 17542
rect 3240 17478 3292 17484
rect 3252 17270 3280 17478
rect 3240 17264 3292 17270
rect 3240 17206 3292 17212
rect 3240 16992 3292 16998
rect 3240 16934 3292 16940
rect 2870 14991 2926 15000
rect 3068 15014 3188 15042
rect 2964 14952 3016 14958
rect 2964 14894 3016 14900
rect 2872 14408 2924 14414
rect 2778 14376 2834 14385
rect 2872 14350 2924 14356
rect 2778 14311 2834 14320
rect 2686 13832 2742 13841
rect 2686 13767 2742 13776
rect 2596 13524 2648 13530
rect 2596 13466 2648 13472
rect 2792 12442 2820 14311
rect 2884 13938 2912 14350
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2884 12850 2912 13874
rect 2976 13870 3004 14894
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 2780 12436 2832 12442
rect 2976 12434 3004 13262
rect 3068 12986 3096 15014
rect 3148 14952 3200 14958
rect 3148 14894 3200 14900
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 2976 12406 3096 12434
rect 2780 12378 2832 12384
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 2976 11898 3004 12174
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2872 11824 2924 11830
rect 2872 11766 2924 11772
rect 2504 11620 2556 11626
rect 2504 11562 2556 11568
rect 2320 11076 2372 11082
rect 2320 11018 2372 11024
rect 2412 11076 2464 11082
rect 2412 11018 2464 11024
rect 2332 10810 2360 11018
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 2424 10742 2452 11018
rect 2412 10736 2464 10742
rect 2412 10678 2464 10684
rect 2516 10606 2544 11562
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2320 10056 2372 10062
rect 2320 9998 2372 10004
rect 2136 9648 2188 9654
rect 2136 9590 2188 9596
rect 2332 9586 2360 9998
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2042 9208 2098 9217
rect 2042 9143 2098 9152
rect 2056 9110 2084 9143
rect 2044 9104 2096 9110
rect 2044 9046 2096 9052
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1766 6896 1822 6905
rect 1766 6831 1822 6840
rect 1780 6798 1808 6831
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 1400 6656 1452 6662
rect 1400 6598 1452 6604
rect 1950 6488 2006 6497
rect 1950 6423 1952 6432
rect 2004 6423 2006 6432
rect 1952 6394 2004 6400
rect 2042 5944 2098 5953
rect 2042 5879 2098 5888
rect 2056 5846 2084 5879
rect 2044 5840 2096 5846
rect 2044 5782 2096 5788
rect 2516 5710 2544 10542
rect 2884 9654 2912 11766
rect 3068 9738 3096 12406
rect 3160 10266 3188 14894
rect 3252 13326 3280 16934
rect 3344 15706 3372 18294
rect 3424 18216 3476 18222
rect 3424 18158 3476 18164
rect 3514 18184 3570 18193
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 3436 14074 3464 18158
rect 3514 18119 3570 18128
rect 3528 17626 3556 18119
rect 3620 17785 3648 31350
rect 4712 31136 4764 31142
rect 4712 31078 4764 31084
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4620 30592 4672 30598
rect 4620 30534 4672 30540
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4068 29232 4120 29238
rect 4066 29200 4068 29209
rect 4120 29200 4122 29209
rect 4066 29135 4122 29144
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 3884 28008 3936 28014
rect 3884 27950 3936 27956
rect 3896 25838 3924 27950
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4632 27062 4660 30534
rect 4724 28966 4752 31078
rect 4816 29646 4844 31726
rect 5276 30546 5304 33390
rect 5460 32502 5488 33594
rect 5828 32910 5856 36094
rect 6460 36042 6512 36048
rect 7380 36100 7432 36106
rect 7380 36042 7432 36048
rect 8300 36100 8352 36106
rect 8300 36042 8352 36048
rect 5908 36032 5960 36038
rect 7392 36009 7420 36042
rect 5908 35974 5960 35980
rect 7378 36000 7434 36009
rect 5920 35834 5948 35974
rect 7378 35935 7434 35944
rect 5908 35828 5960 35834
rect 5908 35770 5960 35776
rect 6828 35692 6880 35698
rect 6828 35634 6880 35640
rect 6840 35290 6868 35634
rect 8206 35592 8262 35601
rect 8206 35527 8262 35536
rect 8220 35494 8248 35527
rect 7012 35488 7064 35494
rect 7012 35430 7064 35436
rect 8208 35488 8260 35494
rect 8208 35430 8260 35436
rect 6828 35284 6880 35290
rect 6828 35226 6880 35232
rect 6920 34400 6972 34406
rect 6920 34342 6972 34348
rect 6932 34202 6960 34342
rect 6920 34196 6972 34202
rect 6920 34138 6972 34144
rect 5906 33960 5962 33969
rect 5906 33895 5908 33904
rect 5960 33895 5962 33904
rect 5908 33866 5960 33872
rect 5920 33658 5948 33866
rect 5908 33652 5960 33658
rect 5908 33594 5960 33600
rect 5816 32904 5868 32910
rect 5816 32846 5868 32852
rect 5448 32496 5500 32502
rect 5448 32438 5500 32444
rect 5460 31482 5488 32438
rect 6552 32428 6604 32434
rect 6552 32370 6604 32376
rect 5540 32224 5592 32230
rect 5540 32166 5592 32172
rect 5552 31890 5580 32166
rect 6092 32020 6144 32026
rect 6092 31962 6144 31968
rect 5540 31884 5592 31890
rect 5540 31826 5592 31832
rect 5448 31476 5500 31482
rect 5448 31418 5500 31424
rect 5356 31408 5408 31414
rect 5354 31376 5356 31385
rect 5408 31376 5410 31385
rect 5354 31311 5410 31320
rect 6104 30802 6132 31962
rect 5448 30796 5500 30802
rect 5448 30738 5500 30744
rect 6092 30796 6144 30802
rect 6092 30738 6144 30744
rect 5356 30728 5408 30734
rect 5354 30696 5356 30705
rect 5408 30696 5410 30705
rect 5354 30631 5410 30640
rect 5276 30518 5396 30546
rect 4804 29640 4856 29646
rect 4804 29582 4856 29588
rect 4712 28960 4764 28966
rect 4712 28902 4764 28908
rect 4620 27056 4672 27062
rect 4620 26998 4672 27004
rect 4632 26926 4660 26998
rect 4620 26920 4672 26926
rect 4620 26862 4672 26868
rect 4620 26784 4672 26790
rect 4620 26726 4672 26732
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 3884 25832 3936 25838
rect 3884 25774 3936 25780
rect 3792 23044 3844 23050
rect 3792 22986 3844 22992
rect 3700 18420 3752 18426
rect 3700 18362 3752 18368
rect 3606 17776 3662 17785
rect 3606 17711 3662 17720
rect 3528 17598 3648 17626
rect 3516 17536 3568 17542
rect 3516 17478 3568 17484
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 3344 13530 3372 13806
rect 3424 13796 3476 13802
rect 3424 13738 3476 13744
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3436 12850 3464 13738
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3436 12306 3464 12786
rect 3424 12300 3476 12306
rect 3424 12242 3476 12248
rect 3528 10674 3556 17478
rect 3620 16794 3648 17598
rect 3608 16788 3660 16794
rect 3608 16730 3660 16736
rect 3620 16046 3648 16730
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3620 14618 3648 14758
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 3712 14498 3740 18362
rect 3620 14470 3740 14498
rect 3620 12434 3648 14470
rect 3700 14000 3752 14006
rect 3700 13942 3752 13948
rect 3712 13530 3740 13942
rect 3700 13524 3752 13530
rect 3700 13466 3752 13472
rect 3804 12986 3832 22986
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3896 12850 3924 25774
rect 4632 25702 4660 26726
rect 4816 26234 4844 29582
rect 4896 29096 4948 29102
rect 4896 29038 4948 29044
rect 4908 28558 4936 29038
rect 5264 28960 5316 28966
rect 5264 28902 5316 28908
rect 4896 28552 4948 28558
rect 4896 28494 4948 28500
rect 4908 27878 4936 28494
rect 4988 28144 5040 28150
rect 4988 28086 5040 28092
rect 4896 27872 4948 27878
rect 4896 27814 4948 27820
rect 4908 27538 4936 27814
rect 5000 27713 5028 28086
rect 4986 27704 5042 27713
rect 4986 27639 5042 27648
rect 4896 27532 4948 27538
rect 4896 27474 4948 27480
rect 4896 26920 4948 26926
rect 4896 26862 4948 26868
rect 5080 26920 5132 26926
rect 5080 26862 5132 26868
rect 4724 26206 4844 26234
rect 4620 25696 4672 25702
rect 4620 25638 4672 25644
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 3976 25152 4028 25158
rect 3976 25094 4028 25100
rect 3988 19922 4016 25094
rect 4632 24750 4660 25638
rect 4620 24744 4672 24750
rect 4620 24686 4672 24692
rect 4068 24608 4120 24614
rect 4068 24550 4120 24556
rect 4080 24290 4108 24550
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4080 24262 4200 24290
rect 4632 24274 4660 24686
rect 4724 24614 4752 26206
rect 4712 24608 4764 24614
rect 4712 24550 4764 24556
rect 4172 23798 4200 24262
rect 4252 24268 4304 24274
rect 4252 24210 4304 24216
rect 4620 24268 4672 24274
rect 4620 24210 4672 24216
rect 4160 23792 4212 23798
rect 4160 23734 4212 23740
rect 4264 23730 4292 24210
rect 4528 24132 4580 24138
rect 4528 24074 4580 24080
rect 4252 23724 4304 23730
rect 4252 23666 4304 23672
rect 4540 23633 4568 24074
rect 4526 23624 4582 23633
rect 4526 23559 4582 23568
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23186 4660 24210
rect 4804 24132 4856 24138
rect 4804 24074 4856 24080
rect 4712 23860 4764 23866
rect 4712 23802 4764 23808
rect 4620 23180 4672 23186
rect 4620 23122 4672 23128
rect 4724 23066 4752 23802
rect 4632 23038 4752 23066
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3976 19916 4028 19922
rect 3976 19858 4028 19864
rect 4160 19712 4212 19718
rect 4160 19654 4212 19660
rect 4172 19446 4200 19654
rect 4252 19508 4304 19514
rect 4252 19450 4304 19456
rect 4160 19440 4212 19446
rect 4160 19382 4212 19388
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 4080 18850 4108 19314
rect 4160 19304 4212 19310
rect 4264 19258 4292 19450
rect 4212 19252 4292 19258
rect 4160 19246 4292 19252
rect 4172 19230 4292 19246
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4436 18896 4488 18902
rect 4080 18822 4200 18850
rect 4436 18838 4488 18844
rect 4172 18766 4200 18822
rect 4160 18760 4212 18766
rect 4160 18702 4212 18708
rect 4172 18170 4200 18702
rect 4448 18358 4476 18838
rect 4436 18352 4488 18358
rect 4436 18294 4488 18300
rect 4080 18142 4200 18170
rect 4080 17746 4108 18142
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4068 17740 4120 17746
rect 4068 17682 4120 17688
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 3976 16448 4028 16454
rect 3976 16390 4028 16396
rect 3988 16250 4016 16390
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 4080 15706 4108 16526
rect 4632 16522 4660 23038
rect 4712 22432 4764 22438
rect 4712 22374 4764 22380
rect 4724 21570 4752 22374
rect 4816 21706 4844 24074
rect 4908 21894 4936 26862
rect 5092 26353 5120 26862
rect 5172 26784 5224 26790
rect 5172 26726 5224 26732
rect 5078 26344 5134 26353
rect 5078 26279 5080 26288
rect 5132 26279 5134 26288
rect 5080 26250 5132 26256
rect 4988 25900 5040 25906
rect 4988 25842 5040 25848
rect 4896 21888 4948 21894
rect 4896 21830 4948 21836
rect 4816 21678 4936 21706
rect 4724 21542 4844 21570
rect 4816 21486 4844 21542
rect 4804 21480 4856 21486
rect 4804 21422 4856 21428
rect 4816 19446 4844 21422
rect 4804 19440 4856 19446
rect 4804 19382 4856 19388
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4724 18698 4752 19110
rect 4804 18828 4856 18834
rect 4804 18770 4856 18776
rect 4712 18692 4764 18698
rect 4712 18634 4764 18640
rect 4724 18426 4752 18634
rect 4712 18420 4764 18426
rect 4712 18362 4764 18368
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 4620 16516 4672 16522
rect 4620 16458 4672 16464
rect 4724 16153 4752 18158
rect 4710 16144 4766 16153
rect 4710 16079 4766 16088
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 3988 13734 4016 15438
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4080 14346 4108 14962
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14340 4120 14346
rect 4068 14282 4120 14288
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 3620 12406 3740 12434
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3620 11665 3648 11698
rect 3606 11656 3662 11665
rect 3606 11591 3662 11600
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3608 10532 3660 10538
rect 3608 10474 3660 10480
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 2976 9710 3096 9738
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 2976 8514 3004 9710
rect 3054 9616 3110 9625
rect 3054 9551 3056 9560
rect 3108 9551 3110 9560
rect 3056 9522 3108 9528
rect 3146 9480 3202 9489
rect 3146 9415 3202 9424
rect 3056 9104 3108 9110
rect 3056 9046 3108 9052
rect 2884 8486 3004 8514
rect 2884 6390 2912 8486
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2976 7478 3004 8366
rect 3068 7954 3096 9046
rect 3160 8974 3188 9415
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3056 7948 3108 7954
rect 3056 7890 3108 7896
rect 3252 7478 3280 10406
rect 3422 10296 3478 10305
rect 3422 10231 3478 10240
rect 3436 10062 3464 10231
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3620 9625 3648 10474
rect 3712 10130 3740 12406
rect 3792 12164 3844 12170
rect 3792 12106 3844 12112
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3606 9616 3662 9625
rect 3712 9586 3740 9862
rect 3804 9654 3832 12106
rect 3988 11218 4016 13670
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 4172 13190 4200 13262
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4632 12986 4660 15098
rect 4724 13530 4752 15982
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4816 13410 4844 18770
rect 4908 15162 4936 21678
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 4894 15056 4950 15065
rect 4894 14991 4950 15000
rect 4724 13382 4844 13410
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4620 12164 4672 12170
rect 4620 12106 4672 12112
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3606 9551 3662 9560
rect 3700 9580 3752 9586
rect 3620 7954 3648 9551
rect 3700 9522 3752 9528
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 9178 4660 12106
rect 4724 10674 4752 13382
rect 4908 12434 4936 14991
rect 5000 14074 5028 25842
rect 5184 23866 5212 26726
rect 5172 23860 5224 23866
rect 5172 23802 5224 23808
rect 5080 23180 5132 23186
rect 5080 23122 5132 23128
rect 5092 22098 5120 23122
rect 5080 22092 5132 22098
rect 5276 22094 5304 28902
rect 5368 22137 5396 30518
rect 5080 22034 5132 22040
rect 5184 22066 5304 22094
rect 5354 22128 5410 22137
rect 5080 21888 5132 21894
rect 5080 21830 5132 21836
rect 5092 17728 5120 21830
rect 5184 18873 5212 22066
rect 5354 22063 5410 22072
rect 5264 21956 5316 21962
rect 5264 21898 5316 21904
rect 5170 18864 5226 18873
rect 5170 18799 5226 18808
rect 5092 17700 5212 17728
rect 5080 17604 5132 17610
rect 5080 17546 5132 17552
rect 5092 16046 5120 17546
rect 5080 16040 5132 16046
rect 5080 15982 5132 15988
rect 5184 15892 5212 17700
rect 5276 16250 5304 21898
rect 5356 20256 5408 20262
rect 5356 20198 5408 20204
rect 5368 19514 5396 20198
rect 5356 19508 5408 19514
rect 5356 19450 5408 19456
rect 5368 18154 5396 19450
rect 5356 18148 5408 18154
rect 5356 18090 5408 18096
rect 5460 17728 5488 30738
rect 6104 30258 6132 30738
rect 6564 30326 6592 32370
rect 7024 31958 7052 35430
rect 8208 34468 8260 34474
rect 8208 34410 8260 34416
rect 7472 33516 7524 33522
rect 7472 33458 7524 33464
rect 7484 32978 7512 33458
rect 7472 32972 7524 32978
rect 7472 32914 7524 32920
rect 7012 31952 7064 31958
rect 7012 31894 7064 31900
rect 6184 30320 6236 30326
rect 6184 30262 6236 30268
rect 6552 30320 6604 30326
rect 6552 30262 6604 30268
rect 6092 30252 6144 30258
rect 6092 30194 6144 30200
rect 6196 29238 6224 30262
rect 7840 30048 7892 30054
rect 7840 29990 7892 29996
rect 6184 29232 6236 29238
rect 6184 29174 6236 29180
rect 7012 29164 7064 29170
rect 7012 29106 7064 29112
rect 6458 28520 6514 28529
rect 6458 28455 6460 28464
rect 6512 28455 6514 28464
rect 6460 28426 6512 28432
rect 5632 27396 5684 27402
rect 5632 27338 5684 27344
rect 5540 22704 5592 22710
rect 5540 22646 5592 22652
rect 5552 19938 5580 22646
rect 5644 20262 5672 27338
rect 5724 26920 5776 26926
rect 5724 26862 5776 26868
rect 6736 26920 6788 26926
rect 6736 26862 6788 26868
rect 5736 22094 5764 26862
rect 6748 26382 6776 26862
rect 7024 26450 7052 29106
rect 7104 27600 7156 27606
rect 7104 27542 7156 27548
rect 7012 26444 7064 26450
rect 7012 26386 7064 26392
rect 6736 26376 6788 26382
rect 7024 26353 7052 26386
rect 6736 26318 6788 26324
rect 7010 26344 7066 26353
rect 6748 25838 6776 26318
rect 7010 26279 7066 26288
rect 6736 25832 6788 25838
rect 6736 25774 6788 25780
rect 6748 25362 6776 25774
rect 6736 25356 6788 25362
rect 6736 25298 6788 25304
rect 6920 24812 6972 24818
rect 6920 24754 6972 24760
rect 6000 24744 6052 24750
rect 6000 24686 6052 24692
rect 6012 22438 6040 24686
rect 6932 24614 6960 24754
rect 6920 24608 6972 24614
rect 6920 24550 6972 24556
rect 6460 24404 6512 24410
rect 6460 24346 6512 24352
rect 6472 24290 6500 24346
rect 6288 24262 6500 24290
rect 6288 24206 6316 24262
rect 6276 24200 6328 24206
rect 6276 24142 6328 24148
rect 6368 24132 6420 24138
rect 6368 24074 6420 24080
rect 6380 23526 6408 24074
rect 6368 23520 6420 23526
rect 6368 23462 6420 23468
rect 6000 22432 6052 22438
rect 5998 22400 6000 22409
rect 6052 22400 6054 22409
rect 5998 22335 6054 22344
rect 5736 22066 6040 22094
rect 5816 21684 5868 21690
rect 5816 21626 5868 21632
rect 5632 20256 5684 20262
rect 5632 20198 5684 20204
rect 5552 19910 5672 19938
rect 5540 19780 5592 19786
rect 5540 19722 5592 19728
rect 5368 17700 5488 17728
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5092 15864 5212 15892
rect 5276 15881 5304 16050
rect 5262 15872 5318 15881
rect 4988 14068 5040 14074
rect 4988 14010 5040 14016
rect 5092 13258 5120 15864
rect 5262 15807 5318 15816
rect 5276 15722 5304 15807
rect 5184 15694 5304 15722
rect 5184 15026 5212 15694
rect 5264 15632 5316 15638
rect 5264 15574 5316 15580
rect 5172 15020 5224 15026
rect 5172 14962 5224 14968
rect 5172 14272 5224 14278
rect 5172 14214 5224 14220
rect 5080 13252 5132 13258
rect 5080 13194 5132 13200
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 4816 12406 4936 12434
rect 4816 10742 4844 12406
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 4908 10810 4936 11018
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4804 10736 4856 10742
rect 4804 10678 4856 10684
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4816 9042 4844 10678
rect 4804 9036 4856 9042
rect 4804 8978 4856 8984
rect 5000 8906 5028 12786
rect 5184 11218 5212 14214
rect 5276 13138 5304 15574
rect 5368 13326 5396 17700
rect 5552 16454 5580 19722
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5644 16266 5672 19910
rect 5724 19304 5776 19310
rect 5724 19246 5776 19252
rect 5736 18902 5764 19246
rect 5724 18896 5776 18902
rect 5724 18838 5776 18844
rect 5724 18692 5776 18698
rect 5724 18634 5776 18640
rect 5460 16238 5672 16266
rect 5460 16182 5488 16238
rect 5448 16176 5500 16182
rect 5448 16118 5500 16124
rect 5538 16144 5594 16153
rect 5538 16079 5594 16088
rect 5632 16108 5684 16114
rect 5446 15464 5502 15473
rect 5446 15399 5502 15408
rect 5460 15366 5488 15399
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5460 15026 5488 15302
rect 5448 15020 5500 15026
rect 5448 14962 5500 14968
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5460 14006 5488 14214
rect 5448 14000 5500 14006
rect 5448 13942 5500 13948
rect 5446 13696 5502 13705
rect 5446 13631 5502 13640
rect 5460 13326 5488 13631
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5552 13258 5580 16079
rect 5632 16050 5684 16056
rect 5644 15502 5672 16050
rect 5632 15496 5684 15502
rect 5632 15438 5684 15444
rect 5736 14550 5764 18634
rect 5828 15706 5856 21626
rect 5908 16448 5960 16454
rect 5908 16390 5960 16396
rect 5816 15700 5868 15706
rect 5816 15642 5868 15648
rect 5920 15502 5948 16390
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 5920 14958 5948 15438
rect 6012 15366 6040 22066
rect 6092 19780 6144 19786
rect 6092 19722 6144 19728
rect 6000 15360 6052 15366
rect 6000 15302 6052 15308
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5724 14544 5776 14550
rect 5724 14486 5776 14492
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 5540 13252 5592 13258
rect 5540 13194 5592 13200
rect 5276 13110 5396 13138
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5368 10606 5396 13110
rect 5538 12336 5594 12345
rect 5538 12271 5594 12280
rect 5552 12238 5580 12271
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3608 7948 3660 7954
rect 3608 7890 3660 7896
rect 5552 7886 5580 12174
rect 5644 11898 5672 14350
rect 5908 14340 5960 14346
rect 5908 14282 5960 14288
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5630 10976 5686 10985
rect 5630 10911 5686 10920
rect 5644 10674 5672 10911
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 3240 7472 3292 7478
rect 3240 7414 3292 7420
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3252 6798 3280 7142
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 2872 6384 2924 6390
rect 2872 6326 2924 6332
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 1766 5536 1822 5545
rect 1766 5471 1822 5480
rect 1780 5234 1808 5471
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 1768 4480 1820 4486
rect 1768 4422 1820 4428
rect 1780 4185 1808 4422
rect 1766 4176 1822 4185
rect 1400 4140 1452 4146
rect 1766 4111 1822 4120
rect 1400 4082 1452 4088
rect 1412 3505 1440 4082
rect 1398 3496 1454 3505
rect 1398 3431 1454 3440
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 20 2916 72 2922
rect 20 2858 72 2864
rect 32 800 60 2858
rect 664 2848 716 2854
rect 664 2790 716 2796
rect 676 800 704 2790
rect 1688 2145 1716 3334
rect 3068 3058 3096 6598
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 3146 3224 3202 3233
rect 3146 3159 3148 3168
rect 3200 3159 3202 3168
rect 3148 3130 3200 3136
rect 4080 3126 4108 6054
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 5644 4010 5672 9522
rect 5736 7478 5764 11494
rect 5920 9926 5948 14282
rect 6104 11150 6132 19722
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 6196 16114 6224 16526
rect 6276 16516 6328 16522
rect 6276 16458 6328 16464
rect 6288 16182 6316 16458
rect 6276 16176 6328 16182
rect 6276 16118 6328 16124
rect 6184 16108 6236 16114
rect 6184 16050 6236 16056
rect 6196 15502 6224 16050
rect 6276 15972 6328 15978
rect 6276 15914 6328 15920
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 6288 14958 6316 15914
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6184 14340 6236 14346
rect 6184 14282 6236 14288
rect 6196 13530 6224 14282
rect 6380 13938 6408 23462
rect 6736 23044 6788 23050
rect 6736 22986 6788 22992
rect 6552 21480 6604 21486
rect 6552 21422 6604 21428
rect 6564 21010 6592 21422
rect 6552 21004 6604 21010
rect 6552 20946 6604 20952
rect 6644 21004 6696 21010
rect 6644 20946 6696 20952
rect 6564 19922 6592 20946
rect 6552 19916 6604 19922
rect 6552 19858 6604 19864
rect 6564 19378 6592 19858
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 6460 18896 6512 18902
rect 6460 18838 6512 18844
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6472 12238 6500 18838
rect 6564 18834 6592 19314
rect 6656 18970 6684 20946
rect 6644 18964 6696 18970
rect 6644 18906 6696 18912
rect 6552 18828 6604 18834
rect 6552 18770 6604 18776
rect 6656 18714 6684 18906
rect 6564 18686 6684 18714
rect 6564 18358 6592 18686
rect 6644 18624 6696 18630
rect 6644 18566 6696 18572
rect 6552 18352 6604 18358
rect 6552 18294 6604 18300
rect 6656 16522 6684 18566
rect 6644 16516 6696 16522
rect 6644 16458 6696 16464
rect 6644 15904 6696 15910
rect 6644 15846 6696 15852
rect 6656 15094 6684 15846
rect 6748 15706 6776 22986
rect 6828 22568 6880 22574
rect 6828 22510 6880 22516
rect 6840 22098 6868 22510
rect 6828 22092 6880 22098
rect 6828 22034 6880 22040
rect 6932 21622 6960 24550
rect 7116 22094 7144 27542
rect 7564 26920 7616 26926
rect 7564 26862 7616 26868
rect 7576 26234 7604 26862
rect 7484 26206 7604 26234
rect 7484 22778 7512 26206
rect 7748 24336 7800 24342
rect 7748 24278 7800 24284
rect 7760 23798 7788 24278
rect 7748 23792 7800 23798
rect 7748 23734 7800 23740
rect 7564 22976 7616 22982
rect 7564 22918 7616 22924
rect 7472 22772 7524 22778
rect 7472 22714 7524 22720
rect 7116 22066 7236 22094
rect 6920 21616 6972 21622
rect 6920 21558 6972 21564
rect 6932 20534 6960 21558
rect 6920 20528 6972 20534
rect 6920 20470 6972 20476
rect 6920 19780 6972 19786
rect 6920 19722 6972 19728
rect 6736 15700 6788 15706
rect 6736 15642 6788 15648
rect 6932 15638 6960 19722
rect 7208 19310 7236 22066
rect 7472 20460 7524 20466
rect 7472 20402 7524 20408
rect 7380 19440 7432 19446
rect 7380 19382 7432 19388
rect 7196 19304 7248 19310
rect 7196 19246 7248 19252
rect 7288 18624 7340 18630
rect 7288 18566 7340 18572
rect 7196 18420 7248 18426
rect 7196 18362 7248 18368
rect 7012 17604 7064 17610
rect 7012 17546 7064 17552
rect 6920 15632 6972 15638
rect 6920 15574 6972 15580
rect 6828 15496 6880 15502
rect 6920 15496 6972 15502
rect 6828 15438 6880 15444
rect 6918 15464 6920 15473
rect 6972 15464 6974 15473
rect 6840 15094 6868 15438
rect 6918 15399 6974 15408
rect 6644 15088 6696 15094
rect 6644 15030 6696 15036
rect 6828 15088 6880 15094
rect 6828 15030 6880 15036
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 6748 13870 6776 14894
rect 7024 14482 7052 17546
rect 7208 15162 7236 18362
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 7300 15042 7328 18566
rect 7392 16250 7420 19382
rect 7484 16590 7512 20402
rect 7576 19174 7604 22918
rect 7748 21888 7800 21894
rect 7748 21830 7800 21836
rect 7760 21622 7788 21830
rect 7748 21616 7800 21622
rect 7748 21558 7800 21564
rect 7748 19780 7800 19786
rect 7748 19722 7800 19728
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7564 18692 7616 18698
rect 7564 18634 7616 18640
rect 7576 18290 7604 18634
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 7564 18148 7616 18154
rect 7564 18090 7616 18096
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7380 16244 7432 16250
rect 7380 16186 7432 16192
rect 7116 15014 7328 15042
rect 7012 14476 7064 14482
rect 7012 14418 7064 14424
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6472 11762 6500 12174
rect 6736 11824 6788 11830
rect 6736 11766 6788 11772
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6748 10810 6776 11766
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6840 11354 6868 11630
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6840 10742 6868 11290
rect 7116 11150 7144 15014
rect 7576 14414 7604 18090
rect 7668 17921 7696 19654
rect 7654 17912 7710 17921
rect 7654 17847 7710 17856
rect 7760 16250 7788 19722
rect 7852 18290 7880 29990
rect 8220 29714 8248 34410
rect 8208 29708 8260 29714
rect 8208 29650 8260 29656
rect 8024 27872 8076 27878
rect 8024 27814 8076 27820
rect 8036 27674 8064 27814
rect 8024 27668 8076 27674
rect 8024 27610 8076 27616
rect 8116 27668 8168 27674
rect 8116 27610 8168 27616
rect 7932 25900 7984 25906
rect 7932 25842 7984 25848
rect 7944 24614 7972 25842
rect 8024 25220 8076 25226
rect 8024 25162 8076 25168
rect 7932 24608 7984 24614
rect 7932 24550 7984 24556
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 7838 18184 7894 18193
rect 7838 18119 7894 18128
rect 7852 17202 7880 18119
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7932 16244 7984 16250
rect 7932 16186 7984 16192
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 7668 15434 7696 16050
rect 7944 16046 7972 16186
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 7656 15428 7708 15434
rect 7656 15370 7708 15376
rect 8036 15094 8064 25162
rect 8128 19718 8156 27610
rect 8404 26314 8432 37198
rect 8772 36718 8800 37334
rect 9048 37126 9076 39200
rect 9692 37126 9720 39200
rect 9956 37256 10008 37262
rect 9956 37198 10008 37204
rect 10048 37256 10100 37262
rect 10048 37198 10100 37204
rect 10980 37210 11008 39200
rect 11978 37360 12034 37369
rect 11978 37295 11980 37304
rect 12032 37295 12034 37304
rect 11980 37266 12032 37272
rect 12268 37262 12296 39200
rect 12256 37256 12308 37262
rect 9036 37120 9088 37126
rect 9036 37062 9088 37068
rect 9680 37120 9732 37126
rect 9680 37062 9732 37068
rect 9680 36780 9732 36786
rect 9680 36722 9732 36728
rect 8760 36712 8812 36718
rect 8760 36654 8812 36660
rect 8484 36372 8536 36378
rect 8484 36314 8536 36320
rect 8496 35154 8524 36314
rect 8668 35488 8720 35494
rect 8668 35430 8720 35436
rect 8484 35148 8536 35154
rect 8484 35090 8536 35096
rect 8496 33454 8524 35090
rect 8576 35080 8628 35086
rect 8576 35022 8628 35028
rect 8588 34746 8616 35022
rect 8576 34740 8628 34746
rect 8576 34682 8628 34688
rect 8680 34610 8708 35430
rect 8668 34604 8720 34610
rect 8668 34546 8720 34552
rect 8484 33448 8536 33454
rect 8484 33390 8536 33396
rect 8484 30592 8536 30598
rect 8484 30534 8536 30540
rect 8392 26308 8444 26314
rect 8392 26250 8444 26256
rect 8392 25832 8444 25838
rect 8392 25774 8444 25780
rect 8404 24818 8432 25774
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 8208 24064 8260 24070
rect 8208 24006 8260 24012
rect 8220 21146 8248 24006
rect 8300 22228 8352 22234
rect 8300 22170 8352 22176
rect 8208 21140 8260 21146
rect 8208 21082 8260 21088
rect 8116 19712 8168 19718
rect 8116 19654 8168 19660
rect 8208 19508 8260 19514
rect 8208 19450 8260 19456
rect 8116 19372 8168 19378
rect 8116 19314 8168 19320
rect 8128 19174 8156 19314
rect 8116 19168 8168 19174
rect 8116 19110 8168 19116
rect 8116 17604 8168 17610
rect 8116 17546 8168 17552
rect 8128 16794 8156 17546
rect 8116 16788 8168 16794
rect 8116 16730 8168 16736
rect 8128 16590 8156 16730
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 8220 16522 8248 19450
rect 8312 19174 8340 22170
rect 8496 22094 8524 30534
rect 8772 26234 8800 36654
rect 9404 36100 9456 36106
rect 9404 36042 9456 36048
rect 9220 36032 9272 36038
rect 9220 35974 9272 35980
rect 9128 35624 9180 35630
rect 9128 35566 9180 35572
rect 8942 35048 8998 35057
rect 8942 34983 8998 34992
rect 8956 34950 8984 34983
rect 8944 34944 8996 34950
rect 8944 34886 8996 34892
rect 9140 34066 9168 35566
rect 9232 35154 9260 35974
rect 9416 35766 9444 36042
rect 9404 35760 9456 35766
rect 9404 35702 9456 35708
rect 9416 35630 9444 35702
rect 9404 35624 9456 35630
rect 9404 35566 9456 35572
rect 9220 35148 9272 35154
rect 9220 35090 9272 35096
rect 9310 35048 9366 35057
rect 9310 34983 9312 34992
rect 9364 34983 9366 34992
rect 9312 34954 9364 34960
rect 9220 34944 9272 34950
rect 9218 34912 9220 34921
rect 9272 34912 9274 34921
rect 9218 34847 9274 34856
rect 9692 34066 9720 36722
rect 9864 35216 9916 35222
rect 9864 35158 9916 35164
rect 9876 35018 9904 35158
rect 9864 35012 9916 35018
rect 9864 34954 9916 34960
rect 9128 34060 9180 34066
rect 9128 34002 9180 34008
rect 9680 34060 9732 34066
rect 9680 34002 9732 34008
rect 9140 33590 9168 34002
rect 9588 33856 9640 33862
rect 9588 33798 9640 33804
rect 9128 33584 9180 33590
rect 9128 33526 9180 33532
rect 9036 33516 9088 33522
rect 9036 33458 9088 33464
rect 9048 33386 9076 33458
rect 9036 33380 9088 33386
rect 9036 33322 9088 33328
rect 9140 32434 9168 33526
rect 9496 33516 9548 33522
rect 9496 33458 9548 33464
rect 9128 32428 9180 32434
rect 9128 32370 9180 32376
rect 9140 31890 9168 32370
rect 9128 31884 9180 31890
rect 9128 31826 9180 31832
rect 9140 31142 9168 31826
rect 9312 31272 9364 31278
rect 9312 31214 9364 31220
rect 9128 31136 9180 31142
rect 9128 31078 9180 31084
rect 9324 30054 9352 31214
rect 9312 30048 9364 30054
rect 9312 29990 9364 29996
rect 9128 29640 9180 29646
rect 9128 29582 9180 29588
rect 9140 29170 9168 29582
rect 9128 29164 9180 29170
rect 9128 29106 9180 29112
rect 9324 28694 9352 29990
rect 9404 29572 9456 29578
rect 9404 29514 9456 29520
rect 9416 29306 9444 29514
rect 9404 29300 9456 29306
rect 9404 29242 9456 29248
rect 9312 28688 9364 28694
rect 9312 28630 9364 28636
rect 9404 27872 9456 27878
rect 9404 27814 9456 27820
rect 8944 26580 8996 26586
rect 8944 26522 8996 26528
rect 8404 22066 8524 22094
rect 8588 26206 8800 26234
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 8312 17338 8340 19110
rect 8404 18834 8432 22066
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 8496 18902 8524 20198
rect 8484 18896 8536 18902
rect 8484 18838 8536 18844
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8484 17060 8536 17066
rect 8484 17002 8536 17008
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8312 16658 8340 16934
rect 8496 16726 8524 17002
rect 8484 16720 8536 16726
rect 8484 16662 8536 16668
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 8208 16516 8260 16522
rect 8208 16458 8260 16464
rect 8300 15632 8352 15638
rect 8300 15574 8352 15580
rect 8312 15502 8340 15574
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8024 15088 8076 15094
rect 8024 15030 8076 15036
rect 8404 15026 8432 16594
rect 8496 16114 8524 16662
rect 8484 16108 8536 16114
rect 8484 16050 8536 16056
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8588 14482 8616 26206
rect 8668 25152 8720 25158
rect 8666 25120 8668 25129
rect 8720 25120 8722 25129
rect 8666 25055 8722 25064
rect 8668 23792 8720 23798
rect 8668 23734 8720 23740
rect 8680 15706 8708 23734
rect 8760 18760 8812 18766
rect 8760 18702 8812 18708
rect 8772 18358 8800 18702
rect 8852 18624 8904 18630
rect 8852 18566 8904 18572
rect 8760 18352 8812 18358
rect 8760 18294 8812 18300
rect 8760 17060 8812 17066
rect 8760 17002 8812 17008
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8772 15638 8800 17002
rect 8760 15632 8812 15638
rect 8760 15574 8812 15580
rect 8772 15026 8800 15574
rect 8864 15570 8892 18566
rect 8852 15564 8904 15570
rect 8852 15506 8904 15512
rect 8760 15020 8812 15026
rect 8760 14962 8812 14968
rect 8576 14476 8628 14482
rect 8576 14418 8628 14424
rect 8956 14414 8984 26522
rect 9128 25832 9180 25838
rect 9128 25774 9180 25780
rect 9140 25362 9168 25774
rect 9128 25356 9180 25362
rect 9128 25298 9180 25304
rect 9220 24132 9272 24138
rect 9220 24074 9272 24080
rect 9128 22568 9180 22574
rect 9128 22510 9180 22516
rect 9140 21486 9168 22510
rect 9128 21480 9180 21486
rect 9128 21422 9180 21428
rect 9140 21010 9168 21422
rect 9128 21004 9180 21010
rect 9128 20946 9180 20952
rect 9036 20936 9088 20942
rect 9036 20878 9088 20884
rect 9048 15706 9076 20878
rect 9140 20534 9168 20946
rect 9128 20528 9180 20534
rect 9128 20470 9180 20476
rect 9140 19378 9168 20470
rect 9128 19372 9180 19378
rect 9128 19314 9180 19320
rect 9232 17882 9260 24074
rect 9312 23112 9364 23118
rect 9312 23054 9364 23060
rect 9324 21962 9352 23054
rect 9312 21956 9364 21962
rect 9312 21898 9364 21904
rect 9324 19854 9352 21898
rect 9416 20330 9444 27814
rect 9404 20324 9456 20330
rect 9404 20266 9456 20272
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9324 18766 9352 19790
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9404 18692 9456 18698
rect 9404 18634 9456 18640
rect 9416 18426 9444 18634
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 9220 17876 9272 17882
rect 9220 17818 9272 17824
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9140 16998 9168 17614
rect 9220 17128 9272 17134
rect 9220 17070 9272 17076
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 9140 15502 9168 16934
rect 9232 16522 9260 17070
rect 9220 16516 9272 16522
rect 9220 16458 9272 16464
rect 9508 16250 9536 33458
rect 9600 32502 9628 33798
rect 9692 33114 9720 34002
rect 9680 33108 9732 33114
rect 9680 33050 9732 33056
rect 9588 32496 9640 32502
rect 9640 32444 9720 32450
rect 9588 32438 9720 32444
rect 9600 32422 9720 32438
rect 9692 32366 9720 32422
rect 9680 32360 9732 32366
rect 9680 32302 9732 32308
rect 9772 31136 9824 31142
rect 9772 31078 9824 31084
rect 9588 30796 9640 30802
rect 9588 30738 9640 30744
rect 9600 28218 9628 30738
rect 9680 30184 9732 30190
rect 9680 30126 9732 30132
rect 9588 28212 9640 28218
rect 9588 28154 9640 28160
rect 9692 28150 9720 30126
rect 9680 28144 9732 28150
rect 9680 28086 9732 28092
rect 9588 28008 9640 28014
rect 9588 27950 9640 27956
rect 9600 27606 9628 27950
rect 9588 27600 9640 27606
rect 9588 27542 9640 27548
rect 9692 27538 9720 28086
rect 9680 27532 9732 27538
rect 9680 27474 9732 27480
rect 9784 26234 9812 31078
rect 9968 26234 9996 37198
rect 10060 36553 10088 37198
rect 10980 37194 11100 37210
rect 12256 37198 12308 37204
rect 13556 37210 13584 39200
rect 14096 37256 14148 37262
rect 10876 37188 10928 37194
rect 10980 37188 11112 37194
rect 10980 37182 11060 37188
rect 10876 37130 10928 37136
rect 13556 37182 13860 37210
rect 14096 37198 14148 37204
rect 11060 37130 11112 37136
rect 10888 36718 10916 37130
rect 13832 37126 13860 37182
rect 12808 37120 12860 37126
rect 12808 37062 12860 37068
rect 13452 37120 13504 37126
rect 13452 37062 13504 37068
rect 13728 37120 13780 37126
rect 13728 37062 13780 37068
rect 13820 37120 13872 37126
rect 13820 37062 13872 37068
rect 12348 36780 12400 36786
rect 12348 36722 12400 36728
rect 10876 36712 10928 36718
rect 10876 36654 10928 36660
rect 10046 36544 10102 36553
rect 10046 36479 10102 36488
rect 12360 36378 12388 36722
rect 12716 36644 12768 36650
rect 12716 36586 12768 36592
rect 12728 36378 12756 36586
rect 12820 36417 12848 37062
rect 13358 36952 13414 36961
rect 13358 36887 13414 36896
rect 13464 36904 13492 37062
rect 13636 36916 13688 36922
rect 13372 36854 13400 36887
rect 13464 36876 13636 36904
rect 13636 36858 13688 36864
rect 13740 36854 13768 37062
rect 13360 36848 13412 36854
rect 13360 36790 13412 36796
rect 13728 36848 13780 36854
rect 13728 36790 13780 36796
rect 12992 36576 13044 36582
rect 12992 36518 13044 36524
rect 13636 36576 13688 36582
rect 13636 36518 13688 36524
rect 12806 36408 12862 36417
rect 12348 36372 12400 36378
rect 12348 36314 12400 36320
rect 12716 36372 12768 36378
rect 12806 36343 12862 36352
rect 12716 36314 12768 36320
rect 11704 36168 11756 36174
rect 11704 36110 11756 36116
rect 11610 35864 11666 35873
rect 11610 35799 11666 35808
rect 11336 35760 11388 35766
rect 11336 35702 11388 35708
rect 10508 35692 10560 35698
rect 10508 35634 10560 35640
rect 10520 35290 10548 35634
rect 10876 35624 10928 35630
rect 10876 35566 10928 35572
rect 10508 35284 10560 35290
rect 10508 35226 10560 35232
rect 10784 32904 10836 32910
rect 10784 32846 10836 32852
rect 10508 32564 10560 32570
rect 10508 32506 10560 32512
rect 10520 31822 10548 32506
rect 10796 31822 10824 32846
rect 10888 32842 10916 35566
rect 11152 35216 11204 35222
rect 11152 35158 11204 35164
rect 11058 34504 11114 34513
rect 11058 34439 11114 34448
rect 11072 33114 11100 34439
rect 11164 33862 11192 35158
rect 11348 34542 11376 35702
rect 11428 35692 11480 35698
rect 11428 35634 11480 35640
rect 11440 35601 11468 35634
rect 11426 35592 11482 35601
rect 11426 35527 11482 35536
rect 11624 35154 11652 35799
rect 11612 35148 11664 35154
rect 11612 35090 11664 35096
rect 11716 35086 11744 36110
rect 12440 35828 12492 35834
rect 12440 35770 12492 35776
rect 12452 35562 12480 35770
rect 13004 35737 13032 36518
rect 12990 35728 13046 35737
rect 12990 35663 13046 35672
rect 12440 35556 12492 35562
rect 12440 35498 12492 35504
rect 13452 35488 13504 35494
rect 13452 35430 13504 35436
rect 11704 35080 11756 35086
rect 11704 35022 11756 35028
rect 12070 35048 12126 35057
rect 11610 34640 11666 34649
rect 11610 34575 11666 34584
rect 11336 34536 11388 34542
rect 11336 34478 11388 34484
rect 11152 33856 11204 33862
rect 11152 33798 11204 33804
rect 11164 33590 11192 33798
rect 11152 33584 11204 33590
rect 11152 33526 11204 33532
rect 11624 33454 11652 34575
rect 11716 34542 11744 35022
rect 12070 34983 12126 34992
rect 12084 34950 12112 34983
rect 12072 34944 12124 34950
rect 12072 34886 12124 34892
rect 13360 34672 13412 34678
rect 13360 34614 13412 34620
rect 11704 34536 11756 34542
rect 11704 34478 11756 34484
rect 11716 34066 11744 34478
rect 11796 34400 11848 34406
rect 13372 34377 13400 34614
rect 11796 34342 11848 34348
rect 13358 34368 13414 34377
rect 11808 34218 11836 34342
rect 13358 34303 13414 34312
rect 12254 34232 12310 34241
rect 11808 34202 12204 34218
rect 11808 34196 12216 34202
rect 11808 34190 12164 34196
rect 12254 34167 12310 34176
rect 12164 34138 12216 34144
rect 11704 34060 11756 34066
rect 11704 34002 11756 34008
rect 11612 33448 11664 33454
rect 11612 33390 11664 33396
rect 11610 33144 11666 33153
rect 11060 33108 11112 33114
rect 11610 33079 11666 33088
rect 11060 33050 11112 33056
rect 10876 32836 10928 32842
rect 10876 32778 10928 32784
rect 11060 32224 11112 32230
rect 11060 32166 11112 32172
rect 10508 31816 10560 31822
rect 10508 31758 10560 31764
rect 10784 31816 10836 31822
rect 10784 31758 10836 31764
rect 10796 30802 10824 31758
rect 10784 30796 10836 30802
rect 10784 30738 10836 30744
rect 10784 30660 10836 30666
rect 10784 30602 10836 30608
rect 10692 28076 10744 28082
rect 10692 28018 10744 28024
rect 10704 27674 10732 28018
rect 10692 27668 10744 27674
rect 10692 27610 10744 27616
rect 9692 26206 9812 26234
rect 9876 26206 9996 26234
rect 9692 25158 9720 26206
rect 9680 25152 9732 25158
rect 9680 25094 9732 25100
rect 9588 24404 9640 24410
rect 9588 24346 9640 24352
rect 9600 24070 9628 24346
rect 9588 24064 9640 24070
rect 9588 24006 9640 24012
rect 9692 22658 9720 25094
rect 9772 24812 9824 24818
rect 9772 24754 9824 24760
rect 9784 24410 9812 24754
rect 9772 24404 9824 24410
rect 9772 24346 9824 24352
rect 9876 22794 9904 26206
rect 10508 25288 10560 25294
rect 10508 25230 10560 25236
rect 10140 24676 10192 24682
rect 10140 24618 10192 24624
rect 10152 23662 10180 24618
rect 10140 23656 10192 23662
rect 10140 23598 10192 23604
rect 9876 22766 10180 22794
rect 9692 22630 10088 22658
rect 9680 21956 9732 21962
rect 9680 21898 9732 21904
rect 9588 19780 9640 19786
rect 9588 19722 9640 19728
rect 9600 19514 9628 19722
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9588 16516 9640 16522
rect 9588 16458 9640 16464
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9404 16176 9456 16182
rect 9404 16118 9456 16124
rect 9310 15872 9366 15881
rect 9310 15807 9366 15816
rect 9324 15638 9352 15807
rect 9312 15632 9364 15638
rect 9312 15574 9364 15580
rect 9416 15570 9444 16118
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 9508 15978 9536 16050
rect 9496 15972 9548 15978
rect 9496 15914 9548 15920
rect 9600 15688 9628 16458
rect 9508 15660 9628 15688
rect 9404 15564 9456 15570
rect 9404 15506 9456 15512
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9404 14884 9456 14890
rect 9404 14826 9456 14832
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 7656 14272 7708 14278
rect 7656 14214 7708 14220
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7668 14006 7696 14214
rect 7656 14000 7708 14006
rect 7656 13942 7708 13948
rect 7852 13870 7880 14214
rect 9416 14006 9444 14826
rect 9508 14074 9536 15660
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9220 14000 9272 14006
rect 9220 13942 9272 13948
rect 9404 14000 9456 14006
rect 9404 13942 9456 13948
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 7196 12912 7248 12918
rect 7196 12854 7248 12860
rect 7208 12442 7236 12854
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7852 11830 7880 13806
rect 8114 13696 8170 13705
rect 8114 13631 8170 13640
rect 8128 13326 8156 13631
rect 9140 13462 9168 13806
rect 9232 13530 9260 13942
rect 9416 13870 9444 13942
rect 9404 13864 9456 13870
rect 9404 13806 9456 13812
rect 9494 13696 9550 13705
rect 9494 13631 9550 13640
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 8300 13456 8352 13462
rect 8300 13398 8352 13404
rect 9128 13456 9180 13462
rect 9128 13398 9180 13404
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8312 12782 8340 13398
rect 9508 13326 9536 13631
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7944 11898 7972 12038
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 8206 11792 8262 11801
rect 8206 11727 8262 11736
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 7944 11082 7972 11562
rect 8220 11218 8248 11727
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8588 11150 8616 12378
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 6828 10736 6880 10742
rect 6828 10678 6880 10684
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 5724 7472 5776 7478
rect 5724 7414 5776 7420
rect 5736 4146 5764 7414
rect 6564 5370 6592 10610
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6656 4622 6684 6598
rect 6748 6322 6776 7142
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 6748 3058 6776 3878
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 2780 2984 2832 2990
rect 2780 2926 2832 2932
rect 1952 2304 2004 2310
rect 1952 2246 2004 2252
rect 1674 2136 1730 2145
rect 1674 2071 1730 2080
rect 1964 800 1992 2246
rect 18 200 74 800
rect 662 200 718 800
rect 1950 200 2006 800
rect 2792 785 2820 2926
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 6564 2446 6592 2790
rect 7300 2650 7328 9998
rect 7944 9518 7972 11018
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 9324 2514 9352 13126
rect 9600 9110 9628 15506
rect 9692 15094 9720 21898
rect 9772 21344 9824 21350
rect 9772 21286 9824 21292
rect 9784 19446 9812 21286
rect 9772 19440 9824 19446
rect 9772 19382 9824 19388
rect 9956 19440 10008 19446
rect 9956 19382 10008 19388
rect 9784 17354 9812 19382
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9876 17542 9904 18634
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9784 17326 9904 17354
rect 9770 15192 9826 15201
rect 9770 15127 9826 15136
rect 9680 15088 9732 15094
rect 9680 15030 9732 15036
rect 9784 15026 9812 15127
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 9784 13841 9812 13942
rect 9770 13832 9826 13841
rect 9770 13767 9826 13776
rect 9772 11824 9824 11830
rect 9772 11766 9824 11772
rect 9784 11558 9812 11766
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9876 11150 9904 17326
rect 9968 14890 9996 19382
rect 10060 17728 10088 22630
rect 10152 21690 10180 22766
rect 10140 21684 10192 21690
rect 10140 21626 10192 21632
rect 10416 20868 10468 20874
rect 10416 20810 10468 20816
rect 10140 19304 10192 19310
rect 10140 19246 10192 19252
rect 10152 18204 10180 19246
rect 10324 18964 10376 18970
rect 10324 18906 10376 18912
rect 10336 18358 10364 18906
rect 10324 18352 10376 18358
rect 10324 18294 10376 18300
rect 10152 18176 10272 18204
rect 10060 17700 10180 17728
rect 9956 14884 10008 14890
rect 9956 14826 10008 14832
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 10060 14346 10088 14758
rect 10048 14340 10100 14346
rect 10048 14282 10100 14288
rect 10152 13326 10180 17700
rect 10244 15994 10272 18176
rect 10428 17882 10456 20810
rect 10416 17876 10468 17882
rect 10416 17818 10468 17824
rect 10416 17264 10468 17270
rect 10416 17206 10468 17212
rect 10324 16584 10376 16590
rect 10324 16526 10376 16532
rect 10336 16114 10364 16526
rect 10428 16114 10456 17206
rect 10520 16250 10548 25230
rect 10600 24608 10652 24614
rect 10600 24550 10652 24556
rect 10612 16454 10640 24550
rect 10796 24070 10824 30602
rect 11072 29102 11100 32166
rect 11624 31754 11652 33079
rect 11716 32366 11744 34002
rect 12268 33930 12296 34167
rect 13268 33992 13320 33998
rect 13268 33934 13320 33940
rect 12256 33924 12308 33930
rect 12256 33866 12308 33872
rect 11886 33824 11942 33833
rect 11886 33759 11942 33768
rect 11900 33386 11928 33759
rect 12622 33688 12678 33697
rect 13280 33658 13308 33934
rect 12622 33623 12678 33632
rect 13268 33652 13320 33658
rect 11980 33516 12032 33522
rect 11980 33458 12032 33464
rect 11888 33380 11940 33386
rect 11888 33322 11940 33328
rect 11992 32774 12020 33458
rect 12348 33448 12400 33454
rect 12348 33390 12400 33396
rect 12164 33312 12216 33318
rect 12164 33254 12216 33260
rect 12176 33096 12204 33254
rect 12256 33108 12308 33114
rect 12176 33068 12256 33096
rect 12256 33050 12308 33056
rect 11888 32768 11940 32774
rect 11888 32710 11940 32716
rect 11980 32768 12032 32774
rect 11980 32710 12032 32716
rect 11900 32473 11928 32710
rect 11992 32502 12020 32710
rect 11980 32496 12032 32502
rect 11886 32464 11942 32473
rect 11980 32438 12032 32444
rect 11886 32399 11942 32408
rect 11704 32360 11756 32366
rect 11704 32302 11756 32308
rect 11888 32360 11940 32366
rect 11888 32302 11940 32308
rect 11796 31884 11848 31890
rect 11796 31826 11848 31832
rect 11612 31748 11664 31754
rect 11612 31690 11664 31696
rect 11624 31278 11652 31690
rect 11704 31340 11756 31346
rect 11704 31282 11756 31288
rect 11152 31272 11204 31278
rect 11152 31214 11204 31220
rect 11612 31272 11664 31278
rect 11612 31214 11664 31220
rect 11060 29096 11112 29102
rect 11060 29038 11112 29044
rect 10968 28960 11020 28966
rect 11020 28908 11100 28914
rect 10968 28902 11100 28908
rect 10980 28886 11100 28902
rect 10968 25832 11020 25838
rect 10968 25774 11020 25780
rect 10876 25764 10928 25770
rect 10876 25706 10928 25712
rect 10888 25498 10916 25706
rect 10876 25492 10928 25498
rect 10876 25434 10928 25440
rect 10784 24064 10836 24070
rect 10784 24006 10836 24012
rect 10784 22092 10836 22098
rect 10784 22034 10836 22040
rect 10692 20596 10744 20602
rect 10692 20538 10744 20544
rect 10704 19854 10732 20538
rect 10692 19848 10744 19854
rect 10692 19790 10744 19796
rect 10796 17202 10824 22034
rect 10980 19786 11008 25774
rect 11072 25702 11100 28886
rect 11060 25696 11112 25702
rect 11060 25638 11112 25644
rect 11072 22953 11100 25638
rect 11058 22944 11114 22953
rect 11058 22879 11114 22888
rect 11060 22772 11112 22778
rect 11060 22714 11112 22720
rect 10968 19780 11020 19786
rect 10968 19722 11020 19728
rect 11072 19718 11100 22714
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 11072 19446 11100 19654
rect 11060 19440 11112 19446
rect 11060 19382 11112 19388
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 10784 17196 10836 17202
rect 10784 17138 10836 17144
rect 10600 16448 10652 16454
rect 10600 16390 10652 16396
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10980 16250 11008 16390
rect 10508 16244 10560 16250
rect 10508 16186 10560 16192
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 11072 16182 11100 19246
rect 11164 16182 11192 31214
rect 11336 30320 11388 30326
rect 11336 30262 11388 30268
rect 11348 29646 11376 30262
rect 11716 30190 11744 31282
rect 11704 30184 11756 30190
rect 11704 30126 11756 30132
rect 11336 29640 11388 29646
rect 11336 29582 11388 29588
rect 11348 27062 11376 29582
rect 11520 29504 11572 29510
rect 11520 29446 11572 29452
rect 11532 29238 11560 29446
rect 11520 29232 11572 29238
rect 11520 29174 11572 29180
rect 11612 29164 11664 29170
rect 11612 29106 11664 29112
rect 11428 29096 11480 29102
rect 11428 29038 11480 29044
rect 11336 27056 11388 27062
rect 11336 26998 11388 27004
rect 11348 24750 11376 26998
rect 11440 25809 11468 29038
rect 11624 28626 11652 29106
rect 11612 28620 11664 28626
rect 11612 28562 11664 28568
rect 11808 27538 11836 31826
rect 11900 31822 11928 32302
rect 11888 31816 11940 31822
rect 11888 31758 11940 31764
rect 11992 30326 12020 32438
rect 12360 32366 12388 33390
rect 12636 32842 12664 33623
rect 13268 33594 13320 33600
rect 13084 33584 13136 33590
rect 13136 33544 13216 33572
rect 13084 33526 13136 33532
rect 12624 32836 12676 32842
rect 12624 32778 12676 32784
rect 12992 32836 13044 32842
rect 12992 32778 13044 32784
rect 13004 32745 13032 32778
rect 12990 32736 13046 32745
rect 12990 32671 13046 32680
rect 12348 32360 12400 32366
rect 12348 32302 12400 32308
rect 12254 31920 12310 31929
rect 12254 31855 12310 31864
rect 12268 31754 12296 31855
rect 12256 31748 12308 31754
rect 12256 31690 12308 31696
rect 12072 31408 12124 31414
rect 12072 31350 12124 31356
rect 12084 31278 12112 31350
rect 12072 31272 12124 31278
rect 12072 31214 12124 31220
rect 13004 30938 13032 32671
rect 12992 30932 13044 30938
rect 12992 30874 13044 30880
rect 11980 30320 12032 30326
rect 11980 30262 12032 30268
rect 11992 30054 12020 30262
rect 12348 30252 12400 30258
rect 12348 30194 12400 30200
rect 12072 30184 12124 30190
rect 12072 30126 12124 30132
rect 11980 30048 12032 30054
rect 11980 29990 12032 29996
rect 12084 29578 12112 30126
rect 12072 29572 12124 29578
rect 12072 29514 12124 29520
rect 12084 29238 12112 29514
rect 12072 29232 12124 29238
rect 12072 29174 12124 29180
rect 12360 29073 12388 30194
rect 12346 29064 12402 29073
rect 12346 28999 12402 29008
rect 13188 28994 13216 33544
rect 13464 33046 13492 35430
rect 13648 35193 13676 36518
rect 14002 36272 14058 36281
rect 14002 36207 14058 36216
rect 13728 36100 13780 36106
rect 13728 36042 13780 36048
rect 13740 35834 13768 36042
rect 13912 36032 13964 36038
rect 13912 35974 13964 35980
rect 13728 35828 13780 35834
rect 13728 35770 13780 35776
rect 13634 35184 13690 35193
rect 13634 35119 13690 35128
rect 13544 35012 13596 35018
rect 13544 34954 13596 34960
rect 13636 35012 13688 35018
rect 13636 34954 13688 34960
rect 13556 34746 13584 34954
rect 13544 34740 13596 34746
rect 13544 34682 13596 34688
rect 13452 33040 13504 33046
rect 13452 32982 13504 32988
rect 13648 31686 13676 34954
rect 13740 34678 13768 35770
rect 13924 35698 13952 35974
rect 14016 35834 14044 36207
rect 14108 36038 14136 37198
rect 14200 36938 14228 39200
rect 15488 37262 15516 39200
rect 15200 37256 15252 37262
rect 15200 37198 15252 37204
rect 15476 37256 15528 37262
rect 15476 37198 15528 37204
rect 14200 36910 14320 36938
rect 14188 36780 14240 36786
rect 14188 36722 14240 36728
rect 14096 36032 14148 36038
rect 14096 35974 14148 35980
rect 14004 35828 14056 35834
rect 14004 35770 14056 35776
rect 13912 35692 13964 35698
rect 13912 35634 13964 35640
rect 14096 35624 14148 35630
rect 14096 35566 14148 35572
rect 13728 34672 13780 34678
rect 13728 34614 13780 34620
rect 13912 34536 13964 34542
rect 13912 34478 13964 34484
rect 13728 34196 13780 34202
rect 13728 34138 13780 34144
rect 13740 33017 13768 34138
rect 13726 33008 13782 33017
rect 13726 32943 13782 32952
rect 13820 32428 13872 32434
rect 13820 32370 13872 32376
rect 13832 32026 13860 32370
rect 13820 32020 13872 32026
rect 13820 31962 13872 31968
rect 13924 31929 13952 34478
rect 13910 31920 13966 31929
rect 13820 31884 13872 31890
rect 13910 31855 13966 31864
rect 13820 31826 13872 31832
rect 13636 31680 13688 31686
rect 13636 31622 13688 31628
rect 13728 31680 13780 31686
rect 13728 31622 13780 31628
rect 13648 30977 13676 31622
rect 13634 30968 13690 30977
rect 13634 30903 13690 30912
rect 13544 29708 13596 29714
rect 13544 29650 13596 29656
rect 13452 29572 13504 29578
rect 13452 29514 13504 29520
rect 13096 28966 13216 28994
rect 12072 28960 12124 28966
rect 12072 28902 12124 28908
rect 11888 28484 11940 28490
rect 11888 28426 11940 28432
rect 11796 27532 11848 27538
rect 11796 27474 11848 27480
rect 11612 26920 11664 26926
rect 11612 26862 11664 26868
rect 11624 26382 11652 26862
rect 11612 26376 11664 26382
rect 11612 26318 11664 26324
rect 11704 26376 11756 26382
rect 11704 26318 11756 26324
rect 11716 25838 11744 26318
rect 11704 25832 11756 25838
rect 11426 25800 11482 25809
rect 11756 25792 11836 25820
rect 11704 25774 11756 25780
rect 11426 25735 11482 25744
rect 11808 25294 11836 25792
rect 11796 25288 11848 25294
rect 11796 25230 11848 25236
rect 11808 24750 11836 25230
rect 11336 24744 11388 24750
rect 11336 24686 11388 24692
rect 11796 24744 11848 24750
rect 11796 24686 11848 24692
rect 11348 23798 11376 24686
rect 11704 24336 11756 24342
rect 11704 24278 11756 24284
rect 11336 23792 11388 23798
rect 11336 23734 11388 23740
rect 11428 22432 11480 22438
rect 11428 22374 11480 22380
rect 11520 22432 11572 22438
rect 11520 22374 11572 22380
rect 11440 22114 11468 22374
rect 11532 22234 11560 22374
rect 11520 22228 11572 22234
rect 11520 22170 11572 22176
rect 11440 22086 11652 22114
rect 11520 19508 11572 19514
rect 11520 19450 11572 19456
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11348 18426 11376 18566
rect 11336 18420 11388 18426
rect 11336 18362 11388 18368
rect 11348 18222 11376 18362
rect 11336 18216 11388 18222
rect 11336 18158 11388 18164
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 11152 16176 11204 16182
rect 11152 16118 11204 16124
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10416 16108 10468 16114
rect 10416 16050 10468 16056
rect 10600 16040 10652 16046
rect 10414 16008 10470 16017
rect 10244 15966 10364 15994
rect 10232 15904 10284 15910
rect 10232 15846 10284 15852
rect 10244 15638 10272 15846
rect 10232 15632 10284 15638
rect 10232 15574 10284 15580
rect 10232 14884 10284 14890
rect 10232 14826 10284 14832
rect 10244 14482 10272 14826
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10336 12170 10364 15966
rect 10600 15982 10652 15988
rect 10414 15943 10470 15952
rect 10428 15502 10456 15943
rect 10612 15706 10640 15982
rect 10600 15700 10652 15706
rect 10520 15660 10600 15688
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10520 13870 10548 15660
rect 10600 15642 10652 15648
rect 11532 15314 11560 19450
rect 11624 15502 11652 22086
rect 11716 19514 11744 24278
rect 11808 23866 11836 24686
rect 11796 23860 11848 23866
rect 11796 23802 11848 23808
rect 11808 22098 11836 23802
rect 11900 22506 11928 28426
rect 12084 26790 12112 28902
rect 13096 28762 13124 28966
rect 13084 28756 13136 28762
rect 13084 28698 13136 28704
rect 12348 27532 12400 27538
rect 12348 27474 12400 27480
rect 12360 27402 12388 27474
rect 12348 27396 12400 27402
rect 12348 27338 12400 27344
rect 13176 27328 13228 27334
rect 13176 27270 13228 27276
rect 12072 26784 12124 26790
rect 12072 26726 12124 26732
rect 11888 22500 11940 22506
rect 11888 22442 11940 22448
rect 11796 22092 11848 22098
rect 11796 22034 11848 22040
rect 11796 21888 11848 21894
rect 11796 21830 11848 21836
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 11808 16658 11836 21830
rect 11980 20392 12032 20398
rect 11980 20334 12032 20340
rect 11992 19922 12020 20334
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 11992 18834 12020 19858
rect 11980 18828 12032 18834
rect 11980 18770 12032 18776
rect 11980 17264 12032 17270
rect 11980 17206 12032 17212
rect 11992 17066 12020 17206
rect 11888 17060 11940 17066
rect 11888 17002 11940 17008
rect 11980 17060 12032 17066
rect 11980 17002 12032 17008
rect 11900 16658 11928 17002
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11980 15360 12032 15366
rect 11532 15286 11652 15314
rect 11980 15302 12032 15308
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 11060 14340 11112 14346
rect 11060 14282 11112 14288
rect 10600 14000 10652 14006
rect 10600 13942 10652 13948
rect 10508 13864 10560 13870
rect 10508 13806 10560 13812
rect 10612 12374 10640 13942
rect 11072 12918 11100 14282
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 10600 12368 10652 12374
rect 10600 12310 10652 12316
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10336 6798 10364 7686
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9312 2508 9364 2514
rect 9312 2450 9364 2456
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 3252 800 3280 2246
rect 3896 800 3924 2382
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 5184 800 5212 2246
rect 5276 2106 5304 2382
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 5264 2100 5316 2106
rect 5264 2042 5316 2048
rect 6472 800 6500 2246
rect 7116 800 7144 2382
rect 8404 800 8432 2382
rect 9692 800 9720 2994
rect 10428 2582 10456 11494
rect 10520 11354 10548 11630
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 10704 11218 10732 11630
rect 11164 11626 11192 14418
rect 11532 13870 11560 14758
rect 11244 13864 11296 13870
rect 11242 13832 11244 13841
rect 11520 13864 11572 13870
rect 11296 13832 11298 13841
rect 11520 13806 11572 13812
rect 11242 13767 11298 13776
rect 11532 12306 11560 13806
rect 11624 12434 11652 15286
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 11716 14793 11744 14894
rect 11702 14784 11758 14793
rect 11702 14719 11758 14728
rect 11900 14618 11928 14894
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 11992 14346 12020 15302
rect 12084 14958 12112 26726
rect 12256 26308 12308 26314
rect 12256 26250 12308 26256
rect 12268 22982 12296 26250
rect 12992 26240 13044 26246
rect 12992 26182 13044 26188
rect 13004 25786 13032 26182
rect 13004 25758 13124 25786
rect 12992 24676 13044 24682
rect 12992 24618 13044 24624
rect 13004 24342 13032 24618
rect 12992 24336 13044 24342
rect 12992 24278 13044 24284
rect 12992 23248 13044 23254
rect 12992 23190 13044 23196
rect 12348 23112 12400 23118
rect 12808 23112 12860 23118
rect 12348 23054 12400 23060
rect 12806 23080 12808 23089
rect 12900 23112 12952 23118
rect 12860 23080 12862 23089
rect 12256 22976 12308 22982
rect 12256 22918 12308 22924
rect 12360 22094 12388 23054
rect 12716 23044 12768 23050
rect 12900 23054 12952 23060
rect 12806 23015 12862 23024
rect 12716 22986 12768 22992
rect 12268 22066 12388 22094
rect 12164 20800 12216 20806
rect 12164 20742 12216 20748
rect 12176 19786 12204 20742
rect 12164 19780 12216 19786
rect 12164 19722 12216 19728
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 12070 14784 12126 14793
rect 12070 14719 12126 14728
rect 12084 14618 12112 14719
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 11980 14340 12032 14346
rect 11980 14282 12032 14288
rect 11888 14000 11940 14006
rect 11888 13942 11940 13948
rect 11900 13530 11928 13942
rect 12084 13870 12112 14418
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11624 12406 11744 12434
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11716 12238 11744 12406
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11152 11620 11204 11626
rect 11152 11562 11204 11568
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10508 11144 10560 11150
rect 10888 11098 10916 11494
rect 11164 11218 11192 11562
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 10560 11092 10916 11098
rect 10508 11086 10916 11092
rect 10520 11070 10916 11086
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10980 7410 11008 8978
rect 11348 8906 11376 12038
rect 11980 11824 12032 11830
rect 11980 11766 12032 11772
rect 11612 11620 11664 11626
rect 11612 11562 11664 11568
rect 11624 11218 11652 11562
rect 11992 11354 12020 11766
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 11244 8900 11296 8906
rect 11244 8842 11296 8848
rect 11336 8900 11388 8906
rect 11336 8842 11388 8848
rect 11152 8424 11204 8430
rect 11152 8366 11204 8372
rect 11164 7410 11192 8366
rect 11256 8022 11284 8842
rect 11244 8016 11296 8022
rect 11244 7958 11296 7964
rect 11900 7478 11928 10406
rect 12176 8498 12204 19722
rect 12268 19378 12296 22066
rect 12624 21956 12676 21962
rect 12624 21898 12676 21904
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 12348 19440 12400 19446
rect 12348 19382 12400 19388
rect 12256 19372 12308 19378
rect 12256 19314 12308 19320
rect 12360 13462 12388 19382
rect 12452 15706 12480 21082
rect 12532 17604 12584 17610
rect 12532 17546 12584 17552
rect 12544 16590 12572 17546
rect 12532 16584 12584 16590
rect 12532 16526 12584 16532
rect 12636 16250 12664 21898
rect 12624 16244 12676 16250
rect 12624 16186 12676 16192
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12440 14544 12492 14550
rect 12440 14486 12492 14492
rect 12452 14278 12480 14486
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12348 13456 12400 13462
rect 12348 13398 12400 13404
rect 12728 13326 12756 22986
rect 12912 22234 12940 23054
rect 12900 22228 12952 22234
rect 12900 22170 12952 22176
rect 12808 18352 12860 18358
rect 12808 18294 12860 18300
rect 12820 15570 12848 18294
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 12912 17746 12940 18158
rect 12900 17740 12952 17746
rect 12900 17682 12952 17688
rect 13004 17542 13032 23190
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12912 14346 12940 14894
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 13004 11150 13032 17478
rect 13096 16153 13124 25758
rect 13188 24818 13216 27270
rect 13268 26512 13320 26518
rect 13268 26454 13320 26460
rect 13176 24812 13228 24818
rect 13176 24754 13228 24760
rect 13280 24698 13308 26454
rect 13464 25838 13492 29514
rect 13556 29306 13584 29650
rect 13544 29300 13596 29306
rect 13544 29242 13596 29248
rect 13636 28688 13688 28694
rect 13636 28630 13688 28636
rect 13648 27713 13676 28630
rect 13740 27878 13768 31622
rect 13832 30938 13860 31826
rect 13820 30932 13872 30938
rect 13820 30874 13872 30880
rect 13910 30832 13966 30841
rect 13910 30767 13966 30776
rect 13924 29646 13952 30767
rect 13912 29640 13964 29646
rect 13912 29582 13964 29588
rect 14108 28937 14136 35566
rect 14200 31686 14228 36722
rect 14292 35086 14320 36910
rect 15212 36786 15240 37198
rect 16776 37126 16804 39200
rect 17224 37664 17276 37670
rect 17224 37606 17276 37612
rect 17236 37398 17264 37606
rect 17224 37392 17276 37398
rect 17224 37334 17276 37340
rect 17316 37392 17368 37398
rect 17316 37334 17368 37340
rect 17328 37262 17356 37334
rect 16856 37256 16908 37262
rect 16856 37198 16908 37204
rect 17316 37256 17368 37262
rect 17316 37198 17368 37204
rect 15292 37120 15344 37126
rect 15292 37062 15344 37068
rect 16764 37120 16816 37126
rect 16764 37062 16816 37068
rect 15200 36780 15252 36786
rect 15200 36722 15252 36728
rect 14556 36712 14608 36718
rect 14556 36654 14608 36660
rect 14464 36644 14516 36650
rect 14464 36586 14516 36592
rect 14476 36242 14504 36586
rect 14464 36236 14516 36242
rect 14464 36178 14516 36184
rect 14372 36168 14424 36174
rect 14372 36110 14424 36116
rect 14280 35080 14332 35086
rect 14280 35022 14332 35028
rect 14384 34406 14412 36110
rect 14464 35556 14516 35562
rect 14464 35498 14516 35504
rect 14476 34950 14504 35498
rect 14464 34944 14516 34950
rect 14464 34886 14516 34892
rect 14372 34400 14424 34406
rect 14372 34342 14424 34348
rect 14464 32428 14516 32434
rect 14464 32370 14516 32376
rect 14370 32328 14426 32337
rect 14370 32263 14426 32272
rect 14384 32230 14412 32263
rect 14476 32230 14504 32370
rect 14372 32224 14424 32230
rect 14372 32166 14424 32172
rect 14464 32224 14516 32230
rect 14464 32166 14516 32172
rect 14568 31890 14596 36654
rect 14832 36576 14884 36582
rect 14832 36518 14884 36524
rect 14924 36576 14976 36582
rect 14924 36518 14976 36524
rect 14844 36378 14872 36518
rect 14740 36372 14792 36378
rect 14740 36314 14792 36320
rect 14832 36372 14884 36378
rect 14832 36314 14884 36320
rect 14752 35601 14780 36314
rect 14832 35624 14884 35630
rect 14738 35592 14794 35601
rect 14832 35566 14884 35572
rect 14738 35527 14794 35536
rect 14740 33108 14792 33114
rect 14740 33050 14792 33056
rect 14752 32502 14780 33050
rect 14740 32496 14792 32502
rect 14660 32456 14740 32484
rect 14556 31884 14608 31890
rect 14556 31826 14608 31832
rect 14188 31680 14240 31686
rect 14188 31622 14240 31628
rect 14556 30048 14608 30054
rect 14556 29990 14608 29996
rect 14464 29640 14516 29646
rect 14464 29582 14516 29588
rect 14476 29034 14504 29582
rect 14568 29481 14596 29990
rect 14554 29472 14610 29481
rect 14554 29407 14610 29416
rect 14464 29028 14516 29034
rect 14464 28970 14516 28976
rect 14094 28928 14150 28937
rect 14094 28863 14150 28872
rect 13728 27872 13780 27878
rect 13728 27814 13780 27820
rect 13634 27704 13690 27713
rect 13634 27639 13690 27648
rect 13728 27056 13780 27062
rect 13728 26998 13780 27004
rect 13452 25832 13504 25838
rect 13452 25774 13504 25780
rect 13188 24670 13308 24698
rect 13188 22438 13216 24670
rect 13268 22500 13320 22506
rect 13268 22442 13320 22448
rect 13176 22432 13228 22438
rect 13176 22374 13228 22380
rect 13188 22166 13216 22374
rect 13280 22234 13308 22442
rect 13268 22228 13320 22234
rect 13268 22170 13320 22176
rect 13176 22160 13228 22166
rect 13176 22102 13228 22108
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 13188 18222 13216 18566
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 13082 16144 13138 16153
rect 13082 16079 13138 16088
rect 13084 15360 13136 15366
rect 13084 15302 13136 15308
rect 13096 14414 13124 15302
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 13004 10742 13032 11086
rect 12992 10736 13044 10742
rect 12992 10678 13044 10684
rect 13188 10198 13216 18158
rect 13360 17536 13412 17542
rect 13360 17478 13412 17484
rect 13372 16726 13400 17478
rect 13360 16720 13412 16726
rect 13360 16662 13412 16668
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13176 10192 13228 10198
rect 13176 10134 13228 10140
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12164 8016 12216 8022
rect 12164 7958 12216 7964
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11716 6798 11744 7142
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11808 6458 11836 7278
rect 12084 7002 12112 7822
rect 12176 7342 12204 7958
rect 12452 7954 12480 8230
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12912 7410 12940 7686
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 13084 7336 13136 7342
rect 13084 7278 13136 7284
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 12360 2582 12388 6734
rect 13096 6458 13124 7278
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 12992 6316 13044 6322
rect 12992 6258 13044 6264
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 12544 2650 12572 5646
rect 13004 2650 13032 6258
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 13280 2582 13308 14214
rect 13464 12374 13492 25774
rect 13740 25498 13768 26998
rect 14660 25974 14688 32456
rect 14740 32438 14792 32444
rect 14740 31884 14792 31890
rect 14740 31826 14792 31832
rect 14752 31346 14780 31826
rect 14844 31414 14872 35566
rect 14936 34066 14964 36518
rect 15212 36174 15240 36722
rect 15016 36168 15068 36174
rect 15014 36136 15016 36145
rect 15200 36168 15252 36174
rect 15068 36136 15070 36145
rect 15200 36110 15252 36116
rect 15014 36071 15070 36080
rect 15200 36032 15252 36038
rect 15200 35974 15252 35980
rect 15212 35834 15240 35974
rect 15200 35828 15252 35834
rect 15200 35770 15252 35776
rect 15108 35760 15160 35766
rect 15304 35714 15332 37062
rect 15384 36848 15436 36854
rect 15382 36816 15384 36825
rect 15436 36816 15438 36825
rect 15382 36751 15438 36760
rect 16764 36780 16816 36786
rect 16868 36768 16896 37198
rect 17420 37126 17448 39200
rect 17500 37256 17552 37262
rect 17500 37198 17552 37204
rect 18604 37256 18656 37262
rect 18604 37198 18656 37204
rect 16948 37120 17000 37126
rect 16948 37062 17000 37068
rect 17408 37120 17460 37126
rect 17408 37062 17460 37068
rect 16816 36740 16896 36768
rect 16764 36722 16816 36728
rect 16488 36712 16540 36718
rect 16488 36654 16540 36660
rect 16212 36576 16264 36582
rect 16212 36518 16264 36524
rect 16028 36100 16080 36106
rect 16028 36042 16080 36048
rect 16120 36100 16172 36106
rect 16120 36042 16172 36048
rect 15384 36032 15436 36038
rect 15384 35974 15436 35980
rect 15160 35708 15332 35714
rect 15108 35702 15332 35708
rect 15120 35686 15332 35702
rect 15200 35624 15252 35630
rect 15028 35572 15200 35578
rect 15028 35566 15252 35572
rect 15028 35550 15240 35566
rect 15028 35222 15056 35550
rect 15200 35488 15252 35494
rect 15200 35430 15252 35436
rect 15016 35216 15068 35222
rect 15016 35158 15068 35164
rect 15212 35154 15240 35430
rect 15200 35148 15252 35154
rect 15200 35090 15252 35096
rect 15212 34066 15240 35090
rect 15290 34232 15346 34241
rect 15290 34167 15292 34176
rect 15344 34167 15346 34176
rect 15292 34138 15344 34144
rect 14924 34060 14976 34066
rect 14924 34002 14976 34008
rect 15200 34060 15252 34066
rect 15200 34002 15252 34008
rect 15212 33522 15240 34002
rect 15292 33856 15344 33862
rect 15292 33798 15344 33804
rect 15200 33516 15252 33522
rect 15200 33458 15252 33464
rect 14924 33040 14976 33046
rect 14924 32982 14976 32988
rect 14936 32881 14964 32982
rect 15212 32978 15240 33458
rect 15200 32972 15252 32978
rect 15200 32914 15252 32920
rect 14922 32872 14978 32881
rect 15304 32842 15332 33798
rect 14922 32807 14978 32816
rect 15292 32836 15344 32842
rect 15292 32778 15344 32784
rect 15396 32026 15424 35974
rect 15934 35320 15990 35329
rect 15934 35255 15990 35264
rect 15948 35018 15976 35255
rect 15936 35012 15988 35018
rect 15936 34954 15988 34960
rect 15474 34912 15530 34921
rect 15474 34847 15530 34856
rect 15488 32337 15516 34847
rect 16040 34785 16068 36042
rect 16132 35170 16160 36042
rect 16224 36009 16252 36518
rect 16500 36242 16528 36654
rect 16488 36236 16540 36242
rect 16488 36178 16540 36184
rect 16764 36236 16816 36242
rect 16764 36178 16816 36184
rect 16210 36000 16266 36009
rect 16210 35935 16266 35944
rect 16304 35760 16356 35766
rect 16304 35702 16356 35708
rect 16316 35562 16344 35702
rect 16500 35698 16528 36178
rect 16488 35692 16540 35698
rect 16488 35634 16540 35640
rect 16304 35556 16356 35562
rect 16304 35498 16356 35504
rect 16132 35142 16252 35170
rect 16500 35154 16528 35634
rect 16672 35488 16724 35494
rect 16672 35430 16724 35436
rect 16684 35154 16712 35430
rect 16120 35012 16172 35018
rect 16120 34954 16172 34960
rect 16132 34921 16160 34954
rect 16118 34912 16174 34921
rect 16118 34847 16174 34856
rect 16026 34776 16082 34785
rect 16026 34711 16082 34720
rect 15568 34604 15620 34610
rect 15568 34546 15620 34552
rect 15580 34241 15608 34546
rect 15566 34232 15622 34241
rect 15566 34167 15622 34176
rect 15844 33924 15896 33930
rect 15844 33866 15896 33872
rect 15856 33454 15884 33866
rect 15844 33448 15896 33454
rect 15842 33416 15844 33425
rect 15896 33416 15898 33425
rect 15842 33351 15898 33360
rect 15856 33325 15884 33351
rect 15566 33280 15622 33289
rect 15566 33215 15622 33224
rect 15474 32328 15530 32337
rect 15474 32263 15530 32272
rect 15384 32020 15436 32026
rect 15384 31962 15436 31968
rect 14924 31680 14976 31686
rect 14924 31622 14976 31628
rect 14936 31414 14964 31622
rect 14832 31408 14884 31414
rect 14832 31350 14884 31356
rect 14924 31408 14976 31414
rect 14924 31350 14976 31356
rect 14740 31340 14792 31346
rect 14740 31282 14792 31288
rect 15580 30870 15608 33215
rect 15844 32224 15896 32230
rect 15844 32166 15896 32172
rect 15568 30864 15620 30870
rect 15568 30806 15620 30812
rect 15856 30802 15884 32166
rect 15936 32020 15988 32026
rect 15936 31962 15988 31968
rect 15948 31754 15976 31962
rect 16040 31754 16068 34711
rect 16224 33289 16252 35142
rect 16488 35148 16540 35154
rect 16488 35090 16540 35096
rect 16672 35148 16724 35154
rect 16672 35090 16724 35096
rect 16580 34128 16632 34134
rect 16580 34070 16632 34076
rect 16592 33862 16620 34070
rect 16580 33856 16632 33862
rect 16580 33798 16632 33804
rect 16488 33516 16540 33522
rect 16488 33458 16540 33464
rect 16210 33280 16266 33289
rect 16210 33215 16266 33224
rect 16212 32972 16264 32978
rect 16212 32914 16264 32920
rect 16224 32366 16252 32914
rect 16396 32836 16448 32842
rect 16396 32778 16448 32784
rect 16212 32360 16264 32366
rect 16212 32302 16264 32308
rect 16304 32360 16356 32366
rect 16304 32302 16356 32308
rect 16212 32224 16264 32230
rect 16212 32166 16264 32172
rect 15936 31748 15988 31754
rect 16040 31726 16160 31754
rect 15936 31690 15988 31696
rect 15844 30796 15896 30802
rect 15844 30738 15896 30744
rect 15108 30592 15160 30598
rect 15108 30534 15160 30540
rect 14740 28960 14792 28966
rect 14740 28902 14792 28908
rect 14752 28801 14780 28902
rect 14738 28792 14794 28801
rect 14738 28727 14794 28736
rect 15014 27568 15070 27577
rect 15014 27503 15070 27512
rect 15028 26353 15056 27503
rect 15014 26344 15070 26353
rect 15014 26279 15070 26288
rect 14648 25968 14700 25974
rect 14648 25910 14700 25916
rect 14832 25900 14884 25906
rect 14832 25842 14884 25848
rect 13728 25492 13780 25498
rect 13648 25452 13728 25480
rect 13544 23044 13596 23050
rect 13544 22986 13596 22992
rect 13556 22574 13584 22986
rect 13544 22568 13596 22574
rect 13544 22510 13596 22516
rect 13648 22098 13676 25452
rect 13728 25434 13780 25440
rect 14844 25362 14872 25842
rect 14832 25356 14884 25362
rect 14832 25298 14884 25304
rect 13912 24404 13964 24410
rect 13912 24346 13964 24352
rect 13728 24064 13780 24070
rect 13728 24006 13780 24012
rect 13740 23730 13768 24006
rect 13728 23724 13780 23730
rect 13728 23666 13780 23672
rect 13636 22094 13688 22098
rect 13556 22092 13688 22094
rect 13556 22066 13636 22092
rect 13452 12368 13504 12374
rect 13452 12310 13504 12316
rect 13556 10674 13584 22066
rect 13636 22034 13688 22040
rect 13740 16658 13768 23666
rect 13924 23526 13952 24346
rect 14740 23588 14792 23594
rect 14740 23530 14792 23536
rect 13912 23520 13964 23526
rect 13912 23462 13964 23468
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 13820 22024 13872 22030
rect 13820 21966 13872 21972
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 13648 15434 13676 16390
rect 13636 15428 13688 15434
rect 13636 15370 13688 15376
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 13648 14385 13676 14894
rect 13634 14376 13690 14385
rect 13634 14311 13690 14320
rect 13648 13870 13676 14311
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13740 11762 13768 13126
rect 13832 12782 13860 21966
rect 14464 21480 14516 21486
rect 14464 21422 14516 21428
rect 14476 20942 14504 21422
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14556 19984 14608 19990
rect 14556 19926 14608 19932
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14476 18834 14504 19110
rect 14464 18828 14516 18834
rect 14464 18770 14516 18776
rect 14372 18692 14424 18698
rect 14372 18634 14424 18640
rect 14004 17604 14056 17610
rect 14004 17546 14056 17552
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13832 9994 13860 12242
rect 13924 10810 13952 13806
rect 14016 12322 14044 17546
rect 14186 17232 14242 17241
rect 14186 17167 14188 17176
rect 14240 17167 14242 17176
rect 14188 17138 14240 17144
rect 14280 16720 14332 16726
rect 14280 16662 14332 16668
rect 14292 16590 14320 16662
rect 14384 16590 14412 18634
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14568 15706 14596 19926
rect 14660 16522 14688 22578
rect 14648 16516 14700 16522
rect 14648 16458 14700 16464
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14752 15162 14780 23530
rect 14832 23180 14884 23186
rect 14832 23122 14884 23128
rect 14844 21078 14872 23122
rect 14832 21072 14884 21078
rect 14832 21014 14884 21020
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 14372 14544 14424 14550
rect 14372 14486 14424 14492
rect 14384 14278 14412 14486
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14096 14000 14148 14006
rect 14096 13942 14148 13948
rect 14108 13870 14136 13942
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14016 12294 14228 12322
rect 14200 11762 14228 12294
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 14200 11354 14228 11494
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 14004 9580 14056 9586
rect 14004 9522 14056 9528
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 13556 7818 13584 9046
rect 13544 7812 13596 7818
rect 13544 7754 13596 7760
rect 13556 7546 13584 7754
rect 13544 7540 13596 7546
rect 13544 7482 13596 7488
rect 14016 6322 14044 9522
rect 14292 7410 14320 13262
rect 14660 12986 14688 14894
rect 14648 12980 14700 12986
rect 14648 12922 14700 12928
rect 14844 12434 14872 21014
rect 15028 18329 15056 26279
rect 15120 26246 15148 30534
rect 15856 30326 15884 30738
rect 15844 30320 15896 30326
rect 15290 30288 15346 30297
rect 15844 30262 15896 30268
rect 15290 30223 15292 30232
rect 15344 30223 15346 30232
rect 15292 30194 15344 30200
rect 15200 30048 15252 30054
rect 15200 29990 15252 29996
rect 15212 29714 15240 29990
rect 15856 29714 15884 30262
rect 15200 29708 15252 29714
rect 15200 29650 15252 29656
rect 15844 29708 15896 29714
rect 15844 29650 15896 29656
rect 15856 29322 15884 29650
rect 15936 29640 15988 29646
rect 15988 29600 16068 29628
rect 15936 29582 15988 29588
rect 15764 29306 15884 29322
rect 16040 29306 16068 29600
rect 15752 29300 15884 29306
rect 15804 29294 15884 29300
rect 16028 29300 16080 29306
rect 15752 29242 15804 29248
rect 16028 29242 16080 29248
rect 15764 28626 15792 29242
rect 15752 28620 15804 28626
rect 15752 28562 15804 28568
rect 15764 28506 15792 28562
rect 15764 28478 15884 28506
rect 15856 28082 15884 28478
rect 15844 28076 15896 28082
rect 15844 28018 15896 28024
rect 15476 28008 15528 28014
rect 15476 27950 15528 27956
rect 15108 26240 15160 26246
rect 15108 26182 15160 26188
rect 15384 25288 15436 25294
rect 15384 25230 15436 25236
rect 15396 24614 15424 25230
rect 15488 25106 15516 27950
rect 15752 26376 15804 26382
rect 15752 26318 15804 26324
rect 15764 25838 15792 26318
rect 15752 25832 15804 25838
rect 15752 25774 15804 25780
rect 15764 25294 15792 25774
rect 15752 25288 15804 25294
rect 15752 25230 15804 25236
rect 15752 25152 15804 25158
rect 15488 25078 15608 25106
rect 15752 25094 15804 25100
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 15488 24721 15516 24754
rect 15474 24712 15530 24721
rect 15474 24647 15530 24656
rect 15384 24608 15436 24614
rect 15384 24550 15436 24556
rect 15396 24206 15424 24550
rect 15384 24200 15436 24206
rect 15384 24142 15436 24148
rect 15396 23662 15424 24142
rect 15384 23656 15436 23662
rect 15384 23598 15436 23604
rect 15200 23316 15252 23322
rect 15200 23258 15252 23264
rect 15212 21486 15240 23258
rect 15292 23112 15344 23118
rect 15396 23100 15424 23598
rect 15476 23112 15528 23118
rect 15396 23072 15476 23100
rect 15292 23054 15344 23060
rect 15476 23054 15528 23060
rect 15304 22710 15332 23054
rect 15488 22778 15516 23054
rect 15476 22772 15528 22778
rect 15476 22714 15528 22720
rect 15292 22704 15344 22710
rect 15292 22646 15344 22652
rect 15200 21480 15252 21486
rect 15200 21422 15252 21428
rect 15108 20868 15160 20874
rect 15108 20810 15160 20816
rect 15120 20398 15148 20810
rect 15108 20392 15160 20398
rect 15108 20334 15160 20340
rect 15120 19854 15148 20334
rect 15108 19848 15160 19854
rect 15108 19790 15160 19796
rect 15120 19446 15148 19790
rect 15384 19780 15436 19786
rect 15384 19722 15436 19728
rect 15108 19440 15160 19446
rect 15108 19382 15160 19388
rect 15120 18766 15148 19382
rect 15108 18760 15160 18766
rect 15108 18702 15160 18708
rect 15014 18320 15070 18329
rect 15120 18290 15148 18702
rect 15014 18255 15070 18264
rect 15108 18284 15160 18290
rect 15108 18226 15160 18232
rect 15120 17746 15148 18226
rect 15396 18222 15424 19722
rect 15580 18698 15608 25078
rect 15764 24954 15792 25094
rect 15752 24948 15804 24954
rect 15752 24890 15804 24896
rect 15764 23050 15792 24890
rect 16132 24698 16160 31726
rect 16224 30190 16252 32166
rect 16212 30184 16264 30190
rect 16212 30126 16264 30132
rect 16316 29034 16344 32302
rect 16408 32230 16436 32778
rect 16500 32434 16528 33458
rect 16776 32502 16804 36178
rect 16856 36032 16908 36038
rect 16856 35974 16908 35980
rect 16868 34202 16896 35974
rect 16856 34196 16908 34202
rect 16856 34138 16908 34144
rect 16764 32496 16816 32502
rect 16764 32438 16816 32444
rect 16488 32428 16540 32434
rect 16488 32370 16540 32376
rect 16396 32224 16448 32230
rect 16396 32166 16448 32172
rect 16500 31906 16528 32370
rect 16868 32042 16896 34138
rect 16960 33930 16988 37062
rect 17132 36576 17184 36582
rect 17184 36536 17264 36564
rect 17132 36518 17184 36524
rect 17236 35766 17264 36536
rect 17512 36310 17540 37198
rect 18510 36952 18566 36961
rect 18510 36887 18512 36896
rect 18564 36887 18566 36896
rect 18512 36858 18564 36864
rect 18616 36802 18644 37198
rect 18524 36774 18644 36802
rect 17592 36712 17644 36718
rect 17592 36654 17644 36660
rect 17684 36712 17736 36718
rect 17684 36654 17736 36660
rect 17500 36304 17552 36310
rect 17500 36246 17552 36252
rect 17406 36000 17462 36009
rect 17406 35935 17462 35944
rect 17420 35766 17448 35935
rect 17224 35760 17276 35766
rect 17224 35702 17276 35708
rect 17408 35760 17460 35766
rect 17408 35702 17460 35708
rect 17236 35630 17264 35702
rect 17132 35624 17184 35630
rect 17132 35566 17184 35572
rect 17224 35624 17276 35630
rect 17224 35566 17276 35572
rect 17144 35222 17172 35566
rect 17604 35290 17632 36654
rect 17408 35284 17460 35290
rect 17408 35226 17460 35232
rect 17592 35284 17644 35290
rect 17592 35226 17644 35232
rect 17132 35216 17184 35222
rect 17132 35158 17184 35164
rect 17316 35148 17368 35154
rect 17316 35090 17368 35096
rect 17130 35048 17186 35057
rect 17130 34983 17186 34992
rect 17144 34202 17172 34983
rect 17328 34474 17356 35090
rect 17420 34610 17448 35226
rect 17696 35018 17724 36654
rect 18524 36174 18552 36774
rect 18604 36576 18656 36582
rect 18604 36518 18656 36524
rect 18512 36168 18564 36174
rect 18510 36136 18512 36145
rect 18564 36136 18566 36145
rect 18510 36071 18566 36080
rect 17960 36032 18012 36038
rect 17960 35974 18012 35980
rect 17684 35012 17736 35018
rect 17684 34954 17736 34960
rect 17776 35012 17828 35018
rect 17776 34954 17828 34960
rect 17684 34672 17736 34678
rect 17684 34614 17736 34620
rect 17408 34604 17460 34610
rect 17408 34546 17460 34552
rect 17500 34536 17552 34542
rect 17500 34478 17552 34484
rect 17316 34468 17368 34474
rect 17316 34410 17368 34416
rect 17132 34196 17184 34202
rect 17132 34138 17184 34144
rect 17144 34066 17172 34138
rect 17132 34060 17184 34066
rect 17132 34002 17184 34008
rect 17408 34060 17460 34066
rect 17408 34002 17460 34008
rect 16948 33924 17000 33930
rect 16948 33866 17000 33872
rect 17040 33924 17092 33930
rect 17040 33866 17092 33872
rect 17052 33658 17080 33866
rect 17040 33652 17092 33658
rect 17040 33594 17092 33600
rect 17420 33590 17448 34002
rect 17512 33697 17540 34478
rect 17498 33688 17554 33697
rect 17498 33623 17554 33632
rect 17408 33584 17460 33590
rect 17408 33526 17460 33532
rect 17696 33454 17724 34614
rect 17592 33448 17644 33454
rect 17592 33390 17644 33396
rect 17684 33448 17736 33454
rect 17684 33390 17736 33396
rect 17316 32972 17368 32978
rect 17316 32914 17368 32920
rect 17328 32881 17356 32914
rect 17408 32904 17460 32910
rect 17314 32872 17370 32881
rect 17408 32846 17460 32852
rect 17314 32807 17370 32816
rect 17132 32768 17184 32774
rect 17132 32710 17184 32716
rect 17040 32496 17092 32502
rect 17040 32438 17092 32444
rect 16948 32224 17000 32230
rect 17052 32178 17080 32438
rect 17144 32230 17172 32710
rect 17420 32502 17448 32846
rect 17604 32774 17632 33390
rect 17684 33108 17736 33114
rect 17684 33050 17736 33056
rect 17592 32768 17644 32774
rect 17592 32710 17644 32716
rect 17408 32496 17460 32502
rect 17408 32438 17460 32444
rect 17224 32360 17276 32366
rect 17224 32302 17276 32308
rect 17000 32172 17080 32178
rect 16948 32166 17080 32172
rect 17132 32224 17184 32230
rect 17132 32166 17184 32172
rect 16960 32150 17080 32166
rect 16868 32014 16988 32042
rect 16408 31890 16528 31906
rect 16396 31884 16528 31890
rect 16448 31878 16528 31884
rect 16672 31884 16724 31890
rect 16396 31826 16448 31832
rect 16672 31826 16724 31832
rect 16684 31754 16712 31826
rect 16580 31748 16712 31754
rect 16632 31726 16712 31748
rect 16580 31690 16632 31696
rect 16408 31198 16712 31226
rect 16408 31142 16436 31198
rect 16396 31136 16448 31142
rect 16396 31078 16448 31084
rect 16488 31136 16540 31142
rect 16488 31078 16540 31084
rect 16396 30048 16448 30054
rect 16396 29990 16448 29996
rect 16304 29028 16356 29034
rect 16304 28970 16356 28976
rect 16212 28756 16264 28762
rect 16212 28698 16264 28704
rect 16224 28490 16252 28698
rect 16212 28484 16264 28490
rect 16212 28426 16264 28432
rect 16224 28393 16252 28426
rect 16210 28384 16266 28393
rect 16210 28319 16266 28328
rect 15856 24670 16160 24698
rect 15752 23044 15804 23050
rect 15752 22986 15804 22992
rect 15856 22438 15884 24670
rect 15936 24608 15988 24614
rect 15936 24550 15988 24556
rect 15844 22432 15896 22438
rect 15844 22374 15896 22380
rect 15856 22094 15884 22374
rect 15764 22066 15884 22094
rect 15568 18692 15620 18698
rect 15568 18634 15620 18640
rect 15476 18352 15528 18358
rect 15476 18294 15528 18300
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 15108 17740 15160 17746
rect 15108 17682 15160 17688
rect 15396 15162 15424 18158
rect 15488 15706 15516 18294
rect 15580 18222 15608 18634
rect 15568 18216 15620 18222
rect 15568 18158 15620 18164
rect 15764 16998 15792 22066
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15856 21146 15884 21490
rect 15844 21140 15896 21146
rect 15844 21082 15896 21088
rect 15948 17882 15976 24550
rect 16304 22160 16356 22166
rect 16304 22102 16356 22108
rect 16212 21684 16264 21690
rect 16212 21626 16264 21632
rect 16120 21616 16172 21622
rect 16120 21558 16172 21564
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 15752 16992 15804 16998
rect 15752 16934 15804 16940
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 15476 15496 15528 15502
rect 15474 15464 15476 15473
rect 15528 15464 15530 15473
rect 15856 15434 15884 15642
rect 15474 15399 15530 15408
rect 15844 15428 15896 15434
rect 15844 15370 15896 15376
rect 15948 15366 15976 17818
rect 15936 15360 15988 15366
rect 16132 15348 16160 21558
rect 16224 19242 16252 21626
rect 16212 19236 16264 19242
rect 16212 19178 16264 19184
rect 16212 18216 16264 18222
rect 16212 18158 16264 18164
rect 15936 15302 15988 15308
rect 16040 15320 16160 15348
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 16040 15026 16068 15320
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 16132 14958 16160 15098
rect 16120 14952 16172 14958
rect 16120 14894 16172 14900
rect 15844 14884 15896 14890
rect 15844 14826 15896 14832
rect 15856 14550 15884 14826
rect 16028 14816 16080 14822
rect 16028 14758 16080 14764
rect 15844 14544 15896 14550
rect 15844 14486 15896 14492
rect 16040 14482 16068 14758
rect 15016 14476 15068 14482
rect 15016 14418 15068 14424
rect 16028 14476 16080 14482
rect 16028 14418 16080 14424
rect 14476 12406 14872 12434
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 14384 11898 14412 12242
rect 14372 11892 14424 11898
rect 14372 11834 14424 11840
rect 14476 9586 14504 12406
rect 14740 12164 14792 12170
rect 14740 12106 14792 12112
rect 14752 11898 14780 12106
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14556 11756 14608 11762
rect 14556 11698 14608 11704
rect 14568 10674 14596 11698
rect 14648 11280 14700 11286
rect 14648 11222 14700 11228
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14476 8974 14504 9318
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14660 8498 14688 11222
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14752 7954 14780 9590
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14752 6866 14780 7890
rect 14832 7812 14884 7818
rect 14832 7754 14884 7760
rect 14844 7546 14872 7754
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 14384 5914 14412 6734
rect 15028 6662 15056 14418
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 15212 13841 15240 14282
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15198 13832 15254 13841
rect 15198 13767 15254 13776
rect 15212 12646 15240 13767
rect 15764 13258 15792 13942
rect 15568 13252 15620 13258
rect 15568 13194 15620 13200
rect 15752 13252 15804 13258
rect 15752 13194 15804 13200
rect 15580 12986 15608 13194
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15384 12844 15436 12850
rect 15384 12786 15436 12792
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 15396 12442 15424 12786
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 15672 11150 15700 11630
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 15764 9994 15792 13194
rect 16132 12238 16160 14894
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16028 11620 16080 11626
rect 16028 11562 16080 11568
rect 15752 9988 15804 9994
rect 15752 9930 15804 9936
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15396 8634 15424 9454
rect 15476 8900 15528 8906
rect 15476 8842 15528 8848
rect 15488 8634 15516 8842
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15660 8356 15712 8362
rect 15660 8298 15712 8304
rect 15672 7886 15700 8298
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 15580 6322 15608 7346
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15672 6458 15700 6734
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 14372 5908 14424 5914
rect 14372 5850 14424 5856
rect 15764 5370 15792 9930
rect 15936 9036 15988 9042
rect 15936 8978 15988 8984
rect 15948 8945 15976 8978
rect 15934 8936 15990 8945
rect 15934 8871 15990 8880
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 16040 5302 16068 11562
rect 16224 9042 16252 18158
rect 16316 16590 16344 22102
rect 16408 21622 16436 29990
rect 16500 29238 16528 31078
rect 16684 30802 16712 31198
rect 16580 30796 16632 30802
rect 16580 30738 16632 30744
rect 16672 30796 16724 30802
rect 16672 30738 16724 30744
rect 16592 30054 16620 30738
rect 16764 30388 16816 30394
rect 16764 30330 16816 30336
rect 16580 30048 16632 30054
rect 16580 29990 16632 29996
rect 16488 29232 16540 29238
rect 16488 29174 16540 29180
rect 16488 29028 16540 29034
rect 16488 28970 16540 28976
rect 16500 27130 16528 28970
rect 16488 27124 16540 27130
rect 16488 27066 16540 27072
rect 16488 26988 16540 26994
rect 16488 26930 16540 26936
rect 16500 23866 16528 26930
rect 16776 25906 16804 30330
rect 16764 25900 16816 25906
rect 16764 25842 16816 25848
rect 16672 25696 16724 25702
rect 16672 25638 16724 25644
rect 16580 25356 16632 25362
rect 16580 25298 16632 25304
rect 16592 24070 16620 25298
rect 16580 24064 16632 24070
rect 16580 24006 16632 24012
rect 16488 23860 16540 23866
rect 16488 23802 16540 23808
rect 16580 22704 16632 22710
rect 16580 22646 16632 22652
rect 16488 22432 16540 22438
rect 16488 22374 16540 22380
rect 16500 22166 16528 22374
rect 16488 22160 16540 22166
rect 16488 22102 16540 22108
rect 16396 21616 16448 21622
rect 16396 21558 16448 21564
rect 16488 19440 16540 19446
rect 16488 19382 16540 19388
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 16408 18630 16436 19110
rect 16396 18624 16448 18630
rect 16396 18566 16448 18572
rect 16408 16998 16436 18566
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16304 16584 16356 16590
rect 16304 16526 16356 16532
rect 16396 16244 16448 16250
rect 16396 16186 16448 16192
rect 16304 15700 16356 15706
rect 16304 15642 16356 15648
rect 16316 15434 16344 15642
rect 16304 15428 16356 15434
rect 16304 15370 16356 15376
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 16316 14074 16344 14418
rect 16408 14346 16436 16186
rect 16500 15162 16528 19382
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16396 14340 16448 14346
rect 16396 14282 16448 14288
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 16396 13456 16448 13462
rect 16396 13398 16448 13404
rect 16304 13252 16356 13258
rect 16304 13194 16356 13200
rect 16316 12306 16344 13194
rect 16408 12714 16436 13398
rect 16396 12708 16448 12714
rect 16396 12650 16448 12656
rect 16304 12300 16356 12306
rect 16304 12242 16356 12248
rect 16212 9036 16264 9042
rect 16212 8978 16264 8984
rect 16224 8498 16252 8978
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 16592 6322 16620 22646
rect 16684 17882 16712 25638
rect 16764 24880 16816 24886
rect 16816 24828 16896 24834
rect 16764 24822 16896 24828
rect 16776 24806 16896 24822
rect 16764 24676 16816 24682
rect 16764 24618 16816 24624
rect 16776 21078 16804 24618
rect 16868 23730 16896 24806
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 16868 23633 16896 23666
rect 16854 23624 16910 23633
rect 16854 23559 16910 23568
rect 16960 23254 16988 32014
rect 16948 23248 17000 23254
rect 16948 23190 17000 23196
rect 17052 22642 17080 32150
rect 17132 30864 17184 30870
rect 17132 30806 17184 30812
rect 17144 30598 17172 30806
rect 17132 30592 17184 30598
rect 17132 30534 17184 30540
rect 17236 30394 17264 32302
rect 17604 31754 17632 32710
rect 17696 31822 17724 33050
rect 17788 32774 17816 34954
rect 17972 32842 18000 35974
rect 18616 35222 18644 36518
rect 18708 35834 18736 39200
rect 19432 37392 19484 37398
rect 19432 37334 19484 37340
rect 19444 37262 19472 37334
rect 18788 37256 18840 37262
rect 18788 37198 18840 37204
rect 19432 37256 19484 37262
rect 19432 37198 19484 37204
rect 18696 35828 18748 35834
rect 18696 35770 18748 35776
rect 18696 35692 18748 35698
rect 18696 35634 18748 35640
rect 18708 35222 18736 35634
rect 18604 35216 18656 35222
rect 18604 35158 18656 35164
rect 18696 35216 18748 35222
rect 18696 35158 18748 35164
rect 18328 34944 18380 34950
rect 18328 34886 18380 34892
rect 18050 34776 18106 34785
rect 18050 34711 18106 34720
rect 18064 34678 18092 34711
rect 18052 34672 18104 34678
rect 18052 34614 18104 34620
rect 18144 34536 18196 34542
rect 18064 34484 18144 34490
rect 18064 34478 18196 34484
rect 18064 34462 18184 34478
rect 18064 33998 18092 34462
rect 18144 34400 18196 34406
rect 18144 34342 18196 34348
rect 18236 34400 18288 34406
rect 18236 34342 18288 34348
rect 18156 33998 18184 34342
rect 18248 34202 18276 34342
rect 18236 34196 18288 34202
rect 18236 34138 18288 34144
rect 18052 33992 18104 33998
rect 18052 33934 18104 33940
rect 18144 33992 18196 33998
rect 18144 33934 18196 33940
rect 17960 32836 18012 32842
rect 17960 32778 18012 32784
rect 17776 32768 17828 32774
rect 17776 32710 17828 32716
rect 17788 32366 17816 32710
rect 17776 32360 17828 32366
rect 17776 32302 17828 32308
rect 17866 31920 17922 31929
rect 17776 31884 17828 31890
rect 17866 31855 17868 31864
rect 17776 31826 17828 31832
rect 17920 31855 17922 31864
rect 17868 31826 17920 31832
rect 17684 31816 17736 31822
rect 17684 31758 17736 31764
rect 17328 31726 17632 31754
rect 17224 30388 17276 30394
rect 17224 30330 17276 30336
rect 17328 30274 17356 31726
rect 17788 31634 17816 31826
rect 17420 31606 17816 31634
rect 17960 31680 18012 31686
rect 17960 31622 18012 31628
rect 17420 30297 17448 31606
rect 17776 31408 17828 31414
rect 17828 31368 17908 31396
rect 17776 31350 17828 31356
rect 17500 31340 17552 31346
rect 17500 31282 17552 31288
rect 17512 30954 17540 31282
rect 17880 31278 17908 31368
rect 17868 31272 17920 31278
rect 17868 31214 17920 31220
rect 17512 30926 17724 30954
rect 17696 30870 17724 30926
rect 17684 30864 17736 30870
rect 17684 30806 17736 30812
rect 17972 30666 18000 31622
rect 18340 31260 18368 34886
rect 18510 34368 18566 34377
rect 18510 34303 18566 34312
rect 18524 34202 18552 34303
rect 18512 34196 18564 34202
rect 18512 34138 18564 34144
rect 18512 33312 18564 33318
rect 18512 33254 18564 33260
rect 18524 31958 18552 33254
rect 18616 32842 18644 35158
rect 18708 34678 18736 35158
rect 18696 34672 18748 34678
rect 18696 34614 18748 34620
rect 18696 34536 18748 34542
rect 18696 34478 18748 34484
rect 18604 32836 18656 32842
rect 18604 32778 18656 32784
rect 18512 31952 18564 31958
rect 18418 31920 18474 31929
rect 18512 31894 18564 31900
rect 18418 31855 18474 31864
rect 18248 31232 18368 31260
rect 17960 30660 18012 30666
rect 17960 30602 18012 30608
rect 18052 30660 18104 30666
rect 18052 30602 18104 30608
rect 17776 30592 17828 30598
rect 17776 30534 17828 30540
rect 17144 30246 17356 30274
rect 17406 30288 17462 30297
rect 17144 29306 17172 30246
rect 17406 30223 17462 30232
rect 17224 30184 17276 30190
rect 17276 30144 17356 30172
rect 17224 30126 17276 30132
rect 17328 29782 17356 30144
rect 17316 29776 17368 29782
rect 17316 29718 17368 29724
rect 17222 29472 17278 29481
rect 17222 29407 17278 29416
rect 17132 29300 17184 29306
rect 17132 29242 17184 29248
rect 17132 26784 17184 26790
rect 17132 26726 17184 26732
rect 17144 26382 17172 26726
rect 17236 26489 17264 29407
rect 17314 28792 17370 28801
rect 17314 28727 17316 28736
rect 17368 28727 17370 28736
rect 17316 28698 17368 28704
rect 17222 26480 17278 26489
rect 17222 26415 17278 26424
rect 17132 26376 17184 26382
rect 17132 26318 17184 26324
rect 17236 26194 17264 26415
rect 17144 26166 17264 26194
rect 17144 25838 17172 26166
rect 17224 25968 17276 25974
rect 17224 25910 17276 25916
rect 17236 25838 17264 25910
rect 17132 25832 17184 25838
rect 17132 25774 17184 25780
rect 17224 25832 17276 25838
rect 17224 25774 17276 25780
rect 17224 24744 17276 24750
rect 17224 24686 17276 24692
rect 17132 24676 17184 24682
rect 17132 24618 17184 24624
rect 17144 24585 17172 24618
rect 17130 24576 17186 24585
rect 17130 24511 17186 24520
rect 17132 24064 17184 24070
rect 17132 24006 17184 24012
rect 17040 22636 17092 22642
rect 17040 22578 17092 22584
rect 17144 21350 17172 24006
rect 17236 23594 17264 24686
rect 17224 23588 17276 23594
rect 17224 23530 17276 23536
rect 17224 22976 17276 22982
rect 17224 22918 17276 22924
rect 17328 22930 17356 28698
rect 17420 25945 17448 30223
rect 17500 30184 17552 30190
rect 17500 30126 17552 30132
rect 17512 28422 17540 30126
rect 17682 29880 17738 29889
rect 17682 29815 17738 29824
rect 17696 29510 17724 29815
rect 17684 29504 17736 29510
rect 17684 29446 17736 29452
rect 17696 29186 17724 29446
rect 17604 29158 17724 29186
rect 17500 28416 17552 28422
rect 17500 28358 17552 28364
rect 17604 28234 17632 29158
rect 17684 28756 17736 28762
rect 17684 28698 17736 28704
rect 17512 28206 17632 28234
rect 17406 25936 17462 25945
rect 17406 25871 17462 25880
rect 17406 24712 17462 24721
rect 17406 24647 17408 24656
rect 17460 24647 17462 24656
rect 17408 24618 17460 24624
rect 17512 24596 17540 28206
rect 17696 28014 17724 28698
rect 17684 28008 17736 28014
rect 17684 27950 17736 27956
rect 17684 27396 17736 27402
rect 17684 27338 17736 27344
rect 17696 27130 17724 27338
rect 17684 27124 17736 27130
rect 17684 27066 17736 27072
rect 17592 26988 17644 26994
rect 17592 26930 17644 26936
rect 17604 26382 17632 26930
rect 17684 26920 17736 26926
rect 17684 26862 17736 26868
rect 17696 26466 17724 26862
rect 17788 26586 17816 30534
rect 18064 30410 18092 30602
rect 17972 30382 18092 30410
rect 17868 29232 17920 29238
rect 17972 29220 18000 30382
rect 18144 30116 18196 30122
rect 18144 30058 18196 30064
rect 18156 29782 18184 30058
rect 18144 29776 18196 29782
rect 18144 29718 18196 29724
rect 18052 29640 18104 29646
rect 18052 29582 18104 29588
rect 18064 29510 18092 29582
rect 18052 29504 18104 29510
rect 18052 29446 18104 29452
rect 18248 29322 18276 31232
rect 18328 30728 18380 30734
rect 18328 30670 18380 30676
rect 17920 29192 18000 29220
rect 18064 29294 18276 29322
rect 17868 29174 17920 29180
rect 17960 27872 18012 27878
rect 17960 27814 18012 27820
rect 17776 26580 17828 26586
rect 17776 26522 17828 26528
rect 17868 26580 17920 26586
rect 17868 26522 17920 26528
rect 17880 26466 17908 26522
rect 17696 26438 17908 26466
rect 17592 26376 17644 26382
rect 17592 26318 17644 26324
rect 17774 26344 17830 26353
rect 17604 24750 17632 26318
rect 17774 26279 17776 26288
rect 17828 26279 17830 26288
rect 17776 26250 17828 26256
rect 17972 26042 18000 27814
rect 17960 26036 18012 26042
rect 17960 25978 18012 25984
rect 17592 24744 17644 24750
rect 17592 24686 17644 24692
rect 17512 24568 17908 24596
rect 18064 24585 18092 29294
rect 18144 29232 18196 29238
rect 18144 29174 18196 29180
rect 18236 29232 18288 29238
rect 18236 29174 18288 29180
rect 18156 29073 18184 29174
rect 18248 29102 18276 29174
rect 18236 29096 18288 29102
rect 18142 29064 18198 29073
rect 18236 29038 18288 29044
rect 18142 28999 18198 29008
rect 18236 28960 18288 28966
rect 18236 28902 18288 28908
rect 18144 28688 18196 28694
rect 18144 28630 18196 28636
rect 18156 27606 18184 28630
rect 18248 28393 18276 28902
rect 18234 28384 18290 28393
rect 18234 28319 18290 28328
rect 18248 27860 18276 28319
rect 18340 28014 18368 30670
rect 18432 29102 18460 31855
rect 18524 29102 18552 31894
rect 18708 30841 18736 34478
rect 18800 33590 18828 37198
rect 19340 37120 19392 37126
rect 19340 37062 19392 37068
rect 19352 36904 19380 37062
rect 19260 36876 19380 36904
rect 19444 36904 19472 37198
rect 19996 37126 20024 39200
rect 21088 37392 21140 37398
rect 21088 37334 21140 37340
rect 20076 37256 20128 37262
rect 20076 37198 20128 37204
rect 20350 37224 20406 37233
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19444 36876 19564 36904
rect 19260 36666 19288 36876
rect 19536 36786 19564 36876
rect 19340 36780 19392 36786
rect 19524 36780 19576 36786
rect 19392 36740 19472 36768
rect 19340 36722 19392 36728
rect 19260 36638 19380 36666
rect 19352 35873 19380 36638
rect 19338 35864 19394 35873
rect 19338 35799 19394 35808
rect 18880 35488 18932 35494
rect 18880 35430 18932 35436
rect 19340 35488 19392 35494
rect 19340 35430 19392 35436
rect 18892 35290 18920 35430
rect 18880 35284 18932 35290
rect 18880 35226 18932 35232
rect 18880 34944 18932 34950
rect 18880 34886 18932 34892
rect 18788 33584 18840 33590
rect 18892 33561 18920 34886
rect 19352 34762 19380 35430
rect 19168 34734 19380 34762
rect 18972 34672 19024 34678
rect 18972 34614 19024 34620
rect 18788 33526 18840 33532
rect 18878 33552 18934 33561
rect 18878 33487 18934 33496
rect 18788 31272 18840 31278
rect 18786 31240 18788 31249
rect 18840 31240 18842 31249
rect 18786 31175 18842 31184
rect 18694 30832 18750 30841
rect 18694 30767 18750 30776
rect 18788 30592 18840 30598
rect 18788 30534 18840 30540
rect 18604 30048 18656 30054
rect 18604 29990 18656 29996
rect 18696 30048 18748 30054
rect 18696 29990 18748 29996
rect 18616 29782 18644 29990
rect 18604 29776 18656 29782
rect 18604 29718 18656 29724
rect 18420 29096 18472 29102
rect 18420 29038 18472 29044
rect 18512 29096 18564 29102
rect 18512 29038 18564 29044
rect 18512 28552 18564 28558
rect 18512 28494 18564 28500
rect 18420 28076 18472 28082
rect 18420 28018 18472 28024
rect 18328 28008 18380 28014
rect 18328 27950 18380 27956
rect 18248 27832 18368 27860
rect 18144 27600 18196 27606
rect 18144 27542 18196 27548
rect 18144 27056 18196 27062
rect 18144 26998 18196 27004
rect 18156 26042 18184 26998
rect 18144 26036 18196 26042
rect 18144 25978 18196 25984
rect 18236 24608 18288 24614
rect 17406 23080 17462 23089
rect 17406 23015 17408 23024
rect 17460 23015 17462 23024
rect 17408 22986 17460 22992
rect 17684 22976 17736 22982
rect 17236 22778 17264 22918
rect 17328 22902 17448 22930
rect 17684 22918 17736 22924
rect 17224 22772 17276 22778
rect 17224 22714 17276 22720
rect 17316 22092 17368 22098
rect 17316 22034 17368 22040
rect 17132 21344 17184 21350
rect 17132 21286 17184 21292
rect 16764 21072 16816 21078
rect 16764 21014 16816 21020
rect 17144 20806 17172 21286
rect 17040 20800 17092 20806
rect 17040 20742 17092 20748
rect 17132 20800 17184 20806
rect 17132 20742 17184 20748
rect 17052 20466 17080 20742
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 16764 19780 16816 19786
rect 16764 19722 16816 19728
rect 16776 19514 16804 19722
rect 16856 19712 16908 19718
rect 16856 19654 16908 19660
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16764 18352 16816 18358
rect 16764 18294 16816 18300
rect 16672 17876 16724 17882
rect 16672 17818 16724 17824
rect 16672 16448 16724 16454
rect 16672 16390 16724 16396
rect 16684 16182 16712 16390
rect 16672 16176 16724 16182
rect 16672 16118 16724 16124
rect 16776 15706 16804 18294
rect 16868 17746 16896 19654
rect 17132 18216 17184 18222
rect 17132 18158 17184 18164
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 17040 17604 17092 17610
rect 17040 17546 17092 17552
rect 17052 16522 17080 17546
rect 17144 16674 17172 18158
rect 17224 17264 17276 17270
rect 17222 17232 17224 17241
rect 17276 17232 17278 17241
rect 17222 17167 17278 17176
rect 17224 17060 17276 17066
rect 17224 17002 17276 17008
rect 17236 16794 17264 17002
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 17144 16646 17264 16674
rect 17040 16516 17092 16522
rect 17040 16458 17092 16464
rect 16764 15700 16816 15706
rect 16764 15642 16816 15648
rect 17040 15496 17092 15502
rect 17038 15464 17040 15473
rect 17092 15464 17094 15473
rect 17038 15399 17094 15408
rect 17052 15026 17080 15399
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 16672 14476 16724 14482
rect 16672 14418 16724 14424
rect 16684 13938 16712 14418
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 17132 13864 17184 13870
rect 17132 13806 17184 13812
rect 16672 13524 16724 13530
rect 16672 13466 16724 13472
rect 16684 13190 16712 13466
rect 16672 13184 16724 13190
rect 16672 13126 16724 13132
rect 16856 13184 16908 13190
rect 16856 13126 16908 13132
rect 16868 12986 16896 13126
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 17052 11898 17080 12786
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 17052 11082 17080 11290
rect 17040 11076 17092 11082
rect 17040 11018 17092 11024
rect 17144 9654 17172 13806
rect 17236 13376 17264 16646
rect 17328 13938 17356 22034
rect 17420 20534 17448 22902
rect 17696 20874 17724 22918
rect 17776 22568 17828 22574
rect 17774 22536 17776 22545
rect 17828 22536 17830 22545
rect 17774 22471 17830 22480
rect 17880 22094 17908 24568
rect 18050 24576 18106 24585
rect 18236 24550 18288 24556
rect 18050 24511 18106 24520
rect 18144 24064 18196 24070
rect 18144 24006 18196 24012
rect 18156 23798 18184 24006
rect 18144 23792 18196 23798
rect 18144 23734 18196 23740
rect 18248 23118 18276 24550
rect 18236 23112 18288 23118
rect 18236 23054 18288 23060
rect 17788 22066 17908 22094
rect 17788 20942 17816 22066
rect 17960 21888 18012 21894
rect 17960 21830 18012 21836
rect 17776 20936 17828 20942
rect 17776 20878 17828 20884
rect 17684 20868 17736 20874
rect 17684 20810 17736 20816
rect 17972 20602 18000 21830
rect 18340 21554 18368 27832
rect 18432 22574 18460 28018
rect 18524 23050 18552 28494
rect 18708 28150 18736 29990
rect 18800 29510 18828 30534
rect 18984 30394 19012 34614
rect 19064 34196 19116 34202
rect 19064 34138 19116 34144
rect 19076 32552 19104 34138
rect 19168 33833 19196 34734
rect 19248 34604 19300 34610
rect 19248 34546 19300 34552
rect 19260 33862 19288 34546
rect 19340 34536 19392 34542
rect 19340 34478 19392 34484
rect 19352 33930 19380 34478
rect 19444 33998 19472 36740
rect 19524 36722 19576 36728
rect 19984 36032 20036 36038
rect 20088 36009 20116 37198
rect 21100 37194 21128 37334
rect 21284 37262 21312 39200
rect 21364 37664 21416 37670
rect 21364 37606 21416 37612
rect 21272 37256 21324 37262
rect 21272 37198 21324 37204
rect 20350 37159 20406 37168
rect 21088 37188 21140 37194
rect 20168 36168 20220 36174
rect 20168 36110 20220 36116
rect 19984 35974 20036 35980
rect 20074 36000 20130 36009
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19800 35760 19852 35766
rect 19800 35702 19852 35708
rect 19706 35456 19762 35465
rect 19706 35391 19762 35400
rect 19720 35154 19748 35391
rect 19708 35148 19760 35154
rect 19708 35090 19760 35096
rect 19812 35086 19840 35702
rect 19892 35216 19944 35222
rect 19892 35158 19944 35164
rect 19904 35086 19932 35158
rect 19800 35080 19852 35086
rect 19800 35022 19852 35028
rect 19892 35080 19944 35086
rect 19892 35022 19944 35028
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19524 34468 19576 34474
rect 19524 34410 19576 34416
rect 19536 33998 19564 34410
rect 19432 33992 19484 33998
rect 19432 33934 19484 33940
rect 19524 33992 19576 33998
rect 19524 33934 19576 33940
rect 19996 33946 20024 35974
rect 20074 35935 20130 35944
rect 20180 35698 20208 36110
rect 20364 35766 20392 37159
rect 21088 37130 21140 37136
rect 21088 36780 21140 36786
rect 21088 36722 21140 36728
rect 20904 36712 20956 36718
rect 20904 36654 20956 36660
rect 20720 36644 20772 36650
rect 20720 36586 20772 36592
rect 20444 36576 20496 36582
rect 20732 36553 20760 36586
rect 20444 36518 20496 36524
rect 20718 36544 20774 36553
rect 20456 36242 20484 36518
rect 20718 36479 20774 36488
rect 20444 36236 20496 36242
rect 20444 36178 20496 36184
rect 20720 36032 20772 36038
rect 20720 35974 20772 35980
rect 20352 35760 20404 35766
rect 20352 35702 20404 35708
rect 20168 35692 20220 35698
rect 20168 35634 20220 35640
rect 20536 35692 20588 35698
rect 20536 35634 20588 35640
rect 20352 35488 20404 35494
rect 20352 35430 20404 35436
rect 20168 35080 20220 35086
rect 20168 35022 20220 35028
rect 20076 35012 20128 35018
rect 20076 34954 20128 34960
rect 20088 34921 20116 34954
rect 20074 34912 20130 34921
rect 20074 34847 20130 34856
rect 19340 33924 19392 33930
rect 19340 33866 19392 33872
rect 19248 33856 19300 33862
rect 19154 33824 19210 33833
rect 19248 33798 19300 33804
rect 19154 33759 19210 33768
rect 19156 33516 19208 33522
rect 19156 33458 19208 33464
rect 19168 33114 19196 33458
rect 19156 33108 19208 33114
rect 19156 33050 19208 33056
rect 19076 32524 19196 32552
rect 19064 32428 19116 32434
rect 19064 32370 19116 32376
rect 19076 31822 19104 32370
rect 19064 31816 19116 31822
rect 19168 31793 19196 32524
rect 19260 32434 19288 33798
rect 19444 33522 19472 33934
rect 19996 33918 20116 33946
rect 19984 33856 20036 33862
rect 19984 33798 20036 33804
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19522 33552 19578 33561
rect 19432 33516 19484 33522
rect 19522 33487 19578 33496
rect 19432 33458 19484 33464
rect 19340 33312 19392 33318
rect 19340 33254 19392 33260
rect 19248 32428 19300 32434
rect 19248 32370 19300 32376
rect 19248 32224 19300 32230
rect 19248 32166 19300 32172
rect 19064 31758 19116 31764
rect 19154 31784 19210 31793
rect 19076 31362 19104 31758
rect 19154 31719 19210 31728
rect 19076 31334 19196 31362
rect 19064 31272 19116 31278
rect 19064 31214 19116 31220
rect 18972 30388 19024 30394
rect 18972 30330 19024 30336
rect 18972 29640 19024 29646
rect 18972 29582 19024 29588
rect 18788 29504 18840 29510
rect 18788 29446 18840 29452
rect 18880 29504 18932 29510
rect 18880 29446 18932 29452
rect 18892 28490 18920 29446
rect 18984 29073 19012 29582
rect 19076 29345 19104 31214
rect 19168 30598 19196 31334
rect 19156 30592 19208 30598
rect 19156 30534 19208 30540
rect 19062 29336 19118 29345
rect 19062 29271 19118 29280
rect 19168 29186 19196 30534
rect 19260 30326 19288 32166
rect 19352 32026 19380 33254
rect 19340 32020 19392 32026
rect 19340 31962 19392 31968
rect 19340 31680 19392 31686
rect 19340 31622 19392 31628
rect 19352 30734 19380 31622
rect 19340 30728 19392 30734
rect 19340 30670 19392 30676
rect 19352 30394 19380 30670
rect 19340 30388 19392 30394
rect 19340 30330 19392 30336
rect 19248 30320 19300 30326
rect 19248 30262 19300 30268
rect 19444 30258 19472 33458
rect 19536 33046 19564 33487
rect 19706 33416 19762 33425
rect 19706 33351 19762 33360
rect 19720 33318 19748 33351
rect 19708 33312 19760 33318
rect 19708 33254 19760 33260
rect 19524 33040 19576 33046
rect 19892 33040 19944 33046
rect 19524 32982 19576 32988
rect 19628 32988 19892 32994
rect 19628 32982 19944 32988
rect 19628 32978 19932 32982
rect 19996 32978 20024 33798
rect 20088 33590 20116 33918
rect 20076 33584 20128 33590
rect 20076 33526 20128 33532
rect 19616 32972 19932 32978
rect 19668 32966 19932 32972
rect 19984 32972 20036 32978
rect 19616 32914 19668 32920
rect 19984 32914 20036 32920
rect 20076 32904 20128 32910
rect 20076 32846 20128 32852
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19616 32496 19668 32502
rect 19668 32456 19840 32484
rect 19616 32438 19668 32444
rect 19616 32360 19668 32366
rect 19616 32302 19668 32308
rect 19628 32201 19656 32302
rect 19614 32192 19670 32201
rect 19614 32127 19670 32136
rect 19812 31668 19840 32456
rect 19892 32360 19944 32366
rect 19892 32302 19944 32308
rect 19904 32230 19932 32302
rect 19892 32224 19944 32230
rect 19892 32166 19944 32172
rect 20088 31686 20116 32846
rect 20076 31680 20128 31686
rect 19812 31640 20024 31668
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19996 31482 20024 31640
rect 20076 31622 20128 31628
rect 19984 31476 20036 31482
rect 19984 31418 20036 31424
rect 19616 31408 19668 31414
rect 19616 31350 19668 31356
rect 19628 30841 19656 31350
rect 20180 31346 20208 35022
rect 20260 34672 20312 34678
rect 20260 34614 20312 34620
rect 20272 34202 20300 34614
rect 20260 34196 20312 34202
rect 20260 34138 20312 34144
rect 20260 32972 20312 32978
rect 20260 32914 20312 32920
rect 20272 32570 20300 32914
rect 20260 32564 20312 32570
rect 20260 32506 20312 32512
rect 20260 32360 20312 32366
rect 20258 32328 20260 32337
rect 20312 32328 20314 32337
rect 20258 32263 20314 32272
rect 20272 31958 20300 32263
rect 20260 31952 20312 31958
rect 20260 31894 20312 31900
rect 19984 31340 20036 31346
rect 19984 31282 20036 31288
rect 20168 31340 20220 31346
rect 20168 31282 20220 31288
rect 19614 30832 19670 30841
rect 19614 30767 19670 30776
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19996 30258 20024 31282
rect 20168 30932 20220 30938
rect 20168 30874 20220 30880
rect 20180 30666 20208 30874
rect 20364 30802 20392 35430
rect 20444 35148 20496 35154
rect 20444 35090 20496 35096
rect 20456 35057 20484 35090
rect 20442 35048 20498 35057
rect 20442 34983 20498 34992
rect 20548 34610 20576 35634
rect 20628 34944 20680 34950
rect 20628 34886 20680 34892
rect 20536 34604 20588 34610
rect 20536 34546 20588 34552
rect 20444 33856 20496 33862
rect 20444 33798 20496 33804
rect 20456 33590 20484 33798
rect 20444 33584 20496 33590
rect 20444 33526 20496 33532
rect 20548 33436 20576 34546
rect 20640 34134 20668 34886
rect 20732 34649 20760 35974
rect 20812 35760 20864 35766
rect 20812 35702 20864 35708
rect 20718 34640 20774 34649
rect 20718 34575 20774 34584
rect 20720 34468 20772 34474
rect 20720 34410 20772 34416
rect 20628 34128 20680 34134
rect 20628 34070 20680 34076
rect 20628 33992 20680 33998
rect 20628 33934 20680 33940
rect 20456 33408 20576 33436
rect 20352 30796 20404 30802
rect 20352 30738 20404 30744
rect 20168 30660 20220 30666
rect 20168 30602 20220 30608
rect 20076 30388 20128 30394
rect 20076 30330 20128 30336
rect 19432 30252 19484 30258
rect 19432 30194 19484 30200
rect 19524 30252 19576 30258
rect 19524 30194 19576 30200
rect 19984 30252 20036 30258
rect 19984 30194 20036 30200
rect 19444 29288 19472 30194
rect 19536 29646 19564 30194
rect 19524 29640 19576 29646
rect 19524 29582 19576 29588
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19982 29336 20038 29345
rect 19444 29260 19748 29288
rect 19982 29271 20038 29280
rect 19076 29158 19196 29186
rect 19340 29232 19392 29238
rect 19392 29192 19472 29220
rect 19340 29174 19392 29180
rect 18970 29064 19026 29073
rect 18970 28999 19026 29008
rect 18880 28484 18932 28490
rect 18880 28426 18932 28432
rect 18696 28144 18748 28150
rect 18696 28086 18748 28092
rect 18696 27396 18748 27402
rect 18696 27338 18748 27344
rect 18604 25900 18656 25906
rect 18604 25842 18656 25848
rect 18616 25702 18644 25842
rect 18604 25696 18656 25702
rect 18604 25638 18656 25644
rect 18616 25158 18644 25638
rect 18604 25152 18656 25158
rect 18604 25094 18656 25100
rect 18512 23044 18564 23050
rect 18512 22986 18564 22992
rect 18512 22636 18564 22642
rect 18512 22578 18564 22584
rect 18420 22568 18472 22574
rect 18420 22510 18472 22516
rect 18524 22030 18552 22578
rect 18512 22024 18564 22030
rect 18512 21966 18564 21972
rect 18328 21548 18380 21554
rect 18328 21490 18380 21496
rect 18420 21344 18472 21350
rect 18420 21286 18472 21292
rect 18328 20800 18380 20806
rect 18328 20742 18380 20748
rect 17960 20596 18012 20602
rect 17960 20538 18012 20544
rect 17408 20528 17460 20534
rect 17408 20470 17460 20476
rect 18144 20460 18196 20466
rect 18144 20402 18196 20408
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17512 18766 17540 20334
rect 17960 19780 18012 19786
rect 17960 19722 18012 19728
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17512 18222 17540 18702
rect 17500 18216 17552 18222
rect 17500 18158 17552 18164
rect 17604 17610 17632 19246
rect 17684 18896 17736 18902
rect 17684 18838 17736 18844
rect 17696 18698 17724 18838
rect 17684 18692 17736 18698
rect 17684 18634 17736 18640
rect 17774 18320 17830 18329
rect 17774 18255 17830 18264
rect 17684 17808 17736 17814
rect 17684 17750 17736 17756
rect 17592 17604 17644 17610
rect 17592 17546 17644 17552
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17512 13938 17540 16526
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17500 13796 17552 13802
rect 17500 13738 17552 13744
rect 17236 13348 17356 13376
rect 17224 13252 17276 13258
rect 17224 13194 17276 13200
rect 17236 12986 17264 13194
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 17328 12866 17356 13348
rect 17512 13258 17540 13738
rect 17500 13252 17552 13258
rect 17500 13194 17552 13200
rect 17236 12838 17356 12866
rect 17512 12850 17540 13194
rect 17500 12844 17552 12850
rect 17236 11762 17264 12838
rect 17500 12786 17552 12792
rect 17604 12434 17632 17546
rect 17696 13326 17724 17750
rect 17788 17202 17816 18255
rect 17868 17876 17920 17882
rect 17868 17818 17920 17824
rect 17880 17202 17908 17818
rect 17972 17338 18000 19722
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 17960 17332 18012 17338
rect 17960 17274 18012 17280
rect 17776 17196 17828 17202
rect 17776 17138 17828 17144
rect 17868 17196 17920 17202
rect 17868 17138 17920 17144
rect 17776 16992 17828 16998
rect 17960 16992 18012 16998
rect 17776 16934 17828 16940
rect 17880 16952 17960 16980
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17788 13002 17816 16934
rect 17880 15502 17908 16952
rect 17960 16934 18012 16940
rect 17960 16176 18012 16182
rect 17960 16118 18012 16124
rect 17972 15706 18000 16118
rect 17960 15700 18012 15706
rect 17960 15642 18012 15648
rect 18064 15502 18092 18906
rect 18156 18222 18184 20402
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 17868 15496 17920 15502
rect 17868 15438 17920 15444
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 18156 15366 18184 15642
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 17788 12974 17908 13002
rect 17880 12918 17908 12974
rect 17868 12912 17920 12918
rect 17868 12854 17920 12860
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17420 12406 17632 12434
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 17132 9648 17184 9654
rect 17132 9590 17184 9596
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 16028 5296 16080 5302
rect 16028 5238 16080 5244
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 10416 2576 10468 2582
rect 10416 2518 10468 2524
rect 12348 2576 12400 2582
rect 12348 2518 12400 2524
rect 13268 2576 13320 2582
rect 13268 2518 13320 2524
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 10980 800 11008 2382
rect 11624 800 11652 2382
rect 12912 800 12940 2382
rect 14200 800 14228 2994
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 14936 2446 14964 2790
rect 16868 2650 16896 8774
rect 17236 8566 17264 11698
rect 17328 11082 17356 12038
rect 17316 11076 17368 11082
rect 17316 11018 17368 11024
rect 17420 9994 17448 12406
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 17696 10810 17724 11154
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17788 10130 17816 10406
rect 17880 10130 17908 12718
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 18248 11082 18276 11494
rect 18236 11076 18288 11082
rect 18236 11018 18288 11024
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 17684 9512 17736 9518
rect 17684 9454 17736 9460
rect 17696 8906 17724 9454
rect 17880 9178 17908 10066
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17684 8900 17736 8906
rect 17684 8842 17736 8848
rect 17224 8560 17276 8566
rect 17224 8502 17276 8508
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17408 7336 17460 7342
rect 17408 7278 17460 7284
rect 17420 6866 17448 7278
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 14844 800 14872 2246
rect 16132 800 16160 2382
rect 17052 2106 17080 2790
rect 17512 2650 17540 7822
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17604 6458 17632 6734
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17788 3058 17816 8910
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 17500 2644 17552 2650
rect 17500 2586 17552 2592
rect 17880 2446 17908 7686
rect 18340 7478 18368 20742
rect 18432 17542 18460 21286
rect 18708 18358 18736 27338
rect 18972 27328 19024 27334
rect 18972 27270 19024 27276
rect 18984 26353 19012 27270
rect 19076 26382 19104 29158
rect 19340 29096 19392 29102
rect 19340 29038 19392 29044
rect 19248 28484 19300 28490
rect 19248 28426 19300 28432
rect 19156 28416 19208 28422
rect 19156 28358 19208 28364
rect 19064 26376 19116 26382
rect 18970 26344 19026 26353
rect 19064 26318 19116 26324
rect 18970 26279 19026 26288
rect 18880 26240 18932 26246
rect 18880 26182 18932 26188
rect 18788 25288 18840 25294
rect 18788 25230 18840 25236
rect 18800 24970 18828 25230
rect 18892 25158 18920 26182
rect 18880 25152 18932 25158
rect 18984 25140 19012 26279
rect 19168 25974 19196 28358
rect 19260 28082 19288 28426
rect 19248 28076 19300 28082
rect 19248 28018 19300 28024
rect 19248 26376 19300 26382
rect 19248 26318 19300 26324
rect 19156 25968 19208 25974
rect 19156 25910 19208 25916
rect 19154 25800 19210 25809
rect 19154 25735 19210 25744
rect 18984 25112 19104 25140
rect 18880 25094 18932 25100
rect 18800 24942 19012 24970
rect 18800 22094 18828 24942
rect 18984 24886 19012 24942
rect 18972 24880 19024 24886
rect 18972 24822 19024 24828
rect 18880 24812 18932 24818
rect 18880 24754 18932 24760
rect 18892 24274 18920 24754
rect 18880 24268 18932 24274
rect 18880 24210 18932 24216
rect 18892 23100 18920 24210
rect 18972 23112 19024 23118
rect 18892 23072 18972 23100
rect 18972 23054 19024 23060
rect 18984 22642 19012 23054
rect 18972 22636 19024 22642
rect 18972 22578 19024 22584
rect 18800 22066 18920 22094
rect 18892 21486 18920 22066
rect 18984 22030 19012 22578
rect 19076 22098 19104 25112
rect 19168 23730 19196 25735
rect 19156 23724 19208 23730
rect 19156 23666 19208 23672
rect 19156 22568 19208 22574
rect 19156 22510 19208 22516
rect 19168 22137 19196 22510
rect 19154 22128 19210 22137
rect 19064 22092 19116 22098
rect 19154 22063 19210 22072
rect 19064 22034 19116 22040
rect 18972 22024 19024 22030
rect 18972 21966 19024 21972
rect 18984 21554 19012 21966
rect 18972 21548 19024 21554
rect 18972 21490 19024 21496
rect 19260 21486 19288 26318
rect 19352 25498 19380 29038
rect 19444 27112 19472 29192
rect 19720 29170 19748 29260
rect 19708 29164 19760 29170
rect 19996 29152 20024 29271
rect 19708 29106 19760 29112
rect 19812 29124 20024 29152
rect 19522 29064 19578 29073
rect 19522 28999 19578 29008
rect 19708 29028 19760 29034
rect 19536 28558 19564 28999
rect 19812 29016 19840 29124
rect 20088 29050 20116 30330
rect 20260 29640 20312 29646
rect 20260 29582 20312 29588
rect 20272 29481 20300 29582
rect 20258 29472 20314 29481
rect 20258 29407 20314 29416
rect 20350 29336 20406 29345
rect 20350 29271 20406 29280
rect 20260 29232 20312 29238
rect 20260 29174 20312 29180
rect 20272 29102 20300 29174
rect 19760 28988 19840 29016
rect 19996 29022 20116 29050
rect 20260 29096 20312 29102
rect 20260 29038 20312 29044
rect 20168 29028 20220 29034
rect 19708 28970 19760 28976
rect 19524 28552 19576 28558
rect 19524 28494 19576 28500
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19798 27432 19854 27441
rect 19798 27367 19800 27376
rect 19852 27367 19854 27376
rect 19800 27338 19852 27344
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19444 27084 19564 27112
rect 19430 27024 19486 27033
rect 19430 26959 19432 26968
rect 19484 26959 19486 26968
rect 19432 26930 19484 26936
rect 19536 26518 19564 27084
rect 19996 26994 20024 29022
rect 20168 28970 20220 28976
rect 20076 28960 20128 28966
rect 20076 28902 20128 28908
rect 20088 28801 20116 28902
rect 20074 28792 20130 28801
rect 20074 28727 20130 28736
rect 20180 28642 20208 28970
rect 20364 28762 20392 29271
rect 20352 28756 20404 28762
rect 20352 28698 20404 28704
rect 20088 28614 20208 28642
rect 19984 26988 20036 26994
rect 19984 26930 20036 26936
rect 19996 26897 20024 26930
rect 19982 26888 20038 26897
rect 19982 26823 20038 26832
rect 19984 26784 20036 26790
rect 19984 26726 20036 26732
rect 19432 26512 19484 26518
rect 19432 26454 19484 26460
rect 19524 26512 19576 26518
rect 19524 26454 19576 26460
rect 19444 25956 19472 26454
rect 19536 26314 19564 26454
rect 19524 26308 19576 26314
rect 19524 26250 19576 26256
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19444 25928 19564 25956
rect 19432 25696 19484 25702
rect 19432 25638 19484 25644
rect 19340 25492 19392 25498
rect 19340 25434 19392 25440
rect 19340 25288 19392 25294
rect 19340 25230 19392 25236
rect 19352 24274 19380 25230
rect 19444 24274 19472 25638
rect 19536 25498 19564 25928
rect 19524 25492 19576 25498
rect 19524 25434 19576 25440
rect 19996 25294 20024 26726
rect 20088 25480 20116 28614
rect 20168 28552 20220 28558
rect 20168 28494 20220 28500
rect 20180 28082 20208 28494
rect 20168 28076 20220 28082
rect 20168 28018 20220 28024
rect 20180 26994 20208 28018
rect 20168 26988 20220 26994
rect 20168 26930 20220 26936
rect 20180 25906 20208 26930
rect 20456 26874 20484 33408
rect 20534 33008 20590 33017
rect 20534 32943 20536 32952
rect 20588 32943 20590 32952
rect 20536 32914 20588 32920
rect 20536 32836 20588 32842
rect 20536 32778 20588 32784
rect 20548 31822 20576 32778
rect 20640 32570 20668 33934
rect 20628 32564 20680 32570
rect 20628 32506 20680 32512
rect 20536 31816 20588 31822
rect 20536 31758 20588 31764
rect 20732 31754 20760 34410
rect 20824 32230 20852 35702
rect 20916 35562 20944 36654
rect 20996 36576 21048 36582
rect 20996 36518 21048 36524
rect 20904 35556 20956 35562
rect 20904 35498 20956 35504
rect 20902 35184 20958 35193
rect 20902 35119 20958 35128
rect 20916 34542 20944 35119
rect 20904 34536 20956 34542
rect 20904 34478 20956 34484
rect 20904 33856 20956 33862
rect 20904 33798 20956 33804
rect 20812 32224 20864 32230
rect 20812 32166 20864 32172
rect 20732 31726 20852 31754
rect 20720 31476 20772 31482
rect 20720 31418 20772 31424
rect 20732 31278 20760 31418
rect 20720 31272 20772 31278
rect 20720 31214 20772 31220
rect 20536 31136 20588 31142
rect 20536 31078 20588 31084
rect 20548 30598 20576 31078
rect 20626 30832 20682 30841
rect 20626 30767 20682 30776
rect 20536 30592 20588 30598
rect 20536 30534 20588 30540
rect 20640 29714 20668 30767
rect 20720 30728 20772 30734
rect 20720 30670 20772 30676
rect 20628 29708 20680 29714
rect 20628 29650 20680 29656
rect 20534 28656 20590 28665
rect 20534 28591 20590 28600
rect 20548 28490 20576 28591
rect 20536 28484 20588 28490
rect 20536 28426 20588 28432
rect 20628 27872 20680 27878
rect 20628 27814 20680 27820
rect 20640 27674 20668 27814
rect 20628 27668 20680 27674
rect 20628 27610 20680 27616
rect 20628 27464 20680 27470
rect 20628 27406 20680 27412
rect 20536 27396 20588 27402
rect 20536 27338 20588 27344
rect 20272 26846 20484 26874
rect 20168 25900 20220 25906
rect 20168 25842 20220 25848
rect 20088 25452 20208 25480
rect 20076 25356 20128 25362
rect 20076 25298 20128 25304
rect 19984 25288 20036 25294
rect 19984 25230 20036 25236
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19982 24848 20038 24857
rect 19982 24783 19984 24792
rect 20036 24783 20038 24792
rect 19984 24754 20036 24760
rect 19340 24268 19392 24274
rect 19340 24210 19392 24216
rect 19432 24268 19484 24274
rect 19432 24210 19484 24216
rect 19432 24132 19484 24138
rect 19432 24074 19484 24080
rect 19340 22432 19392 22438
rect 19340 22374 19392 22380
rect 18880 21480 18932 21486
rect 18880 21422 18932 21428
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 19248 21480 19300 21486
rect 19248 21422 19300 21428
rect 18696 18352 18748 18358
rect 18696 18294 18748 18300
rect 18604 18216 18656 18222
rect 18604 18158 18656 18164
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18420 16040 18472 16046
rect 18420 15982 18472 15988
rect 18432 12374 18460 15982
rect 18616 12442 18644 18158
rect 19076 16726 19104 21422
rect 19260 18442 19288 21422
rect 19352 18630 19380 22374
rect 19340 18624 19392 18630
rect 19340 18566 19392 18572
rect 19260 18414 19380 18442
rect 19156 18080 19208 18086
rect 19156 18022 19208 18028
rect 19064 16720 19116 16726
rect 19064 16662 19116 16668
rect 18970 16144 19026 16153
rect 18970 16079 19026 16088
rect 18788 15632 18840 15638
rect 18788 15574 18840 15580
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 18708 14822 18736 15098
rect 18800 15026 18828 15574
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18984 12986 19012 16079
rect 19064 14952 19116 14958
rect 19064 14894 19116 14900
rect 19076 14006 19104 14894
rect 19064 14000 19116 14006
rect 19064 13942 19116 13948
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 18604 12436 18656 12442
rect 18604 12378 18656 12384
rect 18420 12368 18472 12374
rect 18420 12310 18472 12316
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18708 9926 18736 10610
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 18696 9920 18748 9926
rect 18696 9862 18748 9868
rect 19076 9722 19104 10542
rect 19064 9716 19116 9722
rect 19064 9658 19116 9664
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 18328 7472 18380 7478
rect 18328 7414 18380 7420
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 18248 6866 18276 7278
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 18524 4078 18552 5102
rect 18512 4072 18564 4078
rect 18512 4014 18564 4020
rect 18616 2514 18644 9522
rect 19076 8974 19104 9658
rect 19064 8968 19116 8974
rect 19064 8910 19116 8916
rect 19168 8634 19196 18022
rect 19352 15162 19380 18414
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19246 14512 19302 14521
rect 19246 14447 19248 14456
rect 19300 14447 19302 14456
rect 19248 14418 19300 14424
rect 19352 13870 19380 14894
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19248 12368 19300 12374
rect 19248 12310 19300 12316
rect 19260 9994 19288 12310
rect 19352 11898 19380 13806
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19444 11778 19472 24074
rect 19984 24064 20036 24070
rect 19984 24006 20036 24012
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19616 22568 19668 22574
rect 19616 22510 19668 22516
rect 19628 22166 19656 22510
rect 19996 22506 20024 24006
rect 19984 22500 20036 22506
rect 19984 22442 20036 22448
rect 19616 22160 19668 22166
rect 19616 22102 19668 22108
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19708 21344 19760 21350
rect 19708 21286 19760 21292
rect 19720 20874 19748 21286
rect 19708 20868 19760 20874
rect 19708 20810 19760 20816
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19982 20496 20038 20505
rect 19982 20431 20038 20440
rect 19996 20058 20024 20431
rect 19984 20052 20036 20058
rect 19984 19994 20036 20000
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19996 19378 20024 19994
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 19708 19236 19760 19242
rect 19708 19178 19760 19184
rect 19524 19168 19576 19174
rect 19524 19110 19576 19116
rect 19536 18698 19564 19110
rect 19524 18692 19576 18698
rect 19524 18634 19576 18640
rect 19720 18630 19748 19178
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 19708 18624 19760 18630
rect 19708 18566 19760 18572
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19892 18352 19944 18358
rect 19890 18320 19892 18329
rect 19944 18320 19946 18329
rect 19890 18255 19946 18264
rect 19890 18184 19946 18193
rect 19890 18119 19892 18128
rect 19944 18119 19946 18128
rect 19892 18090 19944 18096
rect 19892 17808 19944 17814
rect 19890 17776 19892 17785
rect 19944 17776 19946 17785
rect 19996 17746 20024 18906
rect 20088 18850 20116 25298
rect 20180 24818 20208 25452
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20168 23792 20220 23798
rect 20168 23734 20220 23740
rect 20180 23594 20208 23734
rect 20168 23588 20220 23594
rect 20168 23530 20220 23536
rect 20168 22432 20220 22438
rect 20168 22374 20220 22380
rect 20180 21010 20208 22374
rect 20272 21962 20300 26846
rect 20352 26580 20404 26586
rect 20352 26522 20404 26528
rect 20364 23526 20392 26522
rect 20548 26314 20576 27338
rect 20536 26308 20588 26314
rect 20536 26250 20588 26256
rect 20536 25492 20588 25498
rect 20536 25434 20588 25440
rect 20444 25288 20496 25294
rect 20444 25230 20496 25236
rect 20352 23520 20404 23526
rect 20352 23462 20404 23468
rect 20352 23112 20404 23118
rect 20352 23054 20404 23060
rect 20364 22098 20392 23054
rect 20352 22092 20404 22098
rect 20352 22034 20404 22040
rect 20260 21956 20312 21962
rect 20260 21898 20312 21904
rect 20168 21004 20220 21010
rect 20168 20946 20220 20952
rect 20272 19530 20300 21898
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20364 20466 20392 21490
rect 20456 20602 20484 25230
rect 20548 24614 20576 25434
rect 20640 25294 20668 27406
rect 20732 25294 20760 30670
rect 20824 30326 20852 31726
rect 20916 31385 20944 33798
rect 20902 31376 20958 31385
rect 20902 31311 20958 31320
rect 21008 31210 21036 36518
rect 21100 36174 21128 36722
rect 21180 36576 21232 36582
rect 21180 36518 21232 36524
rect 21192 36310 21220 36518
rect 21180 36304 21232 36310
rect 21180 36246 21232 36252
rect 21088 36168 21140 36174
rect 21376 36145 21404 37606
rect 21456 37256 21508 37262
rect 21454 37224 21456 37233
rect 21928 37244 21956 39200
rect 23216 37262 23244 39200
rect 24032 37460 24084 37466
rect 24032 37402 24084 37408
rect 23664 37324 23716 37330
rect 23664 37266 23716 37272
rect 22836 37256 22888 37262
rect 21508 37224 21510 37233
rect 21928 37216 22140 37244
rect 21454 37159 21510 37168
rect 21456 37120 21508 37126
rect 21456 37062 21508 37068
rect 21916 37120 21968 37126
rect 21916 37062 21968 37068
rect 22008 37120 22060 37126
rect 22008 37062 22060 37068
rect 21468 36786 21496 37062
rect 21732 36916 21784 36922
rect 21732 36858 21784 36864
rect 21824 36916 21876 36922
rect 21824 36858 21876 36864
rect 21456 36780 21508 36786
rect 21456 36722 21508 36728
rect 21548 36780 21600 36786
rect 21548 36722 21600 36728
rect 21088 36110 21140 36116
rect 21362 36136 21418 36145
rect 21100 34354 21128 36110
rect 21362 36071 21364 36080
rect 21416 36071 21418 36080
rect 21364 36042 21416 36048
rect 21376 36011 21404 36042
rect 21270 35592 21326 35601
rect 21270 35527 21272 35536
rect 21324 35527 21326 35536
rect 21272 35498 21324 35504
rect 21180 35284 21232 35290
rect 21180 35226 21232 35232
rect 21192 34474 21220 35226
rect 21272 34944 21324 34950
rect 21272 34886 21324 34892
rect 21284 34513 21312 34886
rect 21270 34504 21326 34513
rect 21180 34468 21232 34474
rect 21270 34439 21326 34448
rect 21180 34410 21232 34416
rect 21272 34400 21324 34406
rect 21100 34326 21220 34354
rect 21272 34342 21324 34348
rect 21088 33992 21140 33998
rect 21088 33934 21140 33940
rect 21100 33386 21128 33934
rect 21088 33380 21140 33386
rect 21088 33322 21140 33328
rect 21088 32768 21140 32774
rect 21088 32710 21140 32716
rect 21100 32230 21128 32710
rect 21088 32224 21140 32230
rect 21088 32166 21140 32172
rect 21192 32042 21220 34326
rect 21100 32014 21220 32042
rect 20996 31204 21048 31210
rect 20996 31146 21048 31152
rect 21100 30734 21128 32014
rect 21088 30728 21140 30734
rect 21088 30670 21140 30676
rect 21180 30660 21232 30666
rect 21180 30602 21232 30608
rect 20996 30592 21048 30598
rect 20996 30534 21048 30540
rect 20812 30320 20864 30326
rect 20812 30262 20864 30268
rect 20812 30048 20864 30054
rect 20812 29990 20864 29996
rect 20904 30048 20956 30054
rect 20904 29990 20956 29996
rect 20824 26466 20852 29990
rect 20916 29850 20944 29990
rect 20904 29844 20956 29850
rect 20904 29786 20956 29792
rect 21008 29730 21036 30534
rect 20916 29702 21036 29730
rect 20916 28529 20944 29702
rect 21192 29646 21220 30602
rect 21284 30258 21312 34342
rect 21456 32972 21508 32978
rect 21456 32914 21508 32920
rect 21468 31346 21496 32914
rect 21456 31340 21508 31346
rect 21456 31282 21508 31288
rect 21364 30388 21416 30394
rect 21364 30330 21416 30336
rect 21272 30252 21324 30258
rect 21272 30194 21324 30200
rect 20996 29640 21048 29646
rect 20996 29582 21048 29588
rect 21180 29640 21232 29646
rect 21180 29582 21232 29588
rect 20902 28520 20958 28529
rect 20902 28455 20958 28464
rect 21008 28218 21036 29582
rect 21272 29232 21324 29238
rect 21272 29174 21324 29180
rect 21086 28928 21142 28937
rect 21086 28863 21142 28872
rect 21100 28422 21128 28863
rect 21180 28552 21232 28558
rect 21180 28494 21232 28500
rect 21088 28416 21140 28422
rect 21088 28358 21140 28364
rect 21192 28234 21220 28494
rect 20996 28212 21048 28218
rect 20996 28154 21048 28160
rect 21100 28206 21220 28234
rect 21284 28218 21312 29174
rect 21272 28212 21324 28218
rect 21100 28014 21128 28206
rect 21272 28154 21324 28160
rect 21180 28076 21232 28082
rect 21180 28018 21232 28024
rect 21088 28008 21140 28014
rect 21088 27950 21140 27956
rect 20904 27668 20956 27674
rect 20904 27610 20956 27616
rect 20916 27577 20944 27610
rect 20902 27568 20958 27577
rect 20902 27503 20958 27512
rect 20904 27328 20956 27334
rect 20904 27270 20956 27276
rect 20916 27130 20944 27270
rect 20904 27124 20956 27130
rect 20904 27066 20956 27072
rect 21088 26852 21140 26858
rect 21088 26794 21140 26800
rect 21100 26586 21128 26794
rect 21088 26580 21140 26586
rect 21088 26522 21140 26528
rect 20824 26438 20944 26466
rect 20812 26376 20864 26382
rect 20812 26318 20864 26324
rect 20824 25838 20852 26318
rect 20812 25832 20864 25838
rect 20812 25774 20864 25780
rect 20628 25288 20680 25294
rect 20628 25230 20680 25236
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20720 25152 20772 25158
rect 20720 25094 20772 25100
rect 20626 24984 20682 24993
rect 20626 24919 20682 24928
rect 20640 24818 20668 24919
rect 20628 24812 20680 24818
rect 20628 24754 20680 24760
rect 20536 24608 20588 24614
rect 20536 24550 20588 24556
rect 20628 24132 20680 24138
rect 20628 24074 20680 24080
rect 20536 23248 20588 23254
rect 20536 23190 20588 23196
rect 20548 22574 20576 23190
rect 20640 22710 20668 24074
rect 20732 23322 20760 25094
rect 20916 24834 20944 26438
rect 21086 26344 21142 26353
rect 21086 26279 21088 26288
rect 21140 26279 21142 26288
rect 21088 26250 21140 26256
rect 21192 26042 21220 28018
rect 21272 27328 21324 27334
rect 21272 27270 21324 27276
rect 21284 26450 21312 27270
rect 21272 26444 21324 26450
rect 21272 26386 21324 26392
rect 21180 26036 21232 26042
rect 21180 25978 21232 25984
rect 21376 25906 21404 30330
rect 21560 29510 21588 36722
rect 21640 36304 21692 36310
rect 21640 36246 21692 36252
rect 21652 36106 21680 36246
rect 21640 36100 21692 36106
rect 21640 36042 21692 36048
rect 21652 35698 21680 36042
rect 21744 36038 21772 36858
rect 21836 36530 21864 36858
rect 21928 36802 21956 37062
rect 22020 36922 22048 37062
rect 22112 36922 22140 37216
rect 22836 37198 22888 37204
rect 23204 37256 23256 37262
rect 23204 37198 23256 37204
rect 22008 36916 22060 36922
rect 22008 36858 22060 36864
rect 22100 36916 22152 36922
rect 22100 36858 22152 36864
rect 22744 36848 22796 36854
rect 21928 36774 22048 36802
rect 22744 36790 22796 36796
rect 22020 36768 22048 36774
rect 22100 36780 22152 36786
rect 22020 36740 22100 36768
rect 22100 36722 22152 36728
rect 22468 36576 22520 36582
rect 21836 36502 21956 36530
rect 22468 36518 22520 36524
rect 21822 36408 21878 36417
rect 21822 36343 21878 36352
rect 21732 36032 21784 36038
rect 21732 35974 21784 35980
rect 21836 35698 21864 36343
rect 21640 35692 21692 35698
rect 21640 35634 21692 35640
rect 21824 35692 21876 35698
rect 21824 35634 21876 35640
rect 21928 35034 21956 36502
rect 22098 36272 22154 36281
rect 22098 36207 22154 36216
rect 22008 35828 22060 35834
rect 22008 35770 22060 35776
rect 21836 35006 21956 35034
rect 21836 33318 21864 35006
rect 21916 34944 21968 34950
rect 21916 34886 21968 34892
rect 21824 33312 21876 33318
rect 21824 33254 21876 33260
rect 21640 30796 21692 30802
rect 21640 30738 21692 30744
rect 21652 30122 21680 30738
rect 21732 30660 21784 30666
rect 21732 30602 21784 30608
rect 21640 30116 21692 30122
rect 21640 30058 21692 30064
rect 21744 29850 21772 30602
rect 21732 29844 21784 29850
rect 21732 29786 21784 29792
rect 21640 29640 21692 29646
rect 21640 29582 21692 29588
rect 21548 29504 21600 29510
rect 21548 29446 21600 29452
rect 21652 28665 21680 29582
rect 21836 28665 21864 33254
rect 21928 32201 21956 34886
rect 22020 34406 22048 35770
rect 22112 34746 22140 36207
rect 22284 36100 22336 36106
rect 22284 36042 22336 36048
rect 22192 35760 22244 35766
rect 22192 35702 22244 35708
rect 22100 34740 22152 34746
rect 22100 34682 22152 34688
rect 22008 34400 22060 34406
rect 22008 34342 22060 34348
rect 22204 33590 22232 35702
rect 22296 34610 22324 36042
rect 22376 35488 22428 35494
rect 22376 35430 22428 35436
rect 22284 34604 22336 34610
rect 22284 34546 22336 34552
rect 22192 33584 22244 33590
rect 22192 33526 22244 33532
rect 22006 33008 22062 33017
rect 22006 32943 22062 32952
rect 22020 32434 22048 32943
rect 22192 32564 22244 32570
rect 22192 32506 22244 32512
rect 22008 32428 22060 32434
rect 22008 32370 22060 32376
rect 21914 32192 21970 32201
rect 21914 32127 21970 32136
rect 22008 31340 22060 31346
rect 22008 31282 22060 31288
rect 22020 29714 22048 31282
rect 22100 30796 22152 30802
rect 22100 30738 22152 30744
rect 22008 29708 22060 29714
rect 22008 29650 22060 29656
rect 21916 29572 21968 29578
rect 21916 29514 21968 29520
rect 21928 29306 21956 29514
rect 21916 29300 21968 29306
rect 21916 29242 21968 29248
rect 22112 28778 22140 30738
rect 22204 30258 22232 32506
rect 22282 30696 22338 30705
rect 22282 30631 22338 30640
rect 22296 30258 22324 30631
rect 22192 30252 22244 30258
rect 22192 30194 22244 30200
rect 22284 30252 22336 30258
rect 22284 30194 22336 30200
rect 22204 29073 22232 30194
rect 22388 29170 22416 35430
rect 22480 32366 22508 36518
rect 22756 36242 22784 36790
rect 22560 36236 22612 36242
rect 22560 36178 22612 36184
rect 22744 36236 22796 36242
rect 22744 36178 22796 36184
rect 22572 35222 22600 36178
rect 22652 35760 22704 35766
rect 22652 35702 22704 35708
rect 22560 35216 22612 35222
rect 22560 35158 22612 35164
rect 22560 35012 22612 35018
rect 22560 34954 22612 34960
rect 22468 32360 22520 32366
rect 22468 32302 22520 32308
rect 22572 31142 22600 34954
rect 22560 31136 22612 31142
rect 22560 31078 22612 31084
rect 22466 29200 22522 29209
rect 22376 29164 22428 29170
rect 22466 29135 22522 29144
rect 22376 29106 22428 29112
rect 22190 29064 22246 29073
rect 22190 28999 22246 29008
rect 22112 28750 22232 28778
rect 21638 28656 21694 28665
rect 21638 28591 21694 28600
rect 21822 28656 21878 28665
rect 21822 28591 21878 28600
rect 21732 28552 21784 28558
rect 21732 28494 21784 28500
rect 21916 28552 21968 28558
rect 21916 28494 21968 28500
rect 21454 27704 21510 27713
rect 21454 27639 21510 27648
rect 21468 26246 21496 27639
rect 21640 27464 21692 27470
rect 21640 27406 21692 27412
rect 21652 26994 21680 27406
rect 21744 27130 21772 28494
rect 21928 28257 21956 28494
rect 21914 28248 21970 28257
rect 21914 28183 21970 28192
rect 22204 28098 22232 28750
rect 22284 28416 22336 28422
rect 22284 28358 22336 28364
rect 22376 28416 22428 28422
rect 22376 28358 22428 28364
rect 22296 28218 22324 28358
rect 22284 28212 22336 28218
rect 22284 28154 22336 28160
rect 22204 28070 22324 28098
rect 21824 28008 21876 28014
rect 21824 27950 21876 27956
rect 21732 27124 21784 27130
rect 21732 27066 21784 27072
rect 21640 26988 21692 26994
rect 21640 26930 21692 26936
rect 21456 26240 21508 26246
rect 21456 26182 21508 26188
rect 21638 25936 21694 25945
rect 21180 25900 21232 25906
rect 21364 25900 21416 25906
rect 21232 25860 21312 25888
rect 21180 25842 21232 25848
rect 20996 25764 21048 25770
rect 20996 25706 21048 25712
rect 20824 24806 20944 24834
rect 21008 24818 21036 25706
rect 20996 24812 21048 24818
rect 20824 24750 20852 24806
rect 20996 24754 21048 24760
rect 20812 24744 20864 24750
rect 20812 24686 20864 24692
rect 20994 24576 21050 24585
rect 20994 24511 21050 24520
rect 20812 23724 20864 23730
rect 20812 23666 20864 23672
rect 20720 23316 20772 23322
rect 20720 23258 20772 23264
rect 20628 22704 20680 22710
rect 20628 22646 20680 22652
rect 20824 22642 20852 23666
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 21008 22574 21036 24511
rect 20536 22568 20588 22574
rect 20536 22510 20588 22516
rect 20996 22568 21048 22574
rect 20996 22510 21048 22516
rect 20534 22264 20590 22273
rect 20534 22199 20590 22208
rect 20548 22030 20576 22199
rect 20812 22092 20864 22098
rect 20812 22034 20864 22040
rect 20536 22024 20588 22030
rect 20536 21966 20588 21972
rect 20548 21554 20576 21966
rect 20628 21888 20680 21894
rect 20628 21830 20680 21836
rect 20536 21548 20588 21554
rect 20536 21490 20588 21496
rect 20536 21004 20588 21010
rect 20536 20946 20588 20952
rect 20444 20596 20496 20602
rect 20444 20538 20496 20544
rect 20352 20460 20404 20466
rect 20352 20402 20404 20408
rect 20364 19718 20392 20402
rect 20352 19712 20404 19718
rect 20352 19654 20404 19660
rect 20272 19502 20392 19530
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 20088 18822 20208 18850
rect 20076 18692 20128 18698
rect 20076 18634 20128 18640
rect 19890 17711 19946 17720
rect 19984 17740 20036 17746
rect 19984 17682 20036 17688
rect 19614 17640 19670 17649
rect 19892 17604 19944 17610
rect 19614 17575 19616 17584
rect 19668 17575 19670 17584
rect 19616 17546 19668 17552
rect 19812 17564 19892 17592
rect 19708 17536 19760 17542
rect 19812 17524 19840 17564
rect 19892 17546 19944 17552
rect 19760 17496 19840 17524
rect 19708 17478 19760 17484
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19996 16114 20024 17682
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 20088 15994 20116 18634
rect 20180 16250 20208 18822
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 19904 15966 20116 15994
rect 19904 15502 19932 15966
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 19984 15428 20036 15434
rect 19984 15370 20036 15376
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19616 14884 19668 14890
rect 19616 14826 19668 14832
rect 19628 14346 19656 14826
rect 19616 14340 19668 14346
rect 19616 14282 19668 14288
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19892 14000 19944 14006
rect 19892 13942 19944 13948
rect 19904 13802 19932 13942
rect 19892 13796 19944 13802
rect 19892 13738 19944 13744
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 19352 11750 19472 11778
rect 19248 9988 19300 9994
rect 19248 9930 19300 9936
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19168 7478 19196 8570
rect 19156 7472 19208 7478
rect 19156 7414 19208 7420
rect 19352 6662 19380 11750
rect 19536 11676 19564 11834
rect 19444 11648 19564 11676
rect 19444 10606 19472 11648
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19432 9648 19484 9654
rect 19430 9616 19432 9625
rect 19484 9616 19486 9625
rect 19430 9551 19486 9560
rect 19432 9512 19484 9518
rect 19996 9466 20024 15370
rect 20168 14612 20220 14618
rect 20168 14554 20220 14560
rect 20180 14414 20208 14554
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 20088 12170 20116 12582
rect 20076 12164 20128 12170
rect 20076 12106 20128 12112
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 19432 9454 19484 9460
rect 19444 7750 19472 9454
rect 19720 9450 20024 9466
rect 19708 9444 20024 9450
rect 19760 9438 20024 9444
rect 19708 9386 19760 9392
rect 19800 9376 19852 9382
rect 19800 9318 19852 9324
rect 19812 9178 19840 9318
rect 19800 9172 19852 9178
rect 19800 9114 19852 9120
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 20088 8498 20116 10406
rect 20166 9616 20222 9625
rect 20166 9551 20168 9560
rect 20220 9551 20222 9560
rect 20168 9522 20220 9528
rect 20272 8838 20300 19110
rect 20364 15910 20392 19502
rect 20548 18698 20576 20946
rect 20640 20874 20668 21830
rect 20824 21690 20852 22034
rect 21088 21956 21140 21962
rect 21088 21898 21140 21904
rect 21100 21690 21128 21898
rect 20812 21684 20864 21690
rect 20812 21626 20864 21632
rect 21088 21684 21140 21690
rect 21088 21626 21140 21632
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20732 21078 20760 21422
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20720 21072 20772 21078
rect 20720 21014 20772 21020
rect 20628 20868 20680 20874
rect 20628 20810 20680 20816
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 20640 20398 20668 20538
rect 20628 20392 20680 20398
rect 20628 20334 20680 20340
rect 20536 18692 20588 18698
rect 20536 18634 20588 18640
rect 20444 17604 20496 17610
rect 20444 17546 20496 17552
rect 20456 16998 20484 17546
rect 20444 16992 20496 16998
rect 20444 16934 20496 16940
rect 20456 16590 20484 16934
rect 20640 16658 20668 20334
rect 20720 19236 20772 19242
rect 20720 19178 20772 19184
rect 20628 16652 20680 16658
rect 20628 16594 20680 16600
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20732 16182 20760 19178
rect 20824 16454 20852 21286
rect 20812 16448 20864 16454
rect 20812 16390 20864 16396
rect 20720 16176 20772 16182
rect 20720 16118 20772 16124
rect 20352 15904 20404 15910
rect 20352 15846 20404 15852
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20732 15162 20760 15846
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20916 15094 20944 21286
rect 21284 21026 21312 25860
rect 21416 25860 21588 25888
rect 21638 25871 21640 25880
rect 21364 25842 21416 25848
rect 21364 25696 21416 25702
rect 21364 25638 21416 25644
rect 21376 24682 21404 25638
rect 21456 25288 21508 25294
rect 21456 25230 21508 25236
rect 21364 24676 21416 24682
rect 21364 24618 21416 24624
rect 21468 23798 21496 25230
rect 21560 24857 21588 25860
rect 21692 25871 21694 25880
rect 21640 25842 21692 25848
rect 21546 24848 21602 24857
rect 21546 24783 21602 24792
rect 21560 24206 21588 24783
rect 21730 24712 21786 24721
rect 21640 24676 21692 24682
rect 21730 24647 21786 24656
rect 21640 24618 21692 24624
rect 21548 24200 21600 24206
rect 21548 24142 21600 24148
rect 21456 23792 21508 23798
rect 21456 23734 21508 23740
rect 21560 23118 21588 24142
rect 21652 23662 21680 24618
rect 21744 24410 21772 24647
rect 21732 24404 21784 24410
rect 21732 24346 21784 24352
rect 21730 24168 21786 24177
rect 21730 24103 21786 24112
rect 21744 24070 21772 24103
rect 21732 24064 21784 24070
rect 21732 24006 21784 24012
rect 21640 23656 21692 23662
rect 21836 23633 21864 27950
rect 22192 27600 22244 27606
rect 21914 27568 21970 27577
rect 21914 27503 21916 27512
rect 21968 27503 21970 27512
rect 22190 27568 22192 27577
rect 22244 27568 22246 27577
rect 22190 27503 22246 27512
rect 21916 27474 21968 27480
rect 22100 26920 22152 26926
rect 22100 26862 22152 26868
rect 22112 25888 22140 26862
rect 22192 25900 22244 25906
rect 22112 25860 22192 25888
rect 21916 24744 21968 24750
rect 21916 24686 21968 24692
rect 21928 24177 21956 24686
rect 22008 24608 22060 24614
rect 22008 24550 22060 24556
rect 22020 24342 22048 24550
rect 22008 24336 22060 24342
rect 22008 24278 22060 24284
rect 21914 24168 21970 24177
rect 21914 24103 21970 24112
rect 21640 23598 21692 23604
rect 21822 23624 21878 23633
rect 21822 23559 21878 23568
rect 22006 23488 22062 23497
rect 22006 23423 22062 23432
rect 21548 23112 21600 23118
rect 21548 23054 21600 23060
rect 21638 22128 21694 22137
rect 21364 22092 21416 22098
rect 21638 22063 21694 22072
rect 21364 22034 21416 22040
rect 21376 21690 21404 22034
rect 21364 21684 21416 21690
rect 21364 21626 21416 21632
rect 21192 20998 21312 21026
rect 21192 20942 21220 20998
rect 21180 20936 21232 20942
rect 21180 20878 21232 20884
rect 21192 20806 21220 20878
rect 21180 20800 21232 20806
rect 21180 20742 21232 20748
rect 21088 18692 21140 18698
rect 21088 18634 21140 18640
rect 20996 18352 21048 18358
rect 20996 18294 21048 18300
rect 21008 17338 21036 18294
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 21100 16658 21128 18634
rect 21192 17649 21220 20742
rect 21652 19718 21680 22063
rect 21916 20392 21968 20398
rect 21916 20334 21968 20340
rect 21928 19990 21956 20334
rect 21916 19984 21968 19990
rect 21916 19926 21968 19932
rect 21640 19712 21692 19718
rect 21640 19654 21692 19660
rect 21652 18986 21680 19654
rect 21916 19372 21968 19378
rect 21916 19314 21968 19320
rect 21560 18958 21680 18986
rect 21456 18148 21508 18154
rect 21456 18090 21508 18096
rect 21178 17640 21234 17649
rect 21178 17575 21234 17584
rect 21088 16652 21140 16658
rect 21088 16594 21140 16600
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 20996 16040 21048 16046
rect 20996 15982 21048 15988
rect 20904 15088 20956 15094
rect 20904 15030 20956 15036
rect 21008 14074 21036 15982
rect 21180 15428 21232 15434
rect 21180 15370 21232 15376
rect 21088 14952 21140 14958
rect 21088 14894 21140 14900
rect 21100 14482 21128 14894
rect 21192 14618 21220 15370
rect 21180 14612 21232 14618
rect 21180 14554 21232 14560
rect 21088 14476 21140 14482
rect 21088 14418 21140 14424
rect 21100 14074 21128 14418
rect 21284 14278 21312 16390
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21376 14521 21404 14554
rect 21362 14512 21418 14521
rect 21362 14447 21418 14456
rect 21272 14272 21324 14278
rect 21272 14214 21324 14220
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21468 13530 21496 18090
rect 21560 17678 21588 18958
rect 21640 18896 21692 18902
rect 21640 18838 21692 18844
rect 21548 17672 21600 17678
rect 21548 17614 21600 17620
rect 21652 17610 21680 18838
rect 21640 17604 21692 17610
rect 21640 17546 21692 17552
rect 21732 16652 21784 16658
rect 21732 16594 21784 16600
rect 21548 16108 21600 16114
rect 21548 16050 21600 16056
rect 21560 13938 21588 16050
rect 21548 13932 21600 13938
rect 21548 13874 21600 13880
rect 21456 13524 21508 13530
rect 21456 13466 21508 13472
rect 21640 12708 21692 12714
rect 21640 12650 21692 12656
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20536 12300 20588 12306
rect 20536 12242 20588 12248
rect 20548 11082 20576 12242
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20536 11076 20588 11082
rect 20536 11018 20588 11024
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 20548 8090 20576 11018
rect 20732 10674 20760 11698
rect 20824 11082 20852 12582
rect 20812 11076 20864 11082
rect 20812 11018 20864 11024
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 20732 10538 20760 10610
rect 20720 10532 20772 10538
rect 20720 10474 20772 10480
rect 20732 10062 20760 10474
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 20904 10464 20956 10470
rect 20904 10406 20956 10412
rect 20824 10130 20852 10406
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20732 9654 20760 9862
rect 20916 9722 20944 10406
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 20536 8084 20588 8090
rect 20536 8026 20588 8032
rect 21652 7818 21680 12650
rect 20076 7812 20128 7818
rect 20076 7754 20128 7760
rect 21548 7812 21600 7818
rect 21548 7754 21600 7760
rect 21640 7812 21692 7818
rect 21640 7754 21692 7760
rect 19432 7744 19484 7750
rect 19432 7686 19484 7692
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19432 7472 19484 7478
rect 19996 7426 20024 7686
rect 19432 7414 19484 7420
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19444 6458 19472 7414
rect 19904 7398 20024 7426
rect 19904 7342 19932 7398
rect 20088 7342 20116 7754
rect 21560 7546 21588 7754
rect 21548 7540 21600 7546
rect 21548 7482 21600 7488
rect 19892 7336 19944 7342
rect 19892 7278 19944 7284
rect 20076 7336 20128 7342
rect 20076 7278 20128 7284
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 20536 5160 20588 5166
rect 20536 5102 20588 5108
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 20548 4146 20576 5102
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 19444 2650 19472 4082
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 20732 2650 20760 6734
rect 21744 4010 21772 16594
rect 21824 16516 21876 16522
rect 21824 16458 21876 16464
rect 21836 13938 21864 16458
rect 21928 14618 21956 19314
rect 22020 18154 22048 23423
rect 22112 22438 22140 25860
rect 22192 25842 22244 25848
rect 22192 23588 22244 23594
rect 22192 23530 22244 23536
rect 22204 22794 22232 23530
rect 22296 23497 22324 28070
rect 22388 28014 22416 28358
rect 22376 28008 22428 28014
rect 22376 27950 22428 27956
rect 22480 27062 22508 29135
rect 22468 27056 22520 27062
rect 22468 26998 22520 27004
rect 22468 26920 22520 26926
rect 22468 26862 22520 26868
rect 22376 25968 22428 25974
rect 22376 25910 22428 25916
rect 22282 23488 22338 23497
rect 22282 23423 22338 23432
rect 22204 22766 22324 22794
rect 22192 22704 22244 22710
rect 22192 22646 22244 22652
rect 22100 22432 22152 22438
rect 22100 22374 22152 22380
rect 22100 22160 22152 22166
rect 22100 22102 22152 22108
rect 22112 19938 22140 22102
rect 22204 20602 22232 22646
rect 22296 22166 22324 22766
rect 22284 22160 22336 22166
rect 22284 22102 22336 22108
rect 22284 21480 22336 21486
rect 22284 21422 22336 21428
rect 22296 20806 22324 21422
rect 22388 20924 22416 25910
rect 22480 23594 22508 26862
rect 22572 25498 22600 31078
rect 22664 28762 22692 35702
rect 22744 34128 22796 34134
rect 22744 34070 22796 34076
rect 22756 33930 22784 34070
rect 22744 33924 22796 33930
rect 22744 33866 22796 33872
rect 22742 33552 22798 33561
rect 22742 33487 22744 33496
rect 22796 33487 22798 33496
rect 22744 33458 22796 33464
rect 22744 29640 22796 29646
rect 22744 29582 22796 29588
rect 22652 28756 22704 28762
rect 22652 28698 22704 28704
rect 22664 28082 22692 28698
rect 22652 28076 22704 28082
rect 22652 28018 22704 28024
rect 22560 25492 22612 25498
rect 22560 25434 22612 25440
rect 22756 24392 22784 29582
rect 22848 28098 22876 37198
rect 22928 36780 22980 36786
rect 22928 36722 22980 36728
rect 22940 36378 22968 36722
rect 23020 36576 23072 36582
rect 23020 36518 23072 36524
rect 22928 36372 22980 36378
rect 22928 36314 22980 36320
rect 23032 34066 23060 36518
rect 23480 36032 23532 36038
rect 23480 35974 23532 35980
rect 23296 35624 23348 35630
rect 23296 35566 23348 35572
rect 23308 35329 23336 35566
rect 23294 35320 23350 35329
rect 23294 35255 23350 35264
rect 23388 35216 23440 35222
rect 23388 35158 23440 35164
rect 23112 35012 23164 35018
rect 23112 34954 23164 34960
rect 23124 34921 23152 34954
rect 23110 34912 23166 34921
rect 23110 34847 23166 34856
rect 23400 34746 23428 35158
rect 23388 34740 23440 34746
rect 23388 34682 23440 34688
rect 23388 34468 23440 34474
rect 23388 34410 23440 34416
rect 23020 34060 23072 34066
rect 23020 34002 23072 34008
rect 23204 32904 23256 32910
rect 23204 32846 23256 32852
rect 23216 32502 23244 32846
rect 23204 32496 23256 32502
rect 23204 32438 23256 32444
rect 23296 32428 23348 32434
rect 23296 32370 23348 32376
rect 23020 32292 23072 32298
rect 23020 32234 23072 32240
rect 22928 31680 22980 31686
rect 22928 31622 22980 31628
rect 22940 30376 22968 31622
rect 23032 30802 23060 32234
rect 23204 31748 23256 31754
rect 23204 31690 23256 31696
rect 23110 30968 23166 30977
rect 23110 30903 23166 30912
rect 23020 30796 23072 30802
rect 23020 30738 23072 30744
rect 23124 30734 23152 30903
rect 23112 30728 23164 30734
rect 23112 30670 23164 30676
rect 22940 30348 23152 30376
rect 22928 30184 22980 30190
rect 22928 30126 22980 30132
rect 22940 29646 22968 30126
rect 22928 29640 22980 29646
rect 22928 29582 22980 29588
rect 23020 29504 23072 29510
rect 23020 29446 23072 29452
rect 23032 29238 23060 29446
rect 22928 29232 22980 29238
rect 22928 29174 22980 29180
rect 23020 29232 23072 29238
rect 23020 29174 23072 29180
rect 22940 29050 22968 29174
rect 22940 29022 23060 29050
rect 23032 28626 23060 29022
rect 23020 28620 23072 28626
rect 23020 28562 23072 28568
rect 22848 28082 23060 28098
rect 22848 28076 23072 28082
rect 22848 28070 23020 28076
rect 23020 28018 23072 28024
rect 22928 25288 22980 25294
rect 22928 25230 22980 25236
rect 22940 24682 22968 25230
rect 22928 24676 22980 24682
rect 22928 24618 22980 24624
rect 22756 24364 22968 24392
rect 22652 24336 22704 24342
rect 22652 24278 22704 24284
rect 22664 23730 22692 24278
rect 22836 24268 22888 24274
rect 22836 24210 22888 24216
rect 22652 23724 22704 23730
rect 22652 23666 22704 23672
rect 22558 23624 22614 23633
rect 22468 23588 22520 23594
rect 22558 23559 22614 23568
rect 22468 23530 22520 23536
rect 22468 22500 22520 22506
rect 22468 22442 22520 22448
rect 22480 22030 22508 22442
rect 22468 22024 22520 22030
rect 22468 21966 22520 21972
rect 22388 20896 22508 20924
rect 22284 20800 22336 20806
rect 22284 20742 22336 20748
rect 22192 20596 22244 20602
rect 22192 20538 22244 20544
rect 22112 19910 22324 19938
rect 22098 19816 22154 19825
rect 22098 19751 22154 19760
rect 22112 19174 22140 19751
rect 22192 19440 22244 19446
rect 22192 19382 22244 19388
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 22204 18970 22232 19382
rect 22192 18964 22244 18970
rect 22192 18906 22244 18912
rect 22008 18148 22060 18154
rect 22008 18090 22060 18096
rect 22296 17762 22324 19910
rect 22204 17734 22324 17762
rect 22008 16516 22060 16522
rect 22008 16458 22060 16464
rect 22020 15706 22048 16458
rect 22008 15700 22060 15706
rect 22008 15642 22060 15648
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 21824 13932 21876 13938
rect 21824 13874 21876 13880
rect 22008 13932 22060 13938
rect 22008 13874 22060 13880
rect 21916 13320 21968 13326
rect 21916 13262 21968 13268
rect 21928 11830 21956 13262
rect 21916 11824 21968 11830
rect 21916 11766 21968 11772
rect 22020 10674 22048 13874
rect 22204 13870 22232 17734
rect 22284 17604 22336 17610
rect 22284 17546 22336 17552
rect 22376 17604 22428 17610
rect 22376 17546 22428 17552
rect 22296 16640 22324 17546
rect 22388 17270 22416 17546
rect 22376 17264 22428 17270
rect 22376 17206 22428 17212
rect 22376 16652 22428 16658
rect 22296 16612 22376 16640
rect 22376 16594 22428 16600
rect 22192 13864 22244 13870
rect 22192 13806 22244 13812
rect 22388 13530 22416 16594
rect 22376 13524 22428 13530
rect 22376 13466 22428 13472
rect 22480 12850 22508 20896
rect 22572 19786 22600 23559
rect 22652 22500 22704 22506
rect 22652 22442 22704 22448
rect 22560 19780 22612 19786
rect 22560 19722 22612 19728
rect 22560 16584 22612 16590
rect 22560 16526 22612 16532
rect 22572 16250 22600 16526
rect 22560 16244 22612 16250
rect 22560 16186 22612 16192
rect 22664 13258 22692 22442
rect 22744 21412 22796 21418
rect 22744 21354 22796 21360
rect 22756 15858 22784 21354
rect 22848 15978 22876 24210
rect 22940 22094 22968 24364
rect 23032 23798 23060 28018
rect 23124 26858 23152 30348
rect 23216 30190 23244 31690
rect 23204 30184 23256 30190
rect 23204 30126 23256 30132
rect 23204 28144 23256 28150
rect 23204 28086 23256 28092
rect 23112 26852 23164 26858
rect 23112 26794 23164 26800
rect 23110 26480 23166 26489
rect 23110 26415 23166 26424
rect 23124 26382 23152 26415
rect 23112 26376 23164 26382
rect 23112 26318 23164 26324
rect 23216 24274 23244 28086
rect 23308 26330 23336 32370
rect 23400 28150 23428 34410
rect 23492 34134 23520 35974
rect 23480 34128 23532 34134
rect 23480 34070 23532 34076
rect 23572 33992 23624 33998
rect 23572 33934 23624 33940
rect 23584 33810 23612 33934
rect 23492 33782 23612 33810
rect 23492 33318 23520 33782
rect 23572 33652 23624 33658
rect 23572 33594 23624 33600
rect 23480 33312 23532 33318
rect 23480 33254 23532 33260
rect 23584 33046 23612 33594
rect 23572 33040 23624 33046
rect 23572 32982 23624 32988
rect 23572 32496 23624 32502
rect 23572 32438 23624 32444
rect 23480 31476 23532 31482
rect 23480 31418 23532 31424
rect 23388 28144 23440 28150
rect 23388 28086 23440 28092
rect 23388 27940 23440 27946
rect 23388 27882 23440 27888
rect 23400 26994 23428 27882
rect 23388 26988 23440 26994
rect 23388 26930 23440 26936
rect 23492 26874 23520 31418
rect 23584 30326 23612 32438
rect 23572 30320 23624 30326
rect 23572 30262 23624 30268
rect 23570 28656 23626 28665
rect 23570 28591 23626 28600
rect 23584 28082 23612 28591
rect 23572 28076 23624 28082
rect 23572 28018 23624 28024
rect 23572 27464 23624 27470
rect 23572 27406 23624 27412
rect 23584 27130 23612 27406
rect 23572 27124 23624 27130
rect 23572 27066 23624 27072
rect 23492 26846 23612 26874
rect 23308 26302 23428 26330
rect 23296 26240 23348 26246
rect 23296 26182 23348 26188
rect 23308 25906 23336 26182
rect 23296 25900 23348 25906
rect 23296 25842 23348 25848
rect 23204 24268 23256 24274
rect 23204 24210 23256 24216
rect 23020 23792 23072 23798
rect 23020 23734 23072 23740
rect 22940 22066 23336 22094
rect 23204 22024 23256 22030
rect 23204 21966 23256 21972
rect 23216 21622 23244 21966
rect 23204 21616 23256 21622
rect 23204 21558 23256 21564
rect 23308 21554 23336 22066
rect 23296 21548 23348 21554
rect 23296 21490 23348 21496
rect 23020 20868 23072 20874
rect 23020 20810 23072 20816
rect 23112 20868 23164 20874
rect 23112 20810 23164 20816
rect 23032 19446 23060 20810
rect 23020 19440 23072 19446
rect 23020 19382 23072 19388
rect 22928 18760 22980 18766
rect 22928 18702 22980 18708
rect 22940 18193 22968 18702
rect 22926 18184 22982 18193
rect 22926 18119 22982 18128
rect 22928 16516 22980 16522
rect 22928 16458 22980 16464
rect 22836 15972 22888 15978
rect 22836 15914 22888 15920
rect 22756 15830 22876 15858
rect 22744 14816 22796 14822
rect 22744 14758 22796 14764
rect 22756 14385 22784 14758
rect 22742 14376 22798 14385
rect 22742 14311 22798 14320
rect 22652 13252 22704 13258
rect 22652 13194 22704 13200
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22664 12306 22692 13194
rect 22848 12918 22876 15830
rect 22940 15502 22968 16458
rect 22928 15496 22980 15502
rect 22928 15438 22980 15444
rect 22928 14952 22980 14958
rect 22928 14894 22980 14900
rect 22940 14346 22968 14894
rect 22928 14340 22980 14346
rect 22928 14282 22980 14288
rect 22836 12912 22888 12918
rect 22836 12854 22888 12860
rect 22652 12300 22704 12306
rect 22652 12242 22704 12248
rect 22192 11552 22244 11558
rect 22192 11494 22244 11500
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22112 11082 22140 11290
rect 22204 11218 22232 11494
rect 22192 11212 22244 11218
rect 22192 11154 22244 11160
rect 23124 11082 23152 20810
rect 23204 19848 23256 19854
rect 23204 19790 23256 19796
rect 23216 17610 23244 19790
rect 23400 18766 23428 26302
rect 23584 20806 23612 26846
rect 23676 21570 23704 37266
rect 23756 37256 23808 37262
rect 23756 37198 23808 37204
rect 23768 31482 23796 37198
rect 24044 35018 24072 37402
rect 24504 37126 24532 39200
rect 25148 37330 25176 39200
rect 25136 37324 25188 37330
rect 25136 37266 25188 37272
rect 25872 37256 25924 37262
rect 25872 37198 25924 37204
rect 24400 37120 24452 37126
rect 24400 37062 24452 37068
rect 24492 37120 24544 37126
rect 24492 37062 24544 37068
rect 25504 37120 25556 37126
rect 25504 37062 25556 37068
rect 24412 36378 24440 37062
rect 25136 36848 25188 36854
rect 25228 36848 25280 36854
rect 25136 36790 25188 36796
rect 25226 36816 25228 36825
rect 25280 36816 25282 36825
rect 25044 36712 25096 36718
rect 25044 36654 25096 36660
rect 24400 36372 24452 36378
rect 24400 36314 24452 36320
rect 25056 36281 25084 36654
rect 25148 36650 25176 36790
rect 25226 36751 25282 36760
rect 25228 36712 25280 36718
rect 25228 36654 25280 36660
rect 25136 36644 25188 36650
rect 25136 36586 25188 36592
rect 25042 36272 25098 36281
rect 25042 36207 25098 36216
rect 25136 35760 25188 35766
rect 25136 35702 25188 35708
rect 24768 35488 24820 35494
rect 24768 35430 24820 35436
rect 24492 35216 24544 35222
rect 24492 35158 24544 35164
rect 24032 35012 24084 35018
rect 24032 34954 24084 34960
rect 24504 34610 24532 35158
rect 24780 34678 24808 35430
rect 25148 35222 25176 35702
rect 25240 35494 25268 36654
rect 25516 36242 25544 37062
rect 25884 36378 25912 37198
rect 25872 36372 25924 36378
rect 25872 36314 25924 36320
rect 25504 36236 25556 36242
rect 25504 36178 25556 36184
rect 25596 36100 25648 36106
rect 25596 36042 25648 36048
rect 25412 35760 25464 35766
rect 25410 35728 25412 35737
rect 25464 35728 25466 35737
rect 25410 35663 25466 35672
rect 25228 35488 25280 35494
rect 25228 35430 25280 35436
rect 25318 35456 25374 35465
rect 25136 35216 25188 35222
rect 25136 35158 25188 35164
rect 25136 34740 25188 34746
rect 25136 34682 25188 34688
rect 24768 34672 24820 34678
rect 24768 34614 24820 34620
rect 24952 34672 25004 34678
rect 24952 34614 25004 34620
rect 23940 34604 23992 34610
rect 23940 34546 23992 34552
rect 24492 34604 24544 34610
rect 24492 34546 24544 34552
rect 23846 34096 23902 34105
rect 23846 34031 23902 34040
rect 23860 33658 23888 34031
rect 23952 33969 23980 34546
rect 24124 34400 24176 34406
rect 24124 34342 24176 34348
rect 24032 34128 24084 34134
rect 24032 34070 24084 34076
rect 23938 33960 23994 33969
rect 23938 33895 23994 33904
rect 23848 33652 23900 33658
rect 23848 33594 23900 33600
rect 23940 33312 23992 33318
rect 23940 33254 23992 33260
rect 23848 32836 23900 32842
rect 23848 32778 23900 32784
rect 23860 31482 23888 32778
rect 23952 32366 23980 33254
rect 23940 32360 23992 32366
rect 23940 32302 23992 32308
rect 23756 31476 23808 31482
rect 23756 31418 23808 31424
rect 23848 31476 23900 31482
rect 23848 31418 23900 31424
rect 23756 31340 23808 31346
rect 23756 31282 23808 31288
rect 23848 31340 23900 31346
rect 23848 31282 23900 31288
rect 23768 30938 23796 31282
rect 23756 30932 23808 30938
rect 23756 30874 23808 30880
rect 23860 28694 23888 31282
rect 23940 30048 23992 30054
rect 23940 29990 23992 29996
rect 23952 29850 23980 29990
rect 23940 29844 23992 29850
rect 23940 29786 23992 29792
rect 23940 29096 23992 29102
rect 23940 29038 23992 29044
rect 23848 28688 23900 28694
rect 23848 28630 23900 28636
rect 23848 27056 23900 27062
rect 23848 26998 23900 27004
rect 23860 26586 23888 26998
rect 23848 26580 23900 26586
rect 23848 26522 23900 26528
rect 23952 26466 23980 29038
rect 24044 27606 24072 34070
rect 24136 33590 24164 34342
rect 24504 34066 24532 34546
rect 24492 34060 24544 34066
rect 24492 34002 24544 34008
rect 24308 33992 24360 33998
rect 24228 33952 24308 33980
rect 24124 33584 24176 33590
rect 24124 33526 24176 33532
rect 24124 31408 24176 31414
rect 24228 31396 24256 33952
rect 24308 33934 24360 33940
rect 24584 32904 24636 32910
rect 24582 32872 24584 32881
rect 24636 32872 24638 32881
rect 24582 32807 24638 32816
rect 24860 32360 24912 32366
rect 24860 32302 24912 32308
rect 24176 31368 24256 31396
rect 24124 31350 24176 31356
rect 24032 27600 24084 27606
rect 24032 27542 24084 27548
rect 24032 27124 24084 27130
rect 24032 27066 24084 27072
rect 23860 26438 23980 26466
rect 23756 26376 23808 26382
rect 23756 26318 23808 26324
rect 23768 25294 23796 26318
rect 23756 25288 23808 25294
rect 23756 25230 23808 25236
rect 23860 24682 23888 26438
rect 23940 25900 23992 25906
rect 23940 25842 23992 25848
rect 23952 24818 23980 25842
rect 23940 24812 23992 24818
rect 23940 24754 23992 24760
rect 24044 24721 24072 27066
rect 24030 24712 24086 24721
rect 23848 24676 23900 24682
rect 23848 24618 23900 24624
rect 23952 24670 24030 24698
rect 23756 22092 23808 22098
rect 23952 22094 23980 24670
rect 24030 24647 24086 24656
rect 24032 23860 24084 23866
rect 24032 23802 24084 23808
rect 23756 22034 23808 22040
rect 23860 22066 23980 22094
rect 23768 21690 23796 22034
rect 23860 22030 23888 22066
rect 23848 22024 23900 22030
rect 23848 21966 23900 21972
rect 24044 21690 24072 23802
rect 24136 23730 24164 31350
rect 24768 31136 24820 31142
rect 24768 31078 24820 31084
rect 24400 30320 24452 30326
rect 24400 30262 24452 30268
rect 24216 30184 24268 30190
rect 24216 30126 24268 30132
rect 24228 24970 24256 30126
rect 24308 30048 24360 30054
rect 24308 29990 24360 29996
rect 24320 29714 24348 29990
rect 24308 29708 24360 29714
rect 24308 29650 24360 29656
rect 24308 28008 24360 28014
rect 24308 27950 24360 27956
rect 24320 27441 24348 27950
rect 24306 27432 24362 27441
rect 24306 27367 24362 27376
rect 24412 27130 24440 30262
rect 24780 29889 24808 31078
rect 24766 29880 24822 29889
rect 24872 29850 24900 32302
rect 24964 31958 24992 34614
rect 25148 33658 25176 34682
rect 25136 33652 25188 33658
rect 25136 33594 25188 33600
rect 25044 33516 25096 33522
rect 25044 33458 25096 33464
rect 25056 32910 25084 33458
rect 25044 32904 25096 32910
rect 25044 32846 25096 32852
rect 25240 32722 25268 35430
rect 25318 35391 25374 35400
rect 25332 35086 25360 35391
rect 25608 35290 25636 36042
rect 26436 35834 26464 39200
rect 27436 37256 27488 37262
rect 27436 37198 27488 37204
rect 27448 36854 27476 37198
rect 27724 37126 27752 39200
rect 28368 37330 28396 39200
rect 29656 37330 29684 39200
rect 28356 37324 28408 37330
rect 28356 37266 28408 37272
rect 29644 37324 29696 37330
rect 29644 37266 29696 37272
rect 30944 37262 30972 39200
rect 27804 37256 27856 37262
rect 27804 37198 27856 37204
rect 30932 37256 30984 37262
rect 30932 37198 30984 37204
rect 27712 37120 27764 37126
rect 27712 37062 27764 37068
rect 27816 36922 27844 37198
rect 32232 37126 32260 39200
rect 32876 37262 32904 39200
rect 34164 37330 34192 39200
rect 35452 39114 35480 39200
rect 35544 39114 35572 39222
rect 35452 39086 35572 39114
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34152 37324 34204 37330
rect 34152 37266 34204 37272
rect 32864 37256 32916 37262
rect 32864 37198 32916 37204
rect 28540 37120 28592 37126
rect 28540 37062 28592 37068
rect 28908 37120 28960 37126
rect 28908 37062 28960 37068
rect 29828 37120 29880 37126
rect 29828 37062 29880 37068
rect 31024 37120 31076 37126
rect 31024 37062 31076 37068
rect 32220 37120 32272 37126
rect 32220 37062 32272 37068
rect 33048 37120 33100 37126
rect 35820 37108 35848 39222
rect 36082 39200 36138 39800
rect 37370 39200 37426 39800
rect 38658 39200 38714 39800
rect 39302 39200 39358 39800
rect 35900 37120 35952 37126
rect 35820 37080 35900 37108
rect 33048 37062 33100 37068
rect 35900 37062 35952 37068
rect 27804 36916 27856 36922
rect 27804 36858 27856 36864
rect 27436 36848 27488 36854
rect 27436 36790 27488 36796
rect 26976 36780 27028 36786
rect 26976 36722 27028 36728
rect 26988 36038 27016 36722
rect 27528 36712 27580 36718
rect 27528 36654 27580 36660
rect 28356 36712 28408 36718
rect 28356 36654 28408 36660
rect 27252 36644 27304 36650
rect 27252 36586 27304 36592
rect 26792 36032 26844 36038
rect 26792 35974 26844 35980
rect 26976 36032 27028 36038
rect 26976 35974 27028 35980
rect 26424 35828 26476 35834
rect 26424 35770 26476 35776
rect 25780 35556 25832 35562
rect 25780 35498 25832 35504
rect 25596 35284 25648 35290
rect 25596 35226 25648 35232
rect 25320 35080 25372 35086
rect 25320 35022 25372 35028
rect 25792 33289 25820 35498
rect 26332 35488 26384 35494
rect 26332 35430 26384 35436
rect 26344 35154 26372 35430
rect 26804 35154 26832 35974
rect 26332 35148 26384 35154
rect 26332 35090 26384 35096
rect 26792 35148 26844 35154
rect 26792 35090 26844 35096
rect 26424 35012 26476 35018
rect 26424 34954 26476 34960
rect 26436 33658 26464 34954
rect 26516 34944 26568 34950
rect 26516 34886 26568 34892
rect 26528 34746 26556 34886
rect 26516 34740 26568 34746
rect 26516 34682 26568 34688
rect 26424 33652 26476 33658
rect 26424 33594 26476 33600
rect 25964 33516 26016 33522
rect 25964 33458 26016 33464
rect 25778 33280 25834 33289
rect 25778 33215 25834 33224
rect 25504 32836 25556 32842
rect 25504 32778 25556 32784
rect 25056 32694 25268 32722
rect 24952 31952 25004 31958
rect 24952 31894 25004 31900
rect 24952 30320 25004 30326
rect 24952 30262 25004 30268
rect 24766 29815 24822 29824
rect 24860 29844 24912 29850
rect 24860 29786 24912 29792
rect 24768 29708 24820 29714
rect 24872 29696 24900 29786
rect 24820 29668 24900 29696
rect 24768 29650 24820 29656
rect 24860 29300 24912 29306
rect 24860 29242 24912 29248
rect 24492 29232 24544 29238
rect 24872 29209 24900 29242
rect 24492 29174 24544 29180
rect 24858 29200 24914 29209
rect 24400 27124 24452 27130
rect 24400 27066 24452 27072
rect 24400 26988 24452 26994
rect 24400 26930 24452 26936
rect 24412 26382 24440 26930
rect 24504 26790 24532 29174
rect 24858 29135 24914 29144
rect 24584 28688 24636 28694
rect 24584 28630 24636 28636
rect 24596 28558 24624 28630
rect 24964 28558 24992 30262
rect 25056 29170 25084 32694
rect 25136 32496 25188 32502
rect 25136 32438 25188 32444
rect 25148 32026 25176 32438
rect 25412 32292 25464 32298
rect 25412 32234 25464 32240
rect 25228 32224 25280 32230
rect 25228 32166 25280 32172
rect 25136 32020 25188 32026
rect 25136 31962 25188 31968
rect 25240 31278 25268 32166
rect 25424 31958 25452 32234
rect 25412 31952 25464 31958
rect 25412 31894 25464 31900
rect 25320 31680 25372 31686
rect 25320 31622 25372 31628
rect 25332 31414 25360 31622
rect 25320 31408 25372 31414
rect 25320 31350 25372 31356
rect 25228 31272 25280 31278
rect 25228 31214 25280 31220
rect 25044 29164 25096 29170
rect 25044 29106 25096 29112
rect 25240 29102 25268 31214
rect 25320 29708 25372 29714
rect 25320 29650 25372 29656
rect 25228 29096 25280 29102
rect 25228 29038 25280 29044
rect 24584 28552 24636 28558
rect 24584 28494 24636 28500
rect 24952 28552 25004 28558
rect 24952 28494 25004 28500
rect 25136 28552 25188 28558
rect 25136 28494 25188 28500
rect 24768 28416 24820 28422
rect 24768 28358 24820 28364
rect 24584 27464 24636 27470
rect 24584 27406 24636 27412
rect 24596 27130 24624 27406
rect 24676 27328 24728 27334
rect 24676 27270 24728 27276
rect 24584 27124 24636 27130
rect 24584 27066 24636 27072
rect 24492 26784 24544 26790
rect 24492 26726 24544 26732
rect 24688 26518 24716 27270
rect 24780 26858 24808 28358
rect 24950 28248 25006 28257
rect 24950 28183 24952 28192
rect 25004 28183 25006 28192
rect 24952 28154 25004 28160
rect 24952 28076 25004 28082
rect 24952 28018 25004 28024
rect 24964 27674 24992 28018
rect 24952 27668 25004 27674
rect 24952 27610 25004 27616
rect 24768 26852 24820 26858
rect 24768 26794 24820 26800
rect 25044 26784 25096 26790
rect 25044 26726 25096 26732
rect 24676 26512 24728 26518
rect 24676 26454 24728 26460
rect 24400 26376 24452 26382
rect 24400 26318 24452 26324
rect 24228 24942 24624 24970
rect 24216 24608 24268 24614
rect 24216 24550 24268 24556
rect 24124 23724 24176 23730
rect 24124 23666 24176 23672
rect 23756 21684 23808 21690
rect 23756 21626 23808 21632
rect 24032 21684 24084 21690
rect 24032 21626 24084 21632
rect 23676 21542 23980 21570
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23572 20800 23624 20806
rect 23572 20742 23624 20748
rect 23572 19712 23624 19718
rect 23572 19654 23624 19660
rect 23584 19378 23612 19654
rect 23572 19372 23624 19378
rect 23572 19314 23624 19320
rect 23570 19272 23626 19281
rect 23570 19207 23626 19216
rect 23388 18760 23440 18766
rect 23388 18702 23440 18708
rect 23204 17604 23256 17610
rect 23204 17546 23256 17552
rect 23216 11150 23244 17546
rect 23480 17536 23532 17542
rect 23480 17478 23532 17484
rect 23388 15496 23440 15502
rect 23388 15438 23440 15444
rect 23296 14272 23348 14278
rect 23296 14214 23348 14220
rect 23308 13394 23336 14214
rect 23296 13388 23348 13394
rect 23296 13330 23348 13336
rect 23400 13326 23428 15438
rect 23492 15094 23520 17478
rect 23584 16658 23612 19207
rect 23572 16652 23624 16658
rect 23572 16594 23624 16600
rect 23572 16448 23624 16454
rect 23572 16390 23624 16396
rect 23584 16182 23612 16390
rect 23572 16176 23624 16182
rect 23572 16118 23624 16124
rect 23480 15088 23532 15094
rect 23480 15030 23532 15036
rect 23572 14816 23624 14822
rect 23572 14758 23624 14764
rect 23584 14482 23612 14758
rect 23572 14476 23624 14482
rect 23572 14418 23624 14424
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23480 12776 23532 12782
rect 23480 12718 23532 12724
rect 23492 12322 23520 12718
rect 23584 12714 23612 14418
rect 23676 14346 23704 21286
rect 23756 21004 23808 21010
rect 23756 20946 23808 20952
rect 23768 18222 23796 20946
rect 23848 18352 23900 18358
rect 23848 18294 23900 18300
rect 23756 18216 23808 18222
rect 23756 18158 23808 18164
rect 23768 17814 23796 18158
rect 23756 17808 23808 17814
rect 23756 17750 23808 17756
rect 23860 15706 23888 18294
rect 23848 15700 23900 15706
rect 23848 15642 23900 15648
rect 23664 14340 23716 14346
rect 23664 14282 23716 14288
rect 23952 13258 23980 21542
rect 23940 13252 23992 13258
rect 23940 13194 23992 13200
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 23768 12918 23796 13126
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 23572 12708 23624 12714
rect 23572 12650 23624 12656
rect 23756 12436 23808 12442
rect 23756 12378 23808 12384
rect 23308 12294 23520 12322
rect 23572 12300 23624 12306
rect 23308 11898 23336 12294
rect 23572 12242 23624 12248
rect 23296 11892 23348 11898
rect 23296 11834 23348 11840
rect 23204 11144 23256 11150
rect 23204 11086 23256 11092
rect 22100 11076 22152 11082
rect 22100 11018 22152 11024
rect 23112 11076 23164 11082
rect 23112 11018 23164 11024
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 22112 7818 22140 11018
rect 22560 10464 22612 10470
rect 22560 10406 22612 10412
rect 22572 9994 22600 10406
rect 22560 9988 22612 9994
rect 22560 9930 22612 9936
rect 23308 9042 23336 11834
rect 23480 10668 23532 10674
rect 23480 10610 23532 10616
rect 23492 10198 23520 10610
rect 23584 10266 23612 12242
rect 23768 12238 23796 12378
rect 23756 12232 23808 12238
rect 23756 12174 23808 12180
rect 23768 11014 23796 12174
rect 24228 11558 24256 24550
rect 24400 23520 24452 23526
rect 24400 23462 24452 23468
rect 24308 12164 24360 12170
rect 24308 12106 24360 12112
rect 24216 11552 24268 11558
rect 24216 11494 24268 11500
rect 23756 11008 23808 11014
rect 23756 10950 23808 10956
rect 24320 10606 24348 12106
rect 24308 10600 24360 10606
rect 24308 10542 24360 10548
rect 23848 10532 23900 10538
rect 23848 10474 23900 10480
rect 23572 10260 23624 10266
rect 23572 10202 23624 10208
rect 23480 10192 23532 10198
rect 23480 10134 23532 10140
rect 23860 10062 23888 10474
rect 24308 10124 24360 10130
rect 24308 10066 24360 10072
rect 23848 10056 23900 10062
rect 23848 9998 23900 10004
rect 24320 9654 24348 10066
rect 24308 9648 24360 9654
rect 24308 9590 24360 9596
rect 23296 9036 23348 9042
rect 23296 8978 23348 8984
rect 23480 9036 23532 9042
rect 23480 8978 23532 8984
rect 22376 8968 22428 8974
rect 22376 8910 22428 8916
rect 22100 7812 22152 7818
rect 22100 7754 22152 7760
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 21732 4004 21784 4010
rect 21732 3946 21784 3952
rect 21916 3936 21968 3942
rect 21916 3878 21968 3884
rect 21928 3534 21956 3878
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 22020 2650 22048 7346
rect 22388 6798 22416 8910
rect 23492 8430 23520 8978
rect 23480 8424 23532 8430
rect 23480 8366 23532 8372
rect 23388 8356 23440 8362
rect 23388 8298 23440 8304
rect 22376 6792 22428 6798
rect 22376 6734 22428 6740
rect 22652 3392 22704 3398
rect 22652 3334 22704 3340
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 22008 2644 22060 2650
rect 22008 2586 22060 2592
rect 18604 2508 18656 2514
rect 18604 2450 18656 2456
rect 22664 2446 22692 3334
rect 23400 2514 23428 8298
rect 23492 8242 23520 8366
rect 23492 8214 23612 8242
rect 23480 7472 23532 7478
rect 23480 7414 23532 7420
rect 23492 7002 23520 7414
rect 23584 7274 23612 8214
rect 23572 7268 23624 7274
rect 23572 7210 23624 7216
rect 23480 6996 23532 7002
rect 23480 6938 23532 6944
rect 23388 2508 23440 2514
rect 23388 2450 23440 2456
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 22652 2440 22704 2446
rect 22652 2382 22704 2388
rect 23848 2440 23900 2446
rect 23848 2382 23900 2388
rect 17040 2100 17092 2106
rect 17040 2042 17092 2048
rect 17420 800 17448 2382
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 18064 800 18092 2246
rect 19352 800 19380 2382
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 20640 800 20668 2382
rect 21928 800 21956 2382
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 22572 800 22600 2246
rect 23860 800 23888 2382
rect 24412 2106 24440 23462
rect 24596 22778 24624 24942
rect 24584 22772 24636 22778
rect 24584 22714 24636 22720
rect 24596 21554 24624 22714
rect 24676 21956 24728 21962
rect 24676 21898 24728 21904
rect 24584 21548 24636 21554
rect 24584 21490 24636 21496
rect 24688 21010 24716 21898
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 24582 17776 24638 17785
rect 24582 17711 24638 17720
rect 24596 17678 24624 17711
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 24768 16992 24820 16998
rect 24768 16934 24820 16940
rect 24492 16652 24544 16658
rect 24492 16594 24544 16600
rect 24504 2922 24532 16594
rect 24676 16448 24728 16454
rect 24676 16390 24728 16396
rect 24688 15978 24716 16390
rect 24676 15972 24728 15978
rect 24676 15914 24728 15920
rect 24688 15570 24716 15914
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 24780 12170 24808 16934
rect 24872 15162 24900 20742
rect 24860 15156 24912 15162
rect 24860 15098 24912 15104
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 24964 12434 24992 15098
rect 24872 12406 24992 12434
rect 24872 12374 24900 12406
rect 24860 12368 24912 12374
rect 24860 12310 24912 12316
rect 24768 12164 24820 12170
rect 24768 12106 24820 12112
rect 24768 11076 24820 11082
rect 24768 11018 24820 11024
rect 24780 10810 24808 11018
rect 24768 10804 24820 10810
rect 24768 10746 24820 10752
rect 24768 10668 24820 10674
rect 24768 10610 24820 10616
rect 24780 10266 24808 10610
rect 24768 10260 24820 10266
rect 24768 10202 24820 10208
rect 24584 7336 24636 7342
rect 24584 7278 24636 7284
rect 24596 6458 24624 7278
rect 24584 6452 24636 6458
rect 24584 6394 24636 6400
rect 24492 2916 24544 2922
rect 24492 2858 24544 2864
rect 25056 2310 25084 26726
rect 25148 22234 25176 28494
rect 25332 27826 25360 29650
rect 25412 28756 25464 28762
rect 25412 28698 25464 28704
rect 25240 27798 25360 27826
rect 25136 22228 25188 22234
rect 25136 22170 25188 22176
rect 25240 17270 25268 27798
rect 25424 26382 25452 28698
rect 25412 26376 25464 26382
rect 25412 26318 25464 26324
rect 25412 24812 25464 24818
rect 25412 24754 25464 24760
rect 25424 24410 25452 24754
rect 25412 24404 25464 24410
rect 25412 24346 25464 24352
rect 25516 22094 25544 32778
rect 25686 31920 25742 31929
rect 25686 31855 25688 31864
rect 25740 31855 25742 31864
rect 25688 31826 25740 31832
rect 25792 31822 25820 33215
rect 25872 31884 25924 31890
rect 25872 31826 25924 31832
rect 25780 31816 25832 31822
rect 25780 31758 25832 31764
rect 25780 30184 25832 30190
rect 25780 30126 25832 30132
rect 25596 29232 25648 29238
rect 25596 29174 25648 29180
rect 25608 28218 25636 29174
rect 25596 28212 25648 28218
rect 25596 28154 25648 28160
rect 25792 27996 25820 30126
rect 25884 28370 25912 31826
rect 25976 28762 26004 33458
rect 26148 33380 26200 33386
rect 26148 33322 26200 33328
rect 26240 33380 26292 33386
rect 26240 33322 26292 33328
rect 26160 32978 26188 33322
rect 26252 33153 26280 33322
rect 26238 33144 26294 33153
rect 26238 33079 26294 33088
rect 26148 32972 26200 32978
rect 26200 32932 26280 32960
rect 26148 32914 26200 32920
rect 26148 32836 26200 32842
rect 26148 32778 26200 32784
rect 26056 32768 26108 32774
rect 26056 32710 26108 32716
rect 26068 31754 26096 32710
rect 26160 32366 26188 32778
rect 26148 32360 26200 32366
rect 26148 32302 26200 32308
rect 26056 31748 26108 31754
rect 26056 31690 26108 31696
rect 26252 29714 26280 32932
rect 26700 32224 26752 32230
rect 26700 32166 26752 32172
rect 26608 30660 26660 30666
rect 26608 30602 26660 30608
rect 26332 29776 26384 29782
rect 26332 29718 26384 29724
rect 26240 29708 26292 29714
rect 26240 29650 26292 29656
rect 26148 29504 26200 29510
rect 26148 29446 26200 29452
rect 25964 28756 26016 28762
rect 25964 28698 26016 28704
rect 25964 28416 26016 28422
rect 25884 28364 25964 28370
rect 26016 28364 26096 28370
rect 25884 28342 26096 28364
rect 25700 27968 25820 27996
rect 25596 24608 25648 24614
rect 25596 24550 25648 24556
rect 25608 23798 25636 24550
rect 25596 23792 25648 23798
rect 25596 23734 25648 23740
rect 25608 23186 25636 23734
rect 25596 23180 25648 23186
rect 25596 23122 25648 23128
rect 25700 22094 25728 27968
rect 25780 27872 25832 27878
rect 25780 27814 25832 27820
rect 25792 26994 25820 27814
rect 25964 27396 26016 27402
rect 25964 27338 26016 27344
rect 25780 26988 25832 26994
rect 25780 26930 25832 26936
rect 25976 26586 26004 27338
rect 25964 26580 26016 26586
rect 25964 26522 26016 26528
rect 25872 26376 25924 26382
rect 25872 26318 25924 26324
rect 25884 25430 25912 26318
rect 25872 25424 25924 25430
rect 25872 25366 25924 25372
rect 25780 22568 25832 22574
rect 25780 22510 25832 22516
rect 25792 22234 25820 22510
rect 25780 22228 25832 22234
rect 25780 22170 25832 22176
rect 25332 22066 25544 22094
rect 25608 22066 25728 22094
rect 25332 21962 25360 22066
rect 25320 21956 25372 21962
rect 25320 21898 25372 21904
rect 25228 17264 25280 17270
rect 25228 17206 25280 17212
rect 25332 14958 25360 21898
rect 25412 16584 25464 16590
rect 25412 16526 25464 16532
rect 25424 16114 25452 16526
rect 25412 16108 25464 16114
rect 25412 16050 25464 16056
rect 25320 14952 25372 14958
rect 25320 14894 25372 14900
rect 25608 14385 25636 22066
rect 25688 18420 25740 18426
rect 25688 18362 25740 18368
rect 25594 14376 25650 14385
rect 25594 14311 25596 14320
rect 25648 14311 25650 14320
rect 25596 14282 25648 14288
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 25240 13258 25268 13874
rect 25700 13326 25728 18362
rect 25780 16448 25832 16454
rect 25780 16390 25832 16396
rect 25792 16114 25820 16390
rect 25780 16108 25832 16114
rect 25780 16050 25832 16056
rect 25688 13320 25740 13326
rect 25884 13308 25912 25366
rect 25964 22636 26016 22642
rect 25964 22578 26016 22584
rect 25976 22234 26004 22578
rect 25964 22228 26016 22234
rect 25964 22170 26016 22176
rect 26068 15162 26096 28342
rect 26160 28218 26188 29446
rect 26344 28694 26372 29718
rect 26424 29640 26476 29646
rect 26424 29582 26476 29588
rect 26436 28801 26464 29582
rect 26516 29504 26568 29510
rect 26516 29446 26568 29452
rect 26422 28792 26478 28801
rect 26422 28727 26478 28736
rect 26332 28688 26384 28694
rect 26332 28630 26384 28636
rect 26240 28620 26292 28626
rect 26240 28562 26292 28568
rect 26148 28212 26200 28218
rect 26148 28154 26200 28160
rect 26252 27538 26280 28562
rect 26528 28490 26556 29446
rect 26620 29102 26648 30602
rect 26608 29096 26660 29102
rect 26608 29038 26660 29044
rect 26516 28484 26568 28490
rect 26516 28426 26568 28432
rect 26240 27532 26292 27538
rect 26240 27474 26292 27480
rect 26620 27033 26648 29038
rect 26712 27606 26740 32166
rect 26790 29200 26846 29209
rect 26988 29170 27016 35974
rect 27264 35766 27292 36586
rect 27436 36372 27488 36378
rect 27436 36314 27488 36320
rect 27252 35760 27304 35766
rect 27252 35702 27304 35708
rect 27344 35488 27396 35494
rect 27344 35430 27396 35436
rect 27068 35148 27120 35154
rect 27068 35090 27120 35096
rect 27080 32230 27108 35090
rect 27356 34678 27384 35430
rect 27344 34672 27396 34678
rect 27344 34614 27396 34620
rect 27250 34232 27306 34241
rect 27250 34167 27306 34176
rect 27264 34066 27292 34167
rect 27252 34060 27304 34066
rect 27252 34002 27304 34008
rect 27344 33584 27396 33590
rect 27344 33526 27396 33532
rect 27252 33448 27304 33454
rect 27252 33390 27304 33396
rect 27264 32502 27292 33390
rect 27356 33114 27384 33526
rect 27344 33108 27396 33114
rect 27344 33050 27396 33056
rect 27344 32836 27396 32842
rect 27344 32778 27396 32784
rect 27252 32496 27304 32502
rect 27172 32444 27252 32450
rect 27172 32438 27304 32444
rect 27172 32422 27292 32438
rect 27068 32224 27120 32230
rect 27068 32166 27120 32172
rect 27080 31890 27108 32166
rect 27068 31884 27120 31890
rect 27068 31826 27120 31832
rect 27172 30802 27200 32422
rect 27252 31272 27304 31278
rect 27252 31214 27304 31220
rect 27160 30796 27212 30802
rect 27160 30738 27212 30744
rect 27264 30138 27292 31214
rect 27356 30326 27384 32778
rect 27448 32434 27476 36314
rect 27540 36242 27568 36654
rect 27988 36644 28040 36650
rect 27988 36586 28040 36592
rect 27528 36236 27580 36242
rect 27528 36178 27580 36184
rect 27620 36236 27672 36242
rect 27620 36178 27672 36184
rect 27632 36122 27660 36178
rect 27540 36094 27660 36122
rect 28000 36106 28028 36586
rect 27988 36100 28040 36106
rect 27540 36038 27568 36094
rect 27988 36042 28040 36048
rect 27528 36032 27580 36038
rect 27528 35974 27580 35980
rect 28172 35012 28224 35018
rect 28172 34954 28224 34960
rect 28264 35012 28316 35018
rect 28264 34954 28316 34960
rect 28184 34746 28212 34954
rect 28172 34740 28224 34746
rect 28172 34682 28224 34688
rect 27896 34536 27948 34542
rect 27896 34478 27948 34484
rect 27712 33924 27764 33930
rect 27712 33866 27764 33872
rect 27724 33658 27752 33866
rect 27712 33652 27764 33658
rect 27712 33594 27764 33600
rect 27908 33454 27936 34478
rect 28276 34202 28304 34954
rect 28368 34474 28396 36654
rect 28448 35692 28500 35698
rect 28448 35634 28500 35640
rect 28356 34468 28408 34474
rect 28356 34410 28408 34416
rect 28460 34354 28488 35634
rect 28368 34326 28488 34354
rect 28264 34196 28316 34202
rect 28264 34138 28316 34144
rect 28368 33998 28396 34326
rect 28356 33992 28408 33998
rect 28356 33934 28408 33940
rect 27896 33448 27948 33454
rect 27896 33390 27948 33396
rect 27436 32428 27488 32434
rect 27436 32370 27488 32376
rect 27618 31920 27674 31929
rect 27618 31855 27620 31864
rect 27672 31855 27674 31864
rect 27620 31826 27672 31832
rect 27908 31754 27936 33390
rect 27988 32836 28040 32842
rect 27988 32778 28040 32784
rect 27724 31726 27936 31754
rect 27344 30320 27396 30326
rect 27344 30262 27396 30268
rect 27528 30252 27580 30258
rect 27528 30194 27580 30200
rect 27264 30110 27384 30138
rect 27160 29504 27212 29510
rect 27160 29446 27212 29452
rect 26790 29135 26846 29144
rect 26976 29164 27028 29170
rect 26804 28994 26832 29135
rect 26976 29106 27028 29112
rect 26804 28966 26924 28994
rect 26700 27600 26752 27606
rect 26700 27542 26752 27548
rect 26896 27402 26924 28966
rect 27172 28626 27200 29446
rect 27252 29096 27304 29102
rect 27252 29038 27304 29044
rect 27160 28620 27212 28626
rect 27160 28562 27212 28568
rect 26884 27396 26936 27402
rect 26884 27338 26936 27344
rect 26606 27024 26662 27033
rect 26606 26959 26662 26968
rect 26424 26308 26476 26314
rect 26424 26250 26476 26256
rect 26436 26042 26464 26250
rect 26424 26036 26476 26042
rect 26424 25978 26476 25984
rect 26896 23662 26924 27338
rect 27160 25288 27212 25294
rect 27160 25230 27212 25236
rect 27172 24818 27200 25230
rect 27160 24812 27212 24818
rect 27160 24754 27212 24760
rect 27264 24750 27292 29038
rect 27356 28490 27384 30110
rect 27540 29510 27568 30194
rect 27528 29504 27580 29510
rect 27528 29446 27580 29452
rect 27540 28762 27568 29446
rect 27620 29028 27672 29034
rect 27620 28970 27672 28976
rect 27528 28756 27580 28762
rect 27528 28698 27580 28704
rect 27632 28490 27660 28970
rect 27344 28484 27396 28490
rect 27344 28426 27396 28432
rect 27620 28484 27672 28490
rect 27620 28426 27672 28432
rect 27252 24744 27304 24750
rect 27252 24686 27304 24692
rect 26884 23656 26936 23662
rect 26884 23598 26936 23604
rect 26148 23112 26200 23118
rect 26148 23054 26200 23060
rect 26160 22778 26188 23054
rect 26148 22772 26200 22778
rect 26148 22714 26200 22720
rect 26332 22024 26384 22030
rect 26332 21966 26384 21972
rect 26240 21480 26292 21486
rect 26240 21422 26292 21428
rect 26252 20602 26280 21422
rect 26240 20596 26292 20602
rect 26240 20538 26292 20544
rect 26344 20466 26372 21966
rect 26792 20868 26844 20874
rect 26792 20810 26844 20816
rect 26804 20602 26832 20810
rect 26792 20596 26844 20602
rect 26792 20538 26844 20544
rect 26332 20460 26384 20466
rect 26332 20402 26384 20408
rect 26896 20058 26924 23598
rect 27356 21078 27384 28426
rect 27724 28014 27752 31726
rect 28000 30122 28028 32778
rect 28368 32473 28396 33934
rect 28448 33856 28500 33862
rect 28448 33798 28500 33804
rect 28460 32774 28488 33798
rect 28552 33590 28580 37062
rect 28724 36916 28776 36922
rect 28724 36858 28776 36864
rect 28632 36780 28684 36786
rect 28632 36722 28684 36728
rect 28644 35834 28672 36722
rect 28632 35828 28684 35834
rect 28632 35770 28684 35776
rect 28736 34406 28764 36858
rect 28816 36848 28868 36854
rect 28816 36790 28868 36796
rect 28828 35834 28856 36790
rect 28816 35828 28868 35834
rect 28816 35770 28868 35776
rect 28920 35766 28948 37062
rect 29736 36644 29788 36650
rect 29736 36586 29788 36592
rect 28908 35760 28960 35766
rect 28908 35702 28960 35708
rect 29748 35154 29776 36586
rect 29736 35148 29788 35154
rect 29736 35090 29788 35096
rect 28724 34400 28776 34406
rect 28724 34342 28776 34348
rect 28540 33584 28592 33590
rect 28540 33526 28592 33532
rect 28448 32768 28500 32774
rect 28448 32710 28500 32716
rect 28354 32464 28410 32473
rect 28736 32434 28764 34342
rect 29644 33924 29696 33930
rect 29644 33866 29696 33872
rect 29656 33522 29684 33866
rect 29840 33590 29868 37062
rect 31036 36922 31064 37062
rect 31024 36916 31076 36922
rect 31024 36858 31076 36864
rect 33060 36310 33088 37062
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 33048 36304 33100 36310
rect 33048 36246 33100 36252
rect 36096 36174 36124 39200
rect 37186 38856 37242 38865
rect 37186 38791 37242 38800
rect 36176 37256 36228 37262
rect 36176 37198 36228 37204
rect 36084 36168 36136 36174
rect 36084 36110 36136 36116
rect 34520 36032 34572 36038
rect 34520 35974 34572 35980
rect 29828 33584 29880 33590
rect 29828 33526 29880 33532
rect 29644 33516 29696 33522
rect 29644 33458 29696 33464
rect 29092 33312 29144 33318
rect 29092 33254 29144 33260
rect 29184 33312 29236 33318
rect 29184 33254 29236 33260
rect 29104 32978 29132 33254
rect 29092 32972 29144 32978
rect 29092 32914 29144 32920
rect 28354 32399 28410 32408
rect 28724 32428 28776 32434
rect 28080 32224 28132 32230
rect 28080 32166 28132 32172
rect 28092 31482 28120 32166
rect 28264 31816 28316 31822
rect 28264 31758 28316 31764
rect 28172 31680 28224 31686
rect 28172 31622 28224 31628
rect 28080 31476 28132 31482
rect 28080 31418 28132 31424
rect 28092 30870 28120 31418
rect 28184 31346 28212 31622
rect 28172 31340 28224 31346
rect 28172 31282 28224 31288
rect 28080 30864 28132 30870
rect 28080 30806 28132 30812
rect 27988 30116 28040 30122
rect 27988 30058 28040 30064
rect 28172 30048 28224 30054
rect 28172 29990 28224 29996
rect 28184 29714 28212 29990
rect 28172 29708 28224 29714
rect 28172 29650 28224 29656
rect 27988 29096 28040 29102
rect 27988 29038 28040 29044
rect 27804 28620 27856 28626
rect 27804 28562 27856 28568
rect 27712 28008 27764 28014
rect 27712 27950 27764 27956
rect 27724 26858 27752 27950
rect 27816 27946 27844 28562
rect 27804 27940 27856 27946
rect 27804 27882 27856 27888
rect 27712 26852 27764 26858
rect 27712 26794 27764 26800
rect 27528 24880 27580 24886
rect 27528 24822 27580 24828
rect 27540 23730 27568 24822
rect 27724 24138 27752 26794
rect 27816 26518 27844 27882
rect 28000 27606 28028 29038
rect 27988 27600 28040 27606
rect 27988 27542 28040 27548
rect 28080 27328 28132 27334
rect 28080 27270 28132 27276
rect 27896 26784 27948 26790
rect 27896 26726 27948 26732
rect 27804 26512 27856 26518
rect 27804 26454 27856 26460
rect 27712 24132 27764 24138
rect 27712 24074 27764 24080
rect 27908 23798 27936 26726
rect 27896 23792 27948 23798
rect 27896 23734 27948 23740
rect 27528 23724 27580 23730
rect 27528 23666 27580 23672
rect 27988 23656 28040 23662
rect 27988 23598 28040 23604
rect 27804 22704 27856 22710
rect 27804 22646 27856 22652
rect 27436 21344 27488 21350
rect 27436 21286 27488 21292
rect 27344 21072 27396 21078
rect 27344 21014 27396 21020
rect 27448 21010 27476 21286
rect 27436 21004 27488 21010
rect 27436 20946 27488 20952
rect 27252 20460 27304 20466
rect 27252 20402 27304 20408
rect 26884 20052 26936 20058
rect 26884 19994 26936 20000
rect 26148 17128 26200 17134
rect 26148 17070 26200 17076
rect 26160 16250 26188 17070
rect 26240 17060 26292 17066
rect 26240 17002 26292 17008
rect 26252 16590 26280 17002
rect 26332 16992 26384 16998
rect 26332 16934 26384 16940
rect 26240 16584 26292 16590
rect 26240 16526 26292 16532
rect 26344 16522 26372 16934
rect 26332 16516 26384 16522
rect 26332 16458 26384 16464
rect 26148 16244 26200 16250
rect 26148 16186 26200 16192
rect 26344 16046 26372 16458
rect 26332 16040 26384 16046
rect 26332 15982 26384 15988
rect 26896 15570 26924 19994
rect 27264 18766 27292 20402
rect 27448 19922 27476 20946
rect 27528 20256 27580 20262
rect 27528 20198 27580 20204
rect 27436 19916 27488 19922
rect 27436 19858 27488 19864
rect 27540 19786 27568 20198
rect 27712 19984 27764 19990
rect 27712 19926 27764 19932
rect 27528 19780 27580 19786
rect 27528 19722 27580 19728
rect 27252 18760 27304 18766
rect 27252 18702 27304 18708
rect 27528 17808 27580 17814
rect 27528 17750 27580 17756
rect 27160 17672 27212 17678
rect 27160 17614 27212 17620
rect 26976 16992 27028 16998
rect 26976 16934 27028 16940
rect 26884 15564 26936 15570
rect 26884 15506 26936 15512
rect 26516 15428 26568 15434
rect 26516 15370 26568 15376
rect 26528 15162 26556 15370
rect 26056 15156 26108 15162
rect 26056 15098 26108 15104
rect 26516 15156 26568 15162
rect 26516 15098 26568 15104
rect 26068 14770 26096 15098
rect 26068 14742 26188 14770
rect 26056 14612 26108 14618
rect 26056 14554 26108 14560
rect 26068 14006 26096 14554
rect 26160 14550 26188 14742
rect 26148 14544 26200 14550
rect 26148 14486 26200 14492
rect 25964 14000 26016 14006
rect 25964 13942 26016 13948
rect 26056 14000 26108 14006
rect 26056 13942 26108 13948
rect 25976 13530 26004 13942
rect 26528 13870 26556 15098
rect 26516 13864 26568 13870
rect 26516 13806 26568 13812
rect 25964 13524 26016 13530
rect 25964 13466 26016 13472
rect 25964 13320 26016 13326
rect 25884 13280 25964 13308
rect 25688 13262 25740 13268
rect 25964 13262 26016 13268
rect 25228 13252 25280 13258
rect 25228 13194 25280 13200
rect 25320 13184 25372 13190
rect 25320 13126 25372 13132
rect 25332 12986 25360 13126
rect 25320 12980 25372 12986
rect 25320 12922 25372 12928
rect 25700 12434 25728 13262
rect 26056 13184 26108 13190
rect 26056 13126 26108 13132
rect 25700 12406 25912 12434
rect 25780 11688 25832 11694
rect 25780 11630 25832 11636
rect 25792 11218 25820 11630
rect 25780 11212 25832 11218
rect 25780 11154 25832 11160
rect 25504 11144 25556 11150
rect 25504 11086 25556 11092
rect 25320 11076 25372 11082
rect 25320 11018 25372 11024
rect 25228 10736 25280 10742
rect 25228 10678 25280 10684
rect 25240 10266 25268 10678
rect 25228 10260 25280 10266
rect 25228 10202 25280 10208
rect 25228 9580 25280 9586
rect 25228 9522 25280 9528
rect 25240 8974 25268 9522
rect 25332 9518 25360 11018
rect 25412 11008 25464 11014
rect 25412 10950 25464 10956
rect 25424 10674 25452 10950
rect 25412 10668 25464 10674
rect 25412 10610 25464 10616
rect 25516 10538 25544 11086
rect 25884 10810 25912 12406
rect 25872 10804 25924 10810
rect 25872 10746 25924 10752
rect 25504 10532 25556 10538
rect 25504 10474 25556 10480
rect 25412 10464 25464 10470
rect 25412 10406 25464 10412
rect 25424 10062 25452 10406
rect 25412 10056 25464 10062
rect 25412 9998 25464 10004
rect 25688 9920 25740 9926
rect 25688 9862 25740 9868
rect 25700 9586 25728 9862
rect 25688 9580 25740 9586
rect 25688 9522 25740 9528
rect 25320 9512 25372 9518
rect 25320 9454 25372 9460
rect 25228 8968 25280 8974
rect 25228 8910 25280 8916
rect 25240 8566 25268 8910
rect 25228 8560 25280 8566
rect 25228 8502 25280 8508
rect 25332 6322 25360 9454
rect 25964 9444 26016 9450
rect 25964 9386 26016 9392
rect 25976 9178 26004 9386
rect 25964 9172 26016 9178
rect 25964 9114 26016 9120
rect 25596 7880 25648 7886
rect 25596 7822 25648 7828
rect 25320 6316 25372 6322
rect 25320 6258 25372 6264
rect 25228 5568 25280 5574
rect 25228 5510 25280 5516
rect 25240 2446 25268 5510
rect 25608 2582 25636 7822
rect 26068 7818 26096 13126
rect 26988 12170 27016 16934
rect 27172 12434 27200 17614
rect 27252 17536 27304 17542
rect 27252 17478 27304 17484
rect 27264 16182 27292 17478
rect 27344 17196 27396 17202
rect 27344 17138 27396 17144
rect 27356 16454 27384 17138
rect 27344 16448 27396 16454
rect 27344 16390 27396 16396
rect 27436 16448 27488 16454
rect 27436 16390 27488 16396
rect 27252 16176 27304 16182
rect 27252 16118 27304 16124
rect 27448 15434 27476 16390
rect 27436 15428 27488 15434
rect 27436 15370 27488 15376
rect 27436 15020 27488 15026
rect 27436 14962 27488 14968
rect 27172 12406 27292 12434
rect 26516 12164 26568 12170
rect 26516 12106 26568 12112
rect 26976 12164 27028 12170
rect 26976 12106 27028 12112
rect 26528 11354 26556 12106
rect 26516 11348 26568 11354
rect 26516 11290 26568 11296
rect 27264 11234 27292 12406
rect 27344 11552 27396 11558
rect 27344 11494 27396 11500
rect 27356 11354 27384 11494
rect 27344 11348 27396 11354
rect 27344 11290 27396 11296
rect 27264 11206 27384 11234
rect 27252 11144 27304 11150
rect 27252 11086 27304 11092
rect 26332 10600 26384 10606
rect 26332 10542 26384 10548
rect 26344 9586 26372 10542
rect 26332 9580 26384 9586
rect 26332 9522 26384 9528
rect 26344 9382 26372 9522
rect 26516 9512 26568 9518
rect 26516 9454 26568 9460
rect 26240 9376 26292 9382
rect 26240 9318 26292 9324
rect 26332 9376 26384 9382
rect 26332 9318 26384 9324
rect 26252 8974 26280 9318
rect 26528 9178 26556 9454
rect 26516 9172 26568 9178
rect 26516 9114 26568 9120
rect 26240 8968 26292 8974
rect 26240 8910 26292 8916
rect 26240 8492 26292 8498
rect 26240 8434 26292 8440
rect 26056 7812 26108 7818
rect 26056 7754 26108 7760
rect 25688 6112 25740 6118
rect 25688 6054 25740 6060
rect 25700 5710 25728 6054
rect 25688 5704 25740 5710
rect 25688 5646 25740 5652
rect 26252 2650 26280 8434
rect 27264 2922 27292 11086
rect 27356 10674 27384 11206
rect 27344 10668 27396 10674
rect 27344 10610 27396 10616
rect 27356 8906 27384 10610
rect 27344 8900 27396 8906
rect 27344 8842 27396 8848
rect 27344 7880 27396 7886
rect 27344 7822 27396 7828
rect 27252 2916 27304 2922
rect 27252 2858 27304 2864
rect 27356 2650 27384 7822
rect 27448 6118 27476 14962
rect 27540 14958 27568 17750
rect 27620 17264 27672 17270
rect 27620 17206 27672 17212
rect 27632 16250 27660 17206
rect 27620 16244 27672 16250
rect 27620 16186 27672 16192
rect 27724 15162 27752 19926
rect 27816 19922 27844 22646
rect 27896 20460 27948 20466
rect 27896 20402 27948 20408
rect 27804 19916 27856 19922
rect 27804 19858 27856 19864
rect 27816 17814 27844 19858
rect 27908 19446 27936 20402
rect 27896 19440 27948 19446
rect 27896 19382 27948 19388
rect 27804 17808 27856 17814
rect 27804 17750 27856 17756
rect 27908 16590 27936 19382
rect 28000 16794 28028 23598
rect 28092 22710 28120 27270
rect 28276 25906 28304 31758
rect 28368 26994 28396 32399
rect 28724 32370 28776 32376
rect 29000 32360 29052 32366
rect 29000 32302 29052 32308
rect 29012 32026 29040 32302
rect 29000 32020 29052 32026
rect 29000 31962 29052 31968
rect 28540 30592 28592 30598
rect 28540 30534 28592 30540
rect 28552 29850 28580 30534
rect 28540 29844 28592 29850
rect 28540 29786 28592 29792
rect 28552 29714 28580 29786
rect 28540 29708 28592 29714
rect 28540 29650 28592 29656
rect 28448 29640 28500 29646
rect 28448 29582 28500 29588
rect 28460 29034 28488 29582
rect 29196 29578 29224 33254
rect 29276 30728 29328 30734
rect 29276 30670 29328 30676
rect 29288 30394 29316 30670
rect 29276 30388 29328 30394
rect 29276 30330 29328 30336
rect 29184 29572 29236 29578
rect 29184 29514 29236 29520
rect 28448 29028 28500 29034
rect 28448 28970 28500 28976
rect 28356 26988 28408 26994
rect 28356 26930 28408 26936
rect 28264 25900 28316 25906
rect 28264 25842 28316 25848
rect 28172 23112 28224 23118
rect 28172 23054 28224 23060
rect 28080 22704 28132 22710
rect 28080 22646 28132 22652
rect 28080 22568 28132 22574
rect 28080 22510 28132 22516
rect 28092 21554 28120 22510
rect 28080 21548 28132 21554
rect 28080 21490 28132 21496
rect 28092 21146 28120 21490
rect 28080 21140 28132 21146
rect 28080 21082 28132 21088
rect 28080 17536 28132 17542
rect 28080 17478 28132 17484
rect 28092 17202 28120 17478
rect 28080 17196 28132 17202
rect 28080 17138 28132 17144
rect 27988 16788 28040 16794
rect 27988 16730 28040 16736
rect 27896 16584 27948 16590
rect 27896 16526 27948 16532
rect 27896 16040 27948 16046
rect 27896 15982 27948 15988
rect 27712 15156 27764 15162
rect 27712 15098 27764 15104
rect 27908 15094 27936 15982
rect 28184 15978 28212 23054
rect 28276 17678 28304 25842
rect 28356 24744 28408 24750
rect 28356 24686 28408 24692
rect 28368 18329 28396 24686
rect 28460 23322 28488 28970
rect 29460 26580 29512 26586
rect 29460 26522 29512 26528
rect 29092 25764 29144 25770
rect 29092 25706 29144 25712
rect 29184 25764 29236 25770
rect 29184 25706 29236 25712
rect 28540 25696 28592 25702
rect 28540 25638 28592 25644
rect 28552 25294 28580 25638
rect 28540 25288 28592 25294
rect 28540 25230 28592 25236
rect 28632 25152 28684 25158
rect 28632 25094 28684 25100
rect 28540 24744 28592 24750
rect 28540 24686 28592 24692
rect 28552 24274 28580 24686
rect 28540 24268 28592 24274
rect 28540 24210 28592 24216
rect 28644 24138 28672 25094
rect 29104 24818 29132 25706
rect 29196 25294 29224 25706
rect 29184 25288 29236 25294
rect 29184 25230 29236 25236
rect 29196 24954 29224 25230
rect 29184 24948 29236 24954
rect 29184 24890 29236 24896
rect 29092 24812 29144 24818
rect 29092 24754 29144 24760
rect 28632 24132 28684 24138
rect 28632 24074 28684 24080
rect 28908 24064 28960 24070
rect 28908 24006 28960 24012
rect 28448 23316 28500 23322
rect 28448 23258 28500 23264
rect 28724 23112 28776 23118
rect 28724 23054 28776 23060
rect 28448 22976 28500 22982
rect 28448 22918 28500 22924
rect 28460 21418 28488 22918
rect 28736 22778 28764 23054
rect 28724 22772 28776 22778
rect 28724 22714 28776 22720
rect 28920 22642 28948 24006
rect 29092 23860 29144 23866
rect 29092 23802 29144 23808
rect 28908 22636 28960 22642
rect 28908 22578 28960 22584
rect 28448 21412 28500 21418
rect 28448 21354 28500 21360
rect 28460 20874 28488 21354
rect 29104 21146 29132 23802
rect 29092 21140 29144 21146
rect 29092 21082 29144 21088
rect 28632 20936 28684 20942
rect 28632 20878 28684 20884
rect 28448 20868 28500 20874
rect 28448 20810 28500 20816
rect 28644 20466 28672 20878
rect 28632 20460 28684 20466
rect 28632 20402 28684 20408
rect 28354 18320 28410 18329
rect 28354 18255 28410 18264
rect 28264 17672 28316 17678
rect 28264 17614 28316 17620
rect 28368 17338 28396 18255
rect 28356 17332 28408 17338
rect 28356 17274 28408 17280
rect 28540 16992 28592 16998
rect 28540 16934 28592 16940
rect 28172 15972 28224 15978
rect 28172 15914 28224 15920
rect 27896 15088 27948 15094
rect 27896 15030 27948 15036
rect 27528 14952 27580 14958
rect 27528 14894 27580 14900
rect 27528 13864 27580 13870
rect 27528 13806 27580 13812
rect 27540 8634 27568 13806
rect 27908 13326 27936 15030
rect 28448 14272 28500 14278
rect 28448 14214 28500 14220
rect 28460 13938 28488 14214
rect 28448 13932 28500 13938
rect 28448 13874 28500 13880
rect 27896 13320 27948 13326
rect 27896 13262 27948 13268
rect 28172 11688 28224 11694
rect 28172 11630 28224 11636
rect 28356 11688 28408 11694
rect 28356 11630 28408 11636
rect 28184 11218 28212 11630
rect 28172 11212 28224 11218
rect 28172 11154 28224 11160
rect 28368 10810 28396 11630
rect 28552 11626 28580 16934
rect 28540 11620 28592 11626
rect 28540 11562 28592 11568
rect 28552 11082 28580 11562
rect 28540 11076 28592 11082
rect 28540 11018 28592 11024
rect 28356 10804 28408 10810
rect 28356 10746 28408 10752
rect 28644 10130 28672 20402
rect 29472 18426 29500 26522
rect 29656 24410 29684 33458
rect 34152 32904 34204 32910
rect 34152 32846 34204 32852
rect 29920 32292 29972 32298
rect 29920 32234 29972 32240
rect 29828 31340 29880 31346
rect 29828 31282 29880 31288
rect 29736 30252 29788 30258
rect 29736 30194 29788 30200
rect 29748 29850 29776 30194
rect 29736 29844 29788 29850
rect 29736 29786 29788 29792
rect 29736 27464 29788 27470
rect 29840 27452 29868 31282
rect 29788 27424 29868 27452
rect 29736 27406 29788 27412
rect 29644 24404 29696 24410
rect 29644 24346 29696 24352
rect 29748 24342 29776 27406
rect 29932 25838 29960 32234
rect 30012 31816 30064 31822
rect 30012 31758 30064 31764
rect 30024 31346 30052 31758
rect 30012 31340 30064 31346
rect 30012 31282 30064 31288
rect 32956 29232 33008 29238
rect 32956 29174 33008 29180
rect 32968 28490 32996 29174
rect 32956 28484 33008 28490
rect 32956 28426 33008 28432
rect 31944 26988 31996 26994
rect 31944 26930 31996 26936
rect 31956 26586 31984 26930
rect 31944 26580 31996 26586
rect 31944 26522 31996 26528
rect 31852 26376 31904 26382
rect 31852 26318 31904 26324
rect 29920 25832 29972 25838
rect 29920 25774 29972 25780
rect 30104 25832 30156 25838
rect 30104 25774 30156 25780
rect 30472 25832 30524 25838
rect 30472 25774 30524 25780
rect 29736 24336 29788 24342
rect 29736 24278 29788 24284
rect 29932 24274 29960 25774
rect 30116 25498 30144 25774
rect 30104 25492 30156 25498
rect 30104 25434 30156 25440
rect 29920 24268 29972 24274
rect 29920 24210 29972 24216
rect 29828 23656 29880 23662
rect 29828 23598 29880 23604
rect 29840 23186 29868 23598
rect 29920 23588 29972 23594
rect 29920 23530 29972 23536
rect 29828 23180 29880 23186
rect 29828 23122 29880 23128
rect 29932 23050 29960 23530
rect 29920 23044 29972 23050
rect 29920 22986 29972 22992
rect 30380 18624 30432 18630
rect 30380 18566 30432 18572
rect 29460 18420 29512 18426
rect 29460 18362 29512 18368
rect 29368 17672 29420 17678
rect 29368 17614 29420 17620
rect 29000 16652 29052 16658
rect 29000 16594 29052 16600
rect 29012 16114 29040 16594
rect 29000 16108 29052 16114
rect 29000 16050 29052 16056
rect 29380 15026 29408 17614
rect 29472 17134 29500 18362
rect 30196 18216 30248 18222
rect 30196 18158 30248 18164
rect 30208 17678 30236 18158
rect 30196 17672 30248 17678
rect 30196 17614 30248 17620
rect 29920 17536 29972 17542
rect 29920 17478 29972 17484
rect 29460 17128 29512 17134
rect 29460 17070 29512 17076
rect 29736 17060 29788 17066
rect 29736 17002 29788 17008
rect 29748 16590 29776 17002
rect 29932 16658 29960 17478
rect 29920 16652 29972 16658
rect 29920 16594 29972 16600
rect 29736 16584 29788 16590
rect 29736 16526 29788 16532
rect 29748 16250 29776 16526
rect 29736 16244 29788 16250
rect 29736 16186 29788 16192
rect 29368 15020 29420 15026
rect 29368 14962 29420 14968
rect 29000 14816 29052 14822
rect 29000 14758 29052 14764
rect 29012 14414 29040 14758
rect 29184 14476 29236 14482
rect 29184 14418 29236 14424
rect 29000 14408 29052 14414
rect 29000 14350 29052 14356
rect 29196 12986 29224 14418
rect 30392 14346 30420 18566
rect 30484 16590 30512 25774
rect 31864 25770 31892 26318
rect 32588 26308 32640 26314
rect 32588 26250 32640 26256
rect 32600 26042 32628 26250
rect 32588 26036 32640 26042
rect 32588 25978 32640 25984
rect 31852 25764 31904 25770
rect 31852 25706 31904 25712
rect 32968 23050 32996 28426
rect 34164 27130 34192 32846
rect 34532 32570 34560 35974
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34520 32564 34572 32570
rect 34520 32506 34572 32512
rect 35440 32428 35492 32434
rect 35440 32370 35492 32376
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35452 29850 35480 32370
rect 35440 29844 35492 29850
rect 35440 29786 35492 29792
rect 34612 29708 34664 29714
rect 34612 29650 34664 29656
rect 34152 27124 34204 27130
rect 34152 27066 34204 27072
rect 34624 27062 34652 29650
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35900 27872 35952 27878
rect 35900 27814 35952 27820
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34612 27056 34664 27062
rect 34612 26998 34664 27004
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 33232 26512 33284 26518
rect 33232 26454 33284 26460
rect 33244 26314 33272 26454
rect 33232 26308 33284 26314
rect 33232 26250 33284 26256
rect 33244 23730 33272 26250
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34704 24200 34756 24206
rect 34704 24142 34756 24148
rect 33232 23724 33284 23730
rect 33232 23666 33284 23672
rect 34428 23520 34480 23526
rect 34428 23462 34480 23468
rect 32956 23044 33008 23050
rect 32956 22986 33008 22992
rect 30930 22672 30986 22681
rect 34440 22642 34468 23462
rect 34716 22778 34744 24142
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34704 22772 34756 22778
rect 34704 22714 34756 22720
rect 30930 22607 30986 22616
rect 31300 22636 31352 22642
rect 30944 20942 30972 22607
rect 31300 22578 31352 22584
rect 34428 22636 34480 22642
rect 34428 22578 34480 22584
rect 31312 22098 31340 22578
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 31300 22092 31352 22098
rect 31300 22034 31352 22040
rect 35912 21622 35940 27814
rect 36188 25226 36216 37198
rect 36820 37188 36872 37194
rect 36820 37130 36872 37136
rect 36544 36100 36596 36106
rect 36544 36042 36596 36048
rect 36556 35290 36584 36042
rect 36544 35284 36596 35290
rect 36544 35226 36596 35232
rect 36636 34604 36688 34610
rect 36636 34546 36688 34552
rect 36648 34202 36676 34546
rect 36636 34196 36688 34202
rect 36636 34138 36688 34144
rect 36832 33998 36860 37130
rect 37200 36378 37228 38791
rect 37188 36372 37240 36378
rect 37188 36314 37240 36320
rect 37280 36168 37332 36174
rect 37280 36110 37332 36116
rect 36820 33992 36872 33998
rect 36820 33934 36872 33940
rect 36832 30326 36860 33934
rect 36820 30320 36872 30326
rect 36820 30262 36872 30268
rect 36176 25220 36228 25226
rect 36176 25162 36228 25168
rect 35992 23044 36044 23050
rect 35992 22986 36044 22992
rect 35900 21616 35952 21622
rect 35900 21558 35952 21564
rect 31668 21548 31720 21554
rect 31668 21490 31720 21496
rect 30932 20936 30984 20942
rect 30932 20878 30984 20884
rect 30944 20466 30972 20878
rect 31576 20800 31628 20806
rect 31576 20742 31628 20748
rect 31588 20466 31616 20742
rect 30932 20460 30984 20466
rect 30932 20402 30984 20408
rect 31576 20460 31628 20466
rect 31576 20402 31628 20408
rect 31116 20392 31168 20398
rect 31116 20334 31168 20340
rect 31128 19922 31156 20334
rect 31116 19916 31168 19922
rect 31116 19858 31168 19864
rect 31680 19514 31708 21490
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 31760 20936 31812 20942
rect 31760 20878 31812 20884
rect 31772 20602 31800 20878
rect 31852 20868 31904 20874
rect 31852 20810 31904 20816
rect 31760 20596 31812 20602
rect 31760 20538 31812 20544
rect 31864 20466 31892 20810
rect 31852 20460 31904 20466
rect 31852 20402 31904 20408
rect 31668 19508 31720 19514
rect 31668 19450 31720 19456
rect 31864 19378 31892 20402
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 30840 19372 30892 19378
rect 30840 19314 30892 19320
rect 31852 19372 31904 19378
rect 31852 19314 31904 19320
rect 33324 19372 33376 19378
rect 33324 19314 33376 19320
rect 30564 17604 30616 17610
rect 30564 17546 30616 17552
rect 30472 16584 30524 16590
rect 30472 16526 30524 16532
rect 30288 14340 30340 14346
rect 30288 14282 30340 14288
rect 30380 14340 30432 14346
rect 30380 14282 30432 14288
rect 30300 14074 30328 14282
rect 30288 14068 30340 14074
rect 30288 14010 30340 14016
rect 30484 14006 30512 16526
rect 30472 14000 30524 14006
rect 30472 13942 30524 13948
rect 29184 12980 29236 12986
rect 29184 12922 29236 12928
rect 29920 10600 29972 10606
rect 29920 10542 29972 10548
rect 28632 10124 28684 10130
rect 28632 10066 28684 10072
rect 27712 9580 27764 9586
rect 27712 9522 27764 9528
rect 27528 8628 27580 8634
rect 27528 8570 27580 8576
rect 27528 6316 27580 6322
rect 27528 6258 27580 6264
rect 27436 6112 27488 6118
rect 27436 6054 27488 6060
rect 26240 2644 26292 2650
rect 26240 2586 26292 2592
rect 27344 2644 27396 2650
rect 27344 2586 27396 2592
rect 27540 2582 27568 6258
rect 27724 5914 27752 9522
rect 27712 5908 27764 5914
rect 27712 5850 27764 5856
rect 29932 5234 29960 10542
rect 30288 5704 30340 5710
rect 30288 5646 30340 5652
rect 29920 5228 29972 5234
rect 29920 5170 29972 5176
rect 30300 2650 30328 5646
rect 30576 3466 30604 17546
rect 30852 12306 30880 19314
rect 33336 18290 33364 19314
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 33324 18284 33376 18290
rect 33324 18226 33376 18232
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34520 15020 34572 15026
rect 34520 14962 34572 14968
rect 31944 14408 31996 14414
rect 31944 14350 31996 14356
rect 31956 13462 31984 14350
rect 31944 13456 31996 13462
rect 31944 13398 31996 13404
rect 32312 13320 32364 13326
rect 32312 13262 32364 13268
rect 32324 12986 32352 13262
rect 32496 13184 32548 13190
rect 32496 13126 32548 13132
rect 32312 12980 32364 12986
rect 32312 12922 32364 12928
rect 32508 12850 32536 13126
rect 32496 12844 32548 12850
rect 32496 12786 32548 12792
rect 30840 12300 30892 12306
rect 30840 12242 30892 12248
rect 34532 11762 34560 14962
rect 35440 14884 35492 14890
rect 35440 14826 35492 14832
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34520 11756 34572 11762
rect 34520 11698 34572 11704
rect 31668 5024 31720 5030
rect 31668 4966 31720 4972
rect 31680 3534 31708 4966
rect 31668 3528 31720 3534
rect 31668 3470 31720 3476
rect 30564 3460 30616 3466
rect 30564 3402 30616 3408
rect 33784 3392 33836 3398
rect 33784 3334 33836 3340
rect 30288 2644 30340 2650
rect 30288 2586 30340 2592
rect 25596 2576 25648 2582
rect 25596 2518 25648 2524
rect 27528 2576 27580 2582
rect 27528 2518 27580 2524
rect 33796 2446 33824 3334
rect 34532 2582 34560 11698
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34796 3936 34848 3942
rect 34796 3878 34848 3884
rect 34520 2576 34572 2582
rect 34520 2518 34572 2524
rect 34808 2514 34836 3878
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35452 3194 35480 14826
rect 36004 8974 36032 22986
rect 37188 20936 37240 20942
rect 37188 20878 37240 20884
rect 37200 20505 37228 20878
rect 37186 20496 37242 20505
rect 37186 20431 37242 20440
rect 36912 16108 36964 16114
rect 36912 16050 36964 16056
rect 36924 15162 36952 16050
rect 37292 15366 37320 36110
rect 37384 35086 37412 39200
rect 38106 37496 38162 37505
rect 38106 37431 38162 37440
rect 37924 37324 37976 37330
rect 37924 37266 37976 37272
rect 37372 35080 37424 35086
rect 37372 35022 37424 35028
rect 37464 34944 37516 34950
rect 37464 34886 37516 34892
rect 37476 29782 37504 34886
rect 37464 29776 37516 29782
rect 37464 29718 37516 29724
rect 37464 29640 37516 29646
rect 37464 29582 37516 29588
rect 37476 29345 37504 29582
rect 37462 29336 37518 29345
rect 37462 29271 37518 29280
rect 37832 21548 37884 21554
rect 37832 21490 37884 21496
rect 37740 20936 37792 20942
rect 37740 20878 37792 20884
rect 37752 16046 37780 20878
rect 37740 16040 37792 16046
rect 37740 15982 37792 15988
rect 37280 15360 37332 15366
rect 37280 15302 37332 15308
rect 36912 15156 36964 15162
rect 36912 15098 36964 15104
rect 37752 15026 37780 15982
rect 37740 15020 37792 15026
rect 37740 14962 37792 14968
rect 37096 14952 37148 14958
rect 37096 14894 37148 14900
rect 36912 13932 36964 13938
rect 36912 13874 36964 13880
rect 35992 8968 36044 8974
rect 35992 8910 36044 8916
rect 36452 8832 36504 8838
rect 36452 8774 36504 8780
rect 36464 8498 36492 8774
rect 36924 8634 36952 13874
rect 37108 11354 37136 14894
rect 37740 13252 37792 13258
rect 37740 13194 37792 13200
rect 37096 11348 37148 11354
rect 37096 11290 37148 11296
rect 37188 10056 37240 10062
rect 37188 9998 37240 10004
rect 37200 9625 37228 9998
rect 37186 9616 37242 9625
rect 37186 9551 37242 9560
rect 37188 9512 37240 9518
rect 37188 9454 37240 9460
rect 36912 8628 36964 8634
rect 36912 8570 36964 8576
rect 36452 8492 36504 8498
rect 36452 8434 36504 8440
rect 36360 7744 36412 7750
rect 36360 7686 36412 7692
rect 36372 4146 36400 7686
rect 37200 4826 37228 9454
rect 37188 4820 37240 4826
rect 37188 4762 37240 4768
rect 37188 4208 37240 4214
rect 37188 4150 37240 4156
rect 36360 4140 36412 4146
rect 36360 4082 36412 4088
rect 35440 3188 35492 3194
rect 35440 3130 35492 3136
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34796 2508 34848 2514
rect 34796 2450 34848 2456
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 31576 2440 31628 2446
rect 31576 2382 31628 2388
rect 33784 2440 33836 2446
rect 33784 2382 33836 2388
rect 36728 2440 36780 2446
rect 36728 2382 36780 2388
rect 25044 2304 25096 2310
rect 25044 2246 25096 2252
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 25780 2304 25832 2310
rect 25780 2246 25832 2252
rect 24400 2100 24452 2106
rect 24400 2042 24452 2048
rect 25148 800 25176 2246
rect 25792 800 25820 2246
rect 27080 800 27108 2382
rect 28368 800 28396 2382
rect 29828 2372 29880 2378
rect 29828 2314 29880 2320
rect 29644 2304 29696 2310
rect 29644 2246 29696 2252
rect 29656 800 29684 2246
rect 29840 2106 29868 2314
rect 29828 2100 29880 2106
rect 29828 2042 29880 2048
rect 30300 800 30328 2382
rect 31588 800 31616 2382
rect 32864 2372 32916 2378
rect 32864 2314 32916 2320
rect 32876 800 32904 2314
rect 33508 2304 33560 2310
rect 33508 2246 33560 2252
rect 34796 2304 34848 2310
rect 34796 2246 34848 2252
rect 36084 2304 36136 2310
rect 36084 2246 36136 2252
rect 33520 800 33548 2246
rect 34808 800 34836 2246
rect 36096 800 36124 2246
rect 36740 800 36768 2382
rect 37200 1465 37228 4150
rect 37464 3392 37516 3398
rect 37464 3334 37516 3340
rect 37476 3126 37504 3334
rect 37464 3120 37516 3126
rect 37464 3062 37516 3068
rect 37280 3052 37332 3058
rect 37280 2994 37332 3000
rect 37186 1456 37242 1465
rect 37186 1391 37242 1400
rect 2778 776 2834 785
rect 2778 711 2834 720
rect 3238 200 3294 800
rect 3882 200 3938 800
rect 5170 200 5226 800
rect 6458 200 6514 800
rect 7102 200 7158 800
rect 8390 200 8446 800
rect 9678 200 9734 800
rect 10966 200 11022 800
rect 11610 200 11666 800
rect 12898 200 12954 800
rect 14186 200 14242 800
rect 14830 200 14886 800
rect 16118 200 16174 800
rect 17406 200 17462 800
rect 18050 200 18106 800
rect 19338 200 19394 800
rect 20626 200 20682 800
rect 21914 200 21970 800
rect 22558 200 22614 800
rect 23846 200 23902 800
rect 25134 200 25190 800
rect 25778 200 25834 800
rect 27066 200 27122 800
rect 28354 200 28410 800
rect 29642 200 29698 800
rect 30286 200 30342 800
rect 31574 200 31630 800
rect 32862 200 32918 800
rect 33506 200 33562 800
rect 34794 200 34850 800
rect 36082 200 36138 800
rect 36726 200 36782 800
rect 37292 785 37320 2994
rect 37752 2514 37780 13194
rect 37844 11286 37872 21490
rect 37936 18222 37964 37266
rect 38120 37262 38148 37431
rect 38108 37256 38160 37262
rect 38108 37198 38160 37204
rect 38672 36854 38700 39200
rect 39316 36922 39344 39200
rect 39304 36916 39356 36922
rect 39304 36858 39356 36864
rect 38660 36848 38712 36854
rect 38660 36790 38712 36796
rect 38200 36576 38252 36582
rect 38200 36518 38252 36524
rect 38212 36310 38240 36518
rect 38200 36304 38252 36310
rect 38200 36246 38252 36252
rect 38198 36136 38254 36145
rect 38198 36071 38254 36080
rect 38212 36038 38240 36071
rect 38200 36032 38252 36038
rect 38200 35974 38252 35980
rect 38016 35692 38068 35698
rect 38016 35634 38068 35640
rect 38028 31142 38056 35634
rect 38200 35488 38252 35494
rect 38198 35456 38200 35465
rect 38252 35456 38254 35465
rect 38198 35391 38254 35400
rect 38200 34400 38252 34406
rect 38200 34342 38252 34348
rect 38212 34105 38240 34342
rect 38198 34096 38254 34105
rect 38198 34031 38254 34040
rect 38200 32768 38252 32774
rect 38198 32736 38200 32745
rect 38252 32736 38254 32745
rect 38198 32671 38254 32680
rect 38200 32224 38252 32230
rect 38200 32166 38252 32172
rect 38212 32065 38240 32166
rect 38198 32056 38254 32065
rect 38198 31991 38254 32000
rect 38016 31136 38068 31142
rect 38016 31078 38068 31084
rect 38292 30728 38344 30734
rect 38290 30696 38292 30705
rect 38344 30696 38346 30705
rect 38290 30631 38346 30640
rect 38108 30592 38160 30598
rect 38108 30534 38160 30540
rect 38120 28626 38148 30534
rect 38108 28620 38160 28626
rect 38108 28562 38160 28568
rect 38292 28076 38344 28082
rect 38292 28018 38344 28024
rect 38304 27985 38332 28018
rect 38290 27976 38346 27985
rect 38290 27911 38346 27920
rect 38016 27464 38068 27470
rect 38016 27406 38068 27412
rect 38028 21690 38056 27406
rect 38200 27328 38252 27334
rect 38198 27296 38200 27305
rect 38252 27296 38254 27305
rect 38198 27231 38254 27240
rect 38108 26920 38160 26926
rect 38108 26862 38160 26868
rect 38120 26586 38148 26862
rect 38108 26580 38160 26586
rect 38108 26522 38160 26528
rect 38292 26376 38344 26382
rect 38292 26318 38344 26324
rect 38304 25945 38332 26318
rect 38290 25936 38346 25945
rect 38290 25871 38346 25880
rect 38200 24608 38252 24614
rect 38198 24576 38200 24585
rect 38252 24576 38254 24585
rect 38198 24511 38254 24520
rect 38200 24064 38252 24070
rect 38200 24006 38252 24012
rect 38212 23905 38240 24006
rect 38198 23896 38254 23905
rect 38198 23831 38254 23840
rect 38198 22536 38254 22545
rect 38198 22471 38200 22480
rect 38252 22471 38254 22480
rect 38200 22442 38252 22448
rect 38016 21684 38068 21690
rect 38016 21626 38068 21632
rect 38200 21344 38252 21350
rect 38200 21286 38252 21292
rect 38212 21185 38240 21286
rect 38198 21176 38254 21185
rect 38198 21111 38254 21120
rect 38108 21072 38160 21078
rect 38108 21014 38160 21020
rect 38120 19514 38148 21014
rect 38108 19508 38160 19514
rect 38108 19450 38160 19456
rect 38292 19372 38344 19378
rect 38292 19314 38344 19320
rect 38304 19145 38332 19314
rect 38290 19136 38346 19145
rect 38290 19071 38346 19080
rect 37924 18216 37976 18222
rect 37924 18158 37976 18164
rect 38200 18080 38252 18086
rect 38200 18022 38252 18028
rect 38212 17785 38240 18022
rect 38198 17776 38254 17785
rect 38198 17711 38254 17720
rect 38016 16584 38068 16590
rect 38016 16526 38068 16532
rect 38028 15910 38056 16526
rect 38200 16448 38252 16454
rect 38198 16416 38200 16425
rect 38252 16416 38254 16425
rect 38198 16351 38254 16360
rect 38016 15904 38068 15910
rect 38016 15846 38068 15852
rect 38200 15904 38252 15910
rect 38200 15846 38252 15852
rect 38212 15745 38240 15846
rect 38198 15736 38254 15745
rect 38198 15671 38254 15680
rect 37924 14816 37976 14822
rect 37924 14758 37976 14764
rect 37832 11280 37884 11286
rect 37832 11222 37884 11228
rect 37936 3534 37964 14758
rect 38198 14376 38254 14385
rect 38198 14311 38254 14320
rect 38212 14278 38240 14311
rect 38200 14272 38252 14278
rect 38200 14214 38252 14220
rect 38200 13184 38252 13190
rect 38200 13126 38252 13132
rect 38212 13025 38240 13126
rect 38198 13016 38254 13025
rect 38198 12951 38254 12960
rect 38292 12844 38344 12850
rect 38292 12786 38344 12792
rect 38304 12345 38332 12786
rect 38290 12336 38346 12345
rect 38290 12271 38346 12280
rect 38292 11144 38344 11150
rect 38292 11086 38344 11092
rect 38304 10985 38332 11086
rect 38290 10976 38346 10985
rect 38290 10911 38346 10920
rect 38292 8492 38344 8498
rect 38292 8434 38344 8440
rect 38016 8356 38068 8362
rect 38016 8298 38068 8304
rect 38028 5234 38056 8298
rect 38304 8265 38332 8434
rect 38290 8256 38346 8265
rect 38290 8191 38346 8200
rect 38292 7880 38344 7886
rect 38292 7822 38344 7828
rect 38304 7585 38332 7822
rect 38290 7576 38346 7585
rect 38290 7511 38346 7520
rect 38292 6316 38344 6322
rect 38292 6258 38344 6264
rect 38304 6225 38332 6258
rect 38290 6216 38346 6225
rect 38290 6151 38346 6160
rect 38016 5228 38068 5234
rect 38016 5170 38068 5176
rect 38200 5024 38252 5030
rect 38200 4966 38252 4972
rect 38212 4865 38240 4966
rect 38198 4856 38254 4865
rect 38198 4791 38254 4800
rect 38292 4616 38344 4622
rect 38292 4558 38344 4564
rect 38304 4185 38332 4558
rect 38290 4176 38346 4185
rect 38290 4111 38346 4120
rect 37924 3528 37976 3534
rect 37924 3470 37976 3476
rect 38016 3392 38068 3398
rect 38016 3334 38068 3340
rect 38200 3392 38252 3398
rect 38200 3334 38252 3340
rect 37740 2508 37792 2514
rect 37740 2450 37792 2456
rect 38028 800 38056 3334
rect 38212 2825 38240 3334
rect 39304 3052 39356 3058
rect 39304 2994 39356 3000
rect 38198 2816 38254 2825
rect 38198 2751 38254 2760
rect 39316 800 39344 2994
rect 37278 776 37334 785
rect 37278 711 37334 720
rect 38014 200 38070 800
rect 39302 200 39358 800
<< via2 >>
rect 1582 38800 1638 38856
rect 1766 38120 1822 38176
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 1582 36352 1638 36408
rect 1766 35400 1822 35456
rect 1766 34720 1822 34776
rect 2410 34040 2466 34096
rect 1766 33360 1822 33416
rect 1674 32000 1730 32056
rect 1766 31320 1822 31376
rect 1766 29996 1768 30016
rect 1768 29996 1820 30016
rect 1820 29996 1822 30016
rect 1766 29960 1822 29996
rect 1582 29008 1638 29064
rect 1766 28600 1822 28656
rect 1766 27276 1768 27296
rect 1768 27276 1820 27296
rect 1820 27276 1822 27296
rect 1766 27240 1822 27276
rect 1766 26560 1822 26616
rect 1582 26288 1638 26344
rect 1674 25236 1676 25256
rect 1676 25236 1728 25256
rect 1728 25236 1730 25256
rect 1674 25200 1730 25236
rect 1766 23840 1822 23896
rect 1674 21800 1730 21856
rect 1674 20440 1730 20496
rect 1766 19080 1822 19136
rect 1674 18400 1730 18456
rect 1674 17040 1730 17096
rect 1766 15680 1822 15736
rect 1674 13640 1730 13696
rect 1766 12316 1768 12336
rect 1768 12316 1820 12336
rect 1820 12316 1822 12336
rect 1766 12280 1822 12316
rect 1766 8880 1822 8936
rect 1766 7520 1822 7576
rect 2410 31764 2412 31784
rect 2412 31764 2464 31784
rect 2464 31764 2466 31784
rect 2410 31728 2466 31764
rect 3330 36760 3386 36816
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4066 33532 4068 33552
rect 4068 33532 4120 33552
rect 4120 33532 4122 33552
rect 4066 33496 4122 33532
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4894 34856 4950 34912
rect 2226 15952 2282 16008
rect 2502 15000 2558 15056
rect 2318 11872 2374 11928
rect 2778 23160 2834 23216
rect 2870 15000 2926 15056
rect 3422 19352 3478 19408
rect 2778 14320 2834 14376
rect 2686 13776 2742 13832
rect 2042 9152 2098 9208
rect 1766 6840 1822 6896
rect 1950 6452 2006 6488
rect 1950 6432 1952 6452
rect 1952 6432 2004 6452
rect 2004 6432 2006 6452
rect 2042 5888 2098 5944
rect 3514 18128 3570 18184
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4066 29180 4068 29200
rect 4068 29180 4120 29200
rect 4120 29180 4122 29200
rect 4066 29144 4122 29180
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 7378 35944 7434 36000
rect 8206 35536 8262 35592
rect 5906 33924 5962 33960
rect 5906 33904 5908 33924
rect 5908 33904 5960 33924
rect 5960 33904 5962 33924
rect 5354 31356 5356 31376
rect 5356 31356 5408 31376
rect 5408 31356 5410 31376
rect 5354 31320 5410 31356
rect 5354 30676 5356 30696
rect 5356 30676 5408 30696
rect 5408 30676 5410 30696
rect 5354 30640 5410 30676
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 3606 17720 3662 17776
rect 4986 27648 5042 27704
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4526 23568 4582 23624
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 5078 26308 5134 26344
rect 5078 26288 5080 26308
rect 5080 26288 5132 26308
rect 5132 26288 5134 26308
rect 4710 16088 4766 16144
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 3606 11600 3662 11656
rect 3054 9580 3110 9616
rect 3054 9560 3056 9580
rect 3056 9560 3108 9580
rect 3108 9560 3110 9580
rect 3146 9424 3202 9480
rect 3422 10240 3478 10296
rect 3606 9560 3662 9616
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4894 15000 4950 15056
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 5354 22072 5410 22128
rect 5170 18808 5226 18864
rect 6458 28484 6514 28520
rect 6458 28464 6460 28484
rect 6460 28464 6512 28484
rect 6512 28464 6514 28484
rect 7010 26288 7066 26344
rect 5998 22380 6000 22400
rect 6000 22380 6052 22400
rect 6052 22380 6054 22400
rect 5998 22344 6054 22380
rect 5262 15816 5318 15872
rect 5538 16088 5594 16144
rect 5446 15408 5502 15464
rect 5446 13640 5502 13696
rect 5538 12280 5594 12336
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 5630 10920 5686 10976
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 1766 5480 1822 5536
rect 1766 4120 1822 4176
rect 1398 3440 1454 3496
rect 3146 3188 3202 3224
rect 3146 3168 3148 3188
rect 3148 3168 3200 3188
rect 3200 3168 3202 3188
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 6918 15444 6920 15464
rect 6920 15444 6972 15464
rect 6972 15444 6974 15464
rect 6918 15408 6974 15444
rect 7654 17856 7710 17912
rect 7838 18128 7894 18184
rect 11978 37324 12034 37360
rect 11978 37304 11980 37324
rect 11980 37304 12032 37324
rect 12032 37304 12034 37324
rect 8942 34992 8998 35048
rect 9310 35012 9366 35048
rect 9310 34992 9312 35012
rect 9312 34992 9364 35012
rect 9364 34992 9366 35012
rect 9218 34892 9220 34912
rect 9220 34892 9272 34912
rect 9272 34892 9274 34912
rect 9218 34856 9274 34892
rect 8666 25100 8668 25120
rect 8668 25100 8720 25120
rect 8720 25100 8722 25120
rect 8666 25064 8722 25100
rect 10046 36488 10102 36544
rect 13358 36896 13414 36952
rect 12806 36352 12862 36408
rect 11610 35808 11666 35864
rect 11058 34448 11114 34504
rect 11426 35536 11482 35592
rect 12990 35672 13046 35728
rect 11610 34584 11666 34640
rect 12070 34992 12126 35048
rect 13358 34312 13414 34368
rect 12254 34176 12310 34232
rect 11610 33088 11666 33144
rect 9310 15816 9366 15872
rect 8114 13640 8170 13696
rect 9494 13640 9550 13696
rect 8206 11736 8262 11792
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 1674 2080 1730 2136
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 9770 15136 9826 15192
rect 9770 13776 9826 13832
rect 11886 33768 11942 33824
rect 12622 33632 12678 33688
rect 11886 32408 11942 32464
rect 11058 22888 11114 22944
rect 12990 32680 13046 32736
rect 12254 31864 12310 31920
rect 12346 29008 12402 29064
rect 14002 36216 14058 36272
rect 13634 35128 13690 35184
rect 13726 32952 13782 33008
rect 13910 31864 13966 31920
rect 13634 30912 13690 30968
rect 11426 25744 11482 25800
rect 10414 15952 10470 16008
rect 11242 13812 11244 13832
rect 11244 13812 11296 13832
rect 11296 13812 11298 13832
rect 11242 13776 11298 13812
rect 11702 14728 11758 14784
rect 12806 23060 12808 23080
rect 12808 23060 12860 23080
rect 12860 23060 12862 23080
rect 12806 23024 12862 23060
rect 12070 14728 12126 14784
rect 13910 30776 13966 30832
rect 14370 32272 14426 32328
rect 14738 35536 14794 35592
rect 14554 29416 14610 29472
rect 14094 28872 14150 28928
rect 13634 27648 13690 27704
rect 13082 16088 13138 16144
rect 15014 36116 15016 36136
rect 15016 36116 15068 36136
rect 15068 36116 15070 36136
rect 15014 36080 15070 36116
rect 15382 36796 15384 36816
rect 15384 36796 15436 36816
rect 15436 36796 15438 36816
rect 15382 36760 15438 36796
rect 15290 34196 15346 34232
rect 15290 34176 15292 34196
rect 15292 34176 15344 34196
rect 15344 34176 15346 34196
rect 14922 32816 14978 32872
rect 15934 35264 15990 35320
rect 15474 34856 15530 34912
rect 16210 35944 16266 36000
rect 16118 34856 16174 34912
rect 16026 34720 16082 34776
rect 15566 34176 15622 34232
rect 15842 33396 15844 33416
rect 15844 33396 15896 33416
rect 15896 33396 15898 33416
rect 15842 33360 15898 33396
rect 15566 33224 15622 33280
rect 15474 32272 15530 32328
rect 16210 33224 16266 33280
rect 14738 28736 14794 28792
rect 15014 27512 15070 27568
rect 15014 26288 15070 26344
rect 13634 14320 13690 14376
rect 14186 17196 14242 17232
rect 14186 17176 14188 17196
rect 14188 17176 14240 17196
rect 14240 17176 14242 17196
rect 15290 30252 15346 30288
rect 15290 30232 15292 30252
rect 15292 30232 15344 30252
rect 15344 30232 15346 30252
rect 15474 24656 15530 24712
rect 15014 18264 15070 18320
rect 18510 36916 18566 36952
rect 18510 36896 18512 36916
rect 18512 36896 18564 36916
rect 18564 36896 18566 36916
rect 17406 35944 17462 36000
rect 17130 34992 17186 35048
rect 18510 36116 18512 36136
rect 18512 36116 18564 36136
rect 18564 36116 18566 36136
rect 18510 36080 18566 36116
rect 17498 33632 17554 33688
rect 17314 32816 17370 32872
rect 16210 28328 16266 28384
rect 15474 15444 15476 15464
rect 15476 15444 15528 15464
rect 15528 15444 15530 15464
rect 15474 15408 15530 15444
rect 15198 13776 15254 13832
rect 15934 8880 15990 8936
rect 16854 23568 16910 23624
rect 18050 34720 18106 34776
rect 17866 31884 17922 31920
rect 17866 31864 17868 31884
rect 17868 31864 17920 31884
rect 17920 31864 17922 31884
rect 18510 34312 18566 34368
rect 18418 31864 18474 31920
rect 17406 30232 17462 30288
rect 17222 29416 17278 29472
rect 17314 28756 17370 28792
rect 17314 28736 17316 28756
rect 17316 28736 17368 28756
rect 17368 28736 17370 28756
rect 17222 26424 17278 26480
rect 17130 24520 17186 24576
rect 17682 29824 17738 29880
rect 17406 25880 17462 25936
rect 17406 24676 17462 24712
rect 17406 24656 17408 24676
rect 17408 24656 17460 24676
rect 17460 24656 17462 24676
rect 17774 26308 17830 26344
rect 17774 26288 17776 26308
rect 17776 26288 17828 26308
rect 17828 26288 17830 26308
rect 18142 29008 18198 29064
rect 18234 28328 18290 28384
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19338 35808 19394 35864
rect 18878 33496 18934 33552
rect 18786 31220 18788 31240
rect 18788 31220 18840 31240
rect 18840 31220 18842 31240
rect 18786 31184 18842 31220
rect 18694 30776 18750 30832
rect 17406 23044 17462 23080
rect 17406 23024 17408 23044
rect 17408 23024 17460 23044
rect 17460 23024 17462 23044
rect 17222 17212 17224 17232
rect 17224 17212 17276 17232
rect 17276 17212 17278 17232
rect 17222 17176 17278 17212
rect 17038 15444 17040 15464
rect 17040 15444 17092 15464
rect 17092 15444 17094 15464
rect 17038 15408 17094 15444
rect 17774 22516 17776 22536
rect 17776 22516 17828 22536
rect 17828 22516 17830 22536
rect 17774 22480 17830 22516
rect 18050 24520 18106 24576
rect 20350 37168 20406 37224
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19706 35400 19762 35456
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 20074 35944 20130 36000
rect 20718 36488 20774 36544
rect 20074 34856 20130 34912
rect 19154 33768 19210 33824
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19522 33496 19578 33552
rect 19154 31728 19210 31784
rect 19062 29280 19118 29336
rect 19706 33360 19762 33416
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19614 32136 19670 32192
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 20258 32308 20260 32328
rect 20260 32308 20312 32328
rect 20312 32308 20314 32328
rect 20258 32272 20314 32308
rect 19614 30776 19670 30832
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 20442 34992 20498 35048
rect 20718 34584 20774 34640
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19982 29280 20038 29336
rect 18970 29008 19026 29064
rect 17774 18264 17830 18320
rect 18970 26288 19026 26344
rect 19154 25744 19210 25800
rect 19154 22072 19210 22128
rect 19522 29008 19578 29064
rect 20258 29416 20314 29472
rect 20350 29280 20406 29336
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19798 27396 19854 27432
rect 19798 27376 19800 27396
rect 19800 27376 19852 27396
rect 19852 27376 19854 27396
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19430 26988 19486 27024
rect 19430 26968 19432 26988
rect 19432 26968 19484 26988
rect 19484 26968 19486 26988
rect 20074 28736 20130 28792
rect 19982 26832 20038 26888
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 20534 32972 20590 33008
rect 20534 32952 20536 32972
rect 20536 32952 20588 32972
rect 20588 32952 20590 32972
rect 20902 35128 20958 35184
rect 20626 30776 20682 30832
rect 20534 28600 20590 28656
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19982 24812 20038 24848
rect 19982 24792 19984 24812
rect 19984 24792 20036 24812
rect 20036 24792 20038 24812
rect 18970 16088 19026 16144
rect 19246 14476 19302 14512
rect 19246 14456 19248 14476
rect 19248 14456 19300 14476
rect 19300 14456 19302 14476
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19982 20440 20038 20496
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19890 18300 19892 18320
rect 19892 18300 19944 18320
rect 19944 18300 19946 18320
rect 19890 18264 19946 18300
rect 19890 18148 19946 18184
rect 19890 18128 19892 18148
rect 19892 18128 19944 18148
rect 19944 18128 19946 18148
rect 19890 17756 19892 17776
rect 19892 17756 19944 17776
rect 19944 17756 19946 17776
rect 19890 17720 19946 17756
rect 20902 31320 20958 31376
rect 21454 37204 21456 37224
rect 21456 37204 21508 37224
rect 21508 37204 21510 37224
rect 21454 37168 21510 37204
rect 21362 36100 21418 36136
rect 21362 36080 21364 36100
rect 21364 36080 21416 36100
rect 21416 36080 21418 36100
rect 21270 35556 21326 35592
rect 21270 35536 21272 35556
rect 21272 35536 21324 35556
rect 21324 35536 21326 35556
rect 21270 34448 21326 34504
rect 20902 28464 20958 28520
rect 21086 28872 21142 28928
rect 20902 27512 20958 27568
rect 20626 24928 20682 24984
rect 21086 26308 21142 26344
rect 21086 26288 21088 26308
rect 21088 26288 21140 26308
rect 21140 26288 21142 26308
rect 21822 36352 21878 36408
rect 22098 36216 22154 36272
rect 22006 32952 22062 33008
rect 21914 32136 21970 32192
rect 22282 30640 22338 30696
rect 22466 29144 22522 29200
rect 22190 29008 22246 29064
rect 21638 28600 21694 28656
rect 21822 28600 21878 28656
rect 21454 27648 21510 27704
rect 21914 28192 21970 28248
rect 20994 24520 21050 24576
rect 20534 22208 20590 22264
rect 19614 17604 19670 17640
rect 19614 17584 19616 17604
rect 19616 17584 19668 17604
rect 19668 17584 19670 17604
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19430 9596 19432 9616
rect 19432 9596 19484 9616
rect 19484 9596 19486 9616
rect 19430 9560 19486 9596
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 20166 9580 20222 9616
rect 20166 9560 20168 9580
rect 20168 9560 20220 9580
rect 20220 9560 20222 9580
rect 21638 25900 21694 25936
rect 21638 25880 21640 25900
rect 21640 25880 21692 25900
rect 21692 25880 21694 25900
rect 21546 24792 21602 24848
rect 21730 24656 21786 24712
rect 21730 24112 21786 24168
rect 21914 27532 21970 27568
rect 21914 27512 21916 27532
rect 21916 27512 21968 27532
rect 21968 27512 21970 27532
rect 22190 27548 22192 27568
rect 22192 27548 22244 27568
rect 22244 27548 22246 27568
rect 22190 27512 22246 27548
rect 21914 24112 21970 24168
rect 21822 23568 21878 23624
rect 22006 23432 22062 23488
rect 21638 22072 21694 22128
rect 21178 17584 21234 17640
rect 21362 14456 21418 14512
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 22282 23432 22338 23488
rect 22742 33516 22798 33552
rect 22742 33496 22744 33516
rect 22744 33496 22796 33516
rect 22796 33496 22798 33516
rect 23294 35264 23350 35320
rect 23110 34856 23166 34912
rect 23110 30912 23166 30968
rect 22558 23568 22614 23624
rect 22098 19760 22154 19816
rect 23110 26424 23166 26480
rect 23570 28600 23626 28656
rect 22926 18128 22982 18184
rect 22742 14320 22798 14376
rect 25226 36796 25228 36816
rect 25228 36796 25280 36816
rect 25280 36796 25282 36816
rect 25226 36760 25282 36796
rect 25042 36216 25098 36272
rect 25410 35708 25412 35728
rect 25412 35708 25464 35728
rect 25464 35708 25466 35728
rect 25410 35672 25466 35708
rect 23846 34040 23902 34096
rect 23938 33904 23994 33960
rect 24582 32852 24584 32872
rect 24584 32852 24636 32872
rect 24636 32852 24638 32872
rect 24582 32816 24638 32852
rect 24030 24656 24086 24712
rect 24306 27376 24362 27432
rect 24766 29824 24822 29880
rect 25318 35400 25374 35456
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 25778 33224 25834 33280
rect 24858 29144 24914 29200
rect 24950 28212 25006 28248
rect 24950 28192 24952 28212
rect 24952 28192 25004 28212
rect 25004 28192 25006 28212
rect 23570 19216 23626 19272
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 24582 17720 24638 17776
rect 25686 31884 25742 31920
rect 25686 31864 25688 31884
rect 25688 31864 25740 31884
rect 25740 31864 25742 31884
rect 26238 33088 26294 33144
rect 25594 14340 25650 14376
rect 25594 14320 25596 14340
rect 25596 14320 25648 14340
rect 25648 14320 25650 14340
rect 26422 28736 26478 28792
rect 26790 29144 26846 29200
rect 27250 34176 27306 34232
rect 27618 31884 27674 31920
rect 27618 31864 27620 31884
rect 27620 31864 27672 31884
rect 27672 31864 27674 31884
rect 26606 26968 26662 27024
rect 28354 32408 28410 32464
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 37186 38800 37242 38856
rect 28354 18264 28410 18320
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 30930 22616 30986 22672
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 37186 20440 37242 20496
rect 38106 37440 38162 37496
rect 37462 29280 37518 29336
rect 37186 9560 37242 9616
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 37186 1400 37242 1456
rect 2778 720 2834 776
rect 38198 36080 38254 36136
rect 38198 35436 38200 35456
rect 38200 35436 38252 35456
rect 38252 35436 38254 35456
rect 38198 35400 38254 35436
rect 38198 34040 38254 34096
rect 38198 32716 38200 32736
rect 38200 32716 38252 32736
rect 38252 32716 38254 32736
rect 38198 32680 38254 32716
rect 38198 32000 38254 32056
rect 38290 30676 38292 30696
rect 38292 30676 38344 30696
rect 38344 30676 38346 30696
rect 38290 30640 38346 30676
rect 38290 27920 38346 27976
rect 38198 27276 38200 27296
rect 38200 27276 38252 27296
rect 38252 27276 38254 27296
rect 38198 27240 38254 27276
rect 38290 25880 38346 25936
rect 38198 24556 38200 24576
rect 38200 24556 38252 24576
rect 38252 24556 38254 24576
rect 38198 24520 38254 24556
rect 38198 23840 38254 23896
rect 38198 22500 38254 22536
rect 38198 22480 38200 22500
rect 38200 22480 38252 22500
rect 38252 22480 38254 22500
rect 38198 21120 38254 21176
rect 38290 19080 38346 19136
rect 38198 17720 38254 17776
rect 38198 16396 38200 16416
rect 38200 16396 38252 16416
rect 38252 16396 38254 16416
rect 38198 16360 38254 16396
rect 38198 15680 38254 15736
rect 38198 14320 38254 14376
rect 38198 12960 38254 13016
rect 38290 12280 38346 12336
rect 38290 10920 38346 10976
rect 38290 8200 38346 8256
rect 38290 7520 38346 7576
rect 38290 6160 38346 6216
rect 38198 4800 38254 4856
rect 38290 4120 38346 4176
rect 38198 2760 38254 2816
rect 37278 720 37334 776
<< metal3 >>
rect 200 38858 800 38888
rect 1577 38858 1643 38861
rect 200 38856 1643 38858
rect 200 38800 1582 38856
rect 1638 38800 1643 38856
rect 200 38798 1643 38800
rect 200 38768 800 38798
rect 1577 38795 1643 38798
rect 37181 38858 37247 38861
rect 39200 38858 39800 38888
rect 37181 38856 39800 38858
rect 37181 38800 37186 38856
rect 37242 38800 39800 38856
rect 37181 38798 39800 38800
rect 37181 38795 37247 38798
rect 39200 38768 39800 38798
rect 200 38178 800 38208
rect 1761 38178 1827 38181
rect 200 38176 1827 38178
rect 200 38120 1766 38176
rect 1822 38120 1827 38176
rect 200 38118 1827 38120
rect 200 38088 800 38118
rect 1761 38115 1827 38118
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 38101 37498 38167 37501
rect 39200 37498 39800 37528
rect 38101 37496 39800 37498
rect 38101 37440 38106 37496
rect 38162 37440 39800 37496
rect 38101 37438 39800 37440
rect 38101 37435 38167 37438
rect 39200 37408 39800 37438
rect 11973 37364 12039 37365
rect 11973 37362 12020 37364
rect 11892 37360 12020 37362
rect 12084 37362 12090 37364
rect 20662 37362 20668 37364
rect 11892 37304 11978 37360
rect 11892 37302 12020 37304
rect 11973 37300 12020 37302
rect 12084 37302 20668 37362
rect 12084 37300 12090 37302
rect 20662 37300 20668 37302
rect 20732 37300 20738 37364
rect 11973 37299 12039 37300
rect 20345 37226 20411 37229
rect 21449 37226 21515 37229
rect 20345 37224 21515 37226
rect 20345 37168 20350 37224
rect 20406 37168 21454 37224
rect 21510 37168 21515 37224
rect 20345 37166 21515 37168
rect 20345 37163 20411 37166
rect 21449 37163 21515 37166
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 13353 36954 13419 36957
rect 18505 36954 18571 36957
rect 13353 36952 18571 36954
rect 13353 36896 13358 36952
rect 13414 36896 18510 36952
rect 18566 36896 18571 36952
rect 13353 36894 18571 36896
rect 13353 36891 13419 36894
rect 18505 36891 18571 36894
rect 200 36818 800 36848
rect 3325 36818 3391 36821
rect 200 36816 3391 36818
rect 200 36760 3330 36816
rect 3386 36760 3391 36816
rect 200 36758 3391 36760
rect 200 36728 800 36758
rect 3325 36755 3391 36758
rect 15377 36818 15443 36821
rect 25221 36818 25287 36821
rect 15377 36816 25287 36818
rect 15377 36760 15382 36816
rect 15438 36760 25226 36816
rect 25282 36760 25287 36816
rect 15377 36758 25287 36760
rect 15377 36755 15443 36758
rect 25221 36755 25287 36758
rect 10041 36546 10107 36549
rect 20713 36546 20779 36549
rect 10041 36544 20779 36546
rect 10041 36488 10046 36544
rect 10102 36488 20718 36544
rect 20774 36488 20779 36544
rect 10041 36486 20779 36488
rect 10041 36483 10107 36486
rect 20713 36483 20779 36486
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 1577 36410 1643 36413
rect 2078 36410 2084 36412
rect 1577 36408 2084 36410
rect 1577 36352 1582 36408
rect 1638 36352 2084 36408
rect 1577 36350 2084 36352
rect 1577 36347 1643 36350
rect 2078 36348 2084 36350
rect 2148 36348 2154 36412
rect 12801 36410 12867 36413
rect 21817 36410 21883 36413
rect 12801 36408 21883 36410
rect 12801 36352 12806 36408
rect 12862 36352 21822 36408
rect 21878 36352 21883 36408
rect 12801 36350 21883 36352
rect 12801 36347 12867 36350
rect 21817 36347 21883 36350
rect 13997 36274 14063 36277
rect 22093 36274 22159 36277
rect 25037 36274 25103 36277
rect 13997 36272 25103 36274
rect 13997 36216 14002 36272
rect 14058 36216 22098 36272
rect 22154 36216 25042 36272
rect 25098 36216 25103 36272
rect 13997 36214 25103 36216
rect 13997 36211 14063 36214
rect 22093 36211 22159 36214
rect 25037 36211 25103 36214
rect 15009 36138 15075 36141
rect 18505 36138 18571 36141
rect 15009 36136 18571 36138
rect 15009 36080 15014 36136
rect 15070 36080 18510 36136
rect 18566 36080 18571 36136
rect 15009 36078 18571 36080
rect 15009 36075 15075 36078
rect 18505 36075 18571 36078
rect 19374 36076 19380 36140
rect 19444 36138 19450 36140
rect 21357 36138 21423 36141
rect 19444 36136 21423 36138
rect 19444 36080 21362 36136
rect 21418 36080 21423 36136
rect 19444 36078 21423 36080
rect 19444 36076 19450 36078
rect 21357 36075 21423 36078
rect 38193 36138 38259 36141
rect 39200 36138 39800 36168
rect 38193 36136 39800 36138
rect 38193 36080 38198 36136
rect 38254 36080 39800 36136
rect 38193 36078 39800 36080
rect 38193 36075 38259 36078
rect 39200 36048 39800 36078
rect 7373 36004 7439 36005
rect 7373 36000 7420 36004
rect 7484 36002 7490 36004
rect 16205 36002 16271 36005
rect 17401 36002 17467 36005
rect 7373 35944 7378 36000
rect 7373 35940 7420 35944
rect 7484 35942 7530 36002
rect 16205 36000 17467 36002
rect 16205 35944 16210 36000
rect 16266 35944 17406 36000
rect 17462 35944 17467 36000
rect 16205 35942 17467 35944
rect 7484 35940 7490 35942
rect 7373 35939 7439 35940
rect 16205 35939 16271 35942
rect 17401 35939 17467 35942
rect 20069 36004 20135 36005
rect 20069 36000 20116 36004
rect 20180 36002 20186 36004
rect 20069 35944 20074 36000
rect 20069 35940 20116 35944
rect 20180 35942 20226 36002
rect 20180 35940 20186 35942
rect 20069 35939 20135 35940
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 11605 35866 11671 35869
rect 19333 35866 19399 35869
rect 11605 35864 19399 35866
rect 11605 35808 11610 35864
rect 11666 35808 19338 35864
rect 19394 35808 19399 35864
rect 11605 35806 19399 35808
rect 11605 35803 11671 35806
rect 19333 35803 19399 35806
rect 12985 35730 13051 35733
rect 25405 35730 25471 35733
rect 12985 35728 25471 35730
rect 12985 35672 12990 35728
rect 13046 35672 25410 35728
rect 25466 35672 25471 35728
rect 12985 35670 25471 35672
rect 12985 35667 13051 35670
rect 25405 35667 25471 35670
rect 8201 35594 8267 35597
rect 11421 35594 11487 35597
rect 8201 35592 11487 35594
rect 8201 35536 8206 35592
rect 8262 35536 11426 35592
rect 11482 35536 11487 35592
rect 8201 35534 11487 35536
rect 8201 35531 8267 35534
rect 11421 35531 11487 35534
rect 14733 35594 14799 35597
rect 21265 35594 21331 35597
rect 14733 35592 21331 35594
rect 14733 35536 14738 35592
rect 14794 35536 21270 35592
rect 21326 35536 21331 35592
rect 14733 35534 21331 35536
rect 14733 35531 14799 35534
rect 21265 35531 21331 35534
rect 200 35458 800 35488
rect 1761 35458 1827 35461
rect 200 35456 1827 35458
rect 200 35400 1766 35456
rect 1822 35400 1827 35456
rect 200 35398 1827 35400
rect 200 35368 800 35398
rect 1761 35395 1827 35398
rect 19701 35458 19767 35461
rect 25313 35458 25379 35461
rect 19701 35456 25379 35458
rect 19701 35400 19706 35456
rect 19762 35400 25318 35456
rect 25374 35400 25379 35456
rect 19701 35398 25379 35400
rect 19701 35395 19767 35398
rect 25313 35395 25379 35398
rect 38193 35458 38259 35461
rect 39200 35458 39800 35488
rect 38193 35456 39800 35458
rect 38193 35400 38198 35456
rect 38254 35400 39800 35456
rect 38193 35398 39800 35400
rect 38193 35395 38259 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 39200 35368 39800 35398
rect 34930 35327 35246 35328
rect 15929 35322 15995 35325
rect 23289 35322 23355 35325
rect 15929 35320 23355 35322
rect 15929 35264 15934 35320
rect 15990 35264 23294 35320
rect 23350 35264 23355 35320
rect 15929 35262 23355 35264
rect 15929 35259 15995 35262
rect 23289 35259 23355 35262
rect 13629 35186 13695 35189
rect 20897 35186 20963 35189
rect 13629 35184 20963 35186
rect 13629 35128 13634 35184
rect 13690 35128 20902 35184
rect 20958 35128 20963 35184
rect 13629 35126 20963 35128
rect 13629 35123 13695 35126
rect 20897 35123 20963 35126
rect 8937 35050 9003 35053
rect 9305 35050 9371 35053
rect 8937 35048 9371 35050
rect 8937 34992 8942 35048
rect 8998 34992 9310 35048
rect 9366 34992 9371 35048
rect 8937 34990 9371 34992
rect 8937 34987 9003 34990
rect 9305 34987 9371 34990
rect 12065 35050 12131 35053
rect 17125 35050 17191 35053
rect 20437 35050 20503 35053
rect 12065 35048 17191 35050
rect 12065 34992 12070 35048
rect 12126 34992 17130 35048
rect 17186 34992 17191 35048
rect 12065 34990 17191 34992
rect 12065 34987 12131 34990
rect 17125 34987 17191 34990
rect 19382 35048 20503 35050
rect 19382 34992 20442 35048
rect 20498 34992 20503 35048
rect 19382 34990 20503 34992
rect 4889 34914 4955 34917
rect 9213 34914 9279 34917
rect 4889 34912 9279 34914
rect 4889 34856 4894 34912
rect 4950 34856 9218 34912
rect 9274 34856 9279 34912
rect 4889 34854 9279 34856
rect 4889 34851 4955 34854
rect 9213 34851 9279 34854
rect 15469 34914 15535 34917
rect 16113 34914 16179 34917
rect 19382 34914 19442 34990
rect 20437 34987 20503 34990
rect 15469 34912 19442 34914
rect 15469 34856 15474 34912
rect 15530 34856 16118 34912
rect 16174 34856 19442 34912
rect 15469 34854 19442 34856
rect 20069 34914 20135 34917
rect 23105 34914 23171 34917
rect 20069 34912 23171 34914
rect 20069 34856 20074 34912
rect 20130 34856 23110 34912
rect 23166 34856 23171 34912
rect 20069 34854 23171 34856
rect 15469 34851 15535 34854
rect 16113 34851 16179 34854
rect 20069 34851 20135 34854
rect 23105 34851 23171 34854
rect 19570 34848 19886 34849
rect 200 34778 800 34808
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 1761 34778 1827 34781
rect 200 34776 1827 34778
rect 200 34720 1766 34776
rect 1822 34720 1827 34776
rect 200 34718 1827 34720
rect 200 34688 800 34718
rect 1761 34715 1827 34718
rect 16021 34778 16087 34781
rect 18045 34778 18111 34781
rect 16021 34776 18111 34778
rect 16021 34720 16026 34776
rect 16082 34720 18050 34776
rect 18106 34720 18111 34776
rect 16021 34718 18111 34720
rect 16021 34715 16087 34718
rect 18045 34715 18111 34718
rect 11605 34642 11671 34645
rect 20713 34642 20779 34645
rect 11605 34640 20779 34642
rect 11605 34584 11610 34640
rect 11666 34584 20718 34640
rect 20774 34584 20779 34640
rect 11605 34582 20779 34584
rect 11605 34579 11671 34582
rect 20713 34579 20779 34582
rect 11053 34506 11119 34509
rect 21265 34506 21331 34509
rect 11053 34504 21331 34506
rect 11053 34448 11058 34504
rect 11114 34448 21270 34504
rect 21326 34448 21331 34504
rect 11053 34446 21331 34448
rect 11053 34443 11119 34446
rect 21265 34443 21331 34446
rect 13353 34370 13419 34373
rect 18505 34370 18571 34373
rect 13353 34368 18571 34370
rect 13353 34312 13358 34368
rect 13414 34312 18510 34368
rect 18566 34312 18571 34368
rect 13353 34310 18571 34312
rect 13353 34307 13419 34310
rect 18505 34307 18571 34310
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 12249 34234 12315 34237
rect 15285 34234 15351 34237
rect 12249 34232 15351 34234
rect 12249 34176 12254 34232
rect 12310 34176 15290 34232
rect 15346 34176 15351 34232
rect 12249 34174 15351 34176
rect 12249 34171 12315 34174
rect 15285 34171 15351 34174
rect 15561 34234 15627 34237
rect 27245 34234 27311 34237
rect 15561 34232 27311 34234
rect 15561 34176 15566 34232
rect 15622 34176 27250 34232
rect 27306 34176 27311 34232
rect 15561 34174 27311 34176
rect 15561 34171 15627 34174
rect 27245 34171 27311 34174
rect 2405 34098 2471 34101
rect 23841 34098 23907 34101
rect 2405 34096 23907 34098
rect 2405 34040 2410 34096
rect 2466 34040 23846 34096
rect 23902 34040 23907 34096
rect 2405 34038 23907 34040
rect 2405 34035 2471 34038
rect 23841 34035 23907 34038
rect 38193 34098 38259 34101
rect 39200 34098 39800 34128
rect 38193 34096 39800 34098
rect 38193 34040 38198 34096
rect 38254 34040 39800 34096
rect 38193 34038 39800 34040
rect 38193 34035 38259 34038
rect 39200 34008 39800 34038
rect 5901 33962 5967 33965
rect 23933 33962 23999 33965
rect 5901 33960 23999 33962
rect 5901 33904 5906 33960
rect 5962 33904 23938 33960
rect 23994 33904 23999 33960
rect 5901 33902 23999 33904
rect 5901 33899 5967 33902
rect 23933 33899 23999 33902
rect 11881 33826 11947 33829
rect 19149 33826 19215 33829
rect 11881 33824 19215 33826
rect 11881 33768 11886 33824
rect 11942 33768 19154 33824
rect 19210 33768 19215 33824
rect 11881 33766 19215 33768
rect 11881 33763 11947 33766
rect 19149 33763 19215 33766
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 12617 33690 12683 33693
rect 17493 33690 17559 33693
rect 12617 33688 17559 33690
rect 12617 33632 12622 33688
rect 12678 33632 17498 33688
rect 17554 33632 17559 33688
rect 12617 33630 17559 33632
rect 12617 33627 12683 33630
rect 17493 33627 17559 33630
rect 4061 33554 4127 33557
rect 18873 33554 18939 33557
rect 4061 33552 18939 33554
rect 4061 33496 4066 33552
rect 4122 33496 18878 33552
rect 18934 33496 18939 33552
rect 4061 33494 18939 33496
rect 4061 33491 4127 33494
rect 18873 33491 18939 33494
rect 19517 33554 19583 33557
rect 22737 33554 22803 33557
rect 19517 33552 22803 33554
rect 19517 33496 19522 33552
rect 19578 33496 22742 33552
rect 22798 33496 22803 33552
rect 19517 33494 22803 33496
rect 19517 33491 19583 33494
rect 22737 33491 22803 33494
rect 200 33418 800 33448
rect 1761 33418 1827 33421
rect 200 33416 1827 33418
rect 200 33360 1766 33416
rect 1822 33360 1827 33416
rect 200 33358 1827 33360
rect 200 33328 800 33358
rect 1761 33355 1827 33358
rect 15837 33418 15903 33421
rect 19701 33418 19767 33421
rect 15837 33416 19767 33418
rect 15837 33360 15842 33416
rect 15898 33360 19706 33416
rect 19762 33360 19767 33416
rect 15837 33358 19767 33360
rect 15837 33355 15903 33358
rect 19701 33355 19767 33358
rect 15561 33282 15627 33285
rect 16205 33282 16271 33285
rect 25773 33282 25839 33285
rect 15561 33280 25839 33282
rect 15561 33224 15566 33280
rect 15622 33224 16210 33280
rect 16266 33224 25778 33280
rect 25834 33224 25839 33280
rect 15561 33222 25839 33224
rect 15561 33219 15627 33222
rect 16205 33219 16271 33222
rect 25773 33219 25839 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 11605 33146 11671 33149
rect 26233 33146 26299 33149
rect 11605 33144 26299 33146
rect 11605 33088 11610 33144
rect 11666 33088 26238 33144
rect 26294 33088 26299 33144
rect 11605 33086 26299 33088
rect 11605 33083 11671 33086
rect 26233 33083 26299 33086
rect 13721 33010 13787 33013
rect 20529 33010 20595 33013
rect 13721 33008 20595 33010
rect 13721 32952 13726 33008
rect 13782 32952 20534 33008
rect 20590 32952 20595 33008
rect 13721 32950 20595 32952
rect 13721 32947 13787 32950
rect 20529 32947 20595 32950
rect 20662 32948 20668 33012
rect 20732 33010 20738 33012
rect 22001 33010 22067 33013
rect 20732 33008 22067 33010
rect 20732 32952 22006 33008
rect 22062 32952 22067 33008
rect 20732 32950 22067 32952
rect 20732 32948 20738 32950
rect 22001 32947 22067 32950
rect 14917 32874 14983 32877
rect 17309 32874 17375 32877
rect 24577 32874 24643 32877
rect 14917 32872 17375 32874
rect 14917 32816 14922 32872
rect 14978 32816 17314 32872
rect 17370 32816 17375 32872
rect 14917 32814 17375 32816
rect 14917 32811 14983 32814
rect 17309 32811 17375 32814
rect 17542 32872 24643 32874
rect 17542 32816 24582 32872
rect 24638 32816 24643 32872
rect 17542 32814 24643 32816
rect 12985 32738 13051 32741
rect 17542 32738 17602 32814
rect 24577 32811 24643 32814
rect 12985 32736 17602 32738
rect 12985 32680 12990 32736
rect 13046 32680 17602 32736
rect 12985 32678 17602 32680
rect 38193 32738 38259 32741
rect 39200 32738 39800 32768
rect 38193 32736 39800 32738
rect 38193 32680 38198 32736
rect 38254 32680 39800 32736
rect 38193 32678 39800 32680
rect 12985 32675 13051 32678
rect 38193 32675 38259 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 39200 32648 39800 32678
rect 19570 32607 19886 32608
rect 11881 32466 11947 32469
rect 28349 32466 28415 32469
rect 11881 32464 28415 32466
rect 11881 32408 11886 32464
rect 11942 32408 28354 32464
rect 28410 32408 28415 32464
rect 11881 32406 28415 32408
rect 11881 32403 11947 32406
rect 28349 32403 28415 32406
rect 14365 32330 14431 32333
rect 15469 32330 15535 32333
rect 20253 32332 20319 32333
rect 20253 32330 20300 32332
rect 14365 32328 15535 32330
rect 14365 32272 14370 32328
rect 14426 32272 15474 32328
rect 15530 32272 15535 32328
rect 14365 32270 15535 32272
rect 20208 32328 20300 32330
rect 20208 32272 20258 32328
rect 20208 32270 20300 32272
rect 14365 32267 14431 32270
rect 15469 32267 15535 32270
rect 20253 32268 20300 32270
rect 20364 32268 20370 32332
rect 20253 32267 20319 32268
rect 19609 32194 19675 32197
rect 21909 32194 21975 32197
rect 19609 32192 21975 32194
rect 19609 32136 19614 32192
rect 19670 32136 21914 32192
rect 21970 32136 21975 32192
rect 19609 32134 21975 32136
rect 19609 32131 19675 32134
rect 21909 32131 21975 32134
rect 4210 32128 4526 32129
rect 200 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1669 32058 1735 32061
rect 200 32056 1735 32058
rect 200 32000 1674 32056
rect 1730 32000 1735 32056
rect 200 31998 1735 32000
rect 200 31968 800 31998
rect 1669 31995 1735 31998
rect 38193 32058 38259 32061
rect 39200 32058 39800 32088
rect 38193 32056 39800 32058
rect 38193 32000 38198 32056
rect 38254 32000 39800 32056
rect 38193 31998 39800 32000
rect 38193 31995 38259 31998
rect 39200 31968 39800 31998
rect 12249 31922 12315 31925
rect 13905 31922 13971 31925
rect 17861 31922 17927 31925
rect 12249 31920 17927 31922
rect 12249 31864 12254 31920
rect 12310 31864 13910 31920
rect 13966 31864 17866 31920
rect 17922 31864 17927 31920
rect 12249 31862 17927 31864
rect 12249 31859 12315 31862
rect 13905 31859 13971 31862
rect 17861 31859 17927 31862
rect 18413 31922 18479 31925
rect 19374 31922 19380 31924
rect 18413 31920 19380 31922
rect 18413 31864 18418 31920
rect 18474 31864 19380 31920
rect 18413 31862 19380 31864
rect 18413 31859 18479 31862
rect 19374 31860 19380 31862
rect 19444 31860 19450 31924
rect 25681 31922 25747 31925
rect 27613 31922 27679 31925
rect 25681 31920 27679 31922
rect 25681 31864 25686 31920
rect 25742 31864 27618 31920
rect 27674 31864 27679 31920
rect 25681 31862 27679 31864
rect 25681 31859 25747 31862
rect 27613 31859 27679 31862
rect 2405 31786 2471 31789
rect 19149 31786 19215 31789
rect 2405 31784 19215 31786
rect 2405 31728 2410 31784
rect 2466 31728 19154 31784
rect 19210 31728 19215 31784
rect 2405 31726 19215 31728
rect 2405 31723 2471 31726
rect 19149 31723 19215 31726
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 200 31378 800 31408
rect 1761 31378 1827 31381
rect 200 31376 1827 31378
rect 200 31320 1766 31376
rect 1822 31320 1827 31376
rect 200 31318 1827 31320
rect 200 31288 800 31318
rect 1761 31315 1827 31318
rect 5349 31378 5415 31381
rect 20897 31378 20963 31381
rect 5349 31376 20963 31378
rect 5349 31320 5354 31376
rect 5410 31320 20902 31376
rect 20958 31320 20963 31376
rect 5349 31318 20963 31320
rect 5349 31315 5415 31318
rect 20897 31315 20963 31318
rect 18781 31244 18847 31245
rect 18781 31242 18828 31244
rect 18736 31240 18828 31242
rect 18736 31184 18786 31240
rect 18736 31182 18828 31184
rect 18781 31180 18828 31182
rect 18892 31180 18898 31244
rect 18781 31179 18847 31180
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 13629 30970 13695 30973
rect 23105 30970 23171 30973
rect 13629 30968 23171 30970
rect 13629 30912 13634 30968
rect 13690 30912 23110 30968
rect 23166 30912 23171 30968
rect 13629 30910 23171 30912
rect 13629 30907 13695 30910
rect 23105 30907 23171 30910
rect 13905 30834 13971 30837
rect 18689 30834 18755 30837
rect 13905 30832 18755 30834
rect 13905 30776 13910 30832
rect 13966 30776 18694 30832
rect 18750 30776 18755 30832
rect 13905 30774 18755 30776
rect 13905 30771 13971 30774
rect 18689 30771 18755 30774
rect 19609 30834 19675 30837
rect 20621 30834 20687 30837
rect 19609 30832 20687 30834
rect 19609 30776 19614 30832
rect 19670 30776 20626 30832
rect 20682 30776 20687 30832
rect 19609 30774 20687 30776
rect 19609 30771 19675 30774
rect 20621 30771 20687 30774
rect 5349 30698 5415 30701
rect 22277 30698 22343 30701
rect 5349 30696 22343 30698
rect 5349 30640 5354 30696
rect 5410 30640 22282 30696
rect 22338 30640 22343 30696
rect 5349 30638 22343 30640
rect 5349 30635 5415 30638
rect 22277 30635 22343 30638
rect 38285 30698 38351 30701
rect 39200 30698 39800 30728
rect 38285 30696 39800 30698
rect 38285 30640 38290 30696
rect 38346 30640 39800 30696
rect 38285 30638 39800 30640
rect 38285 30635 38351 30638
rect 39200 30608 39800 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 15285 30290 15351 30293
rect 17401 30290 17467 30293
rect 15285 30288 17467 30290
rect 15285 30232 15290 30288
rect 15346 30232 17406 30288
rect 17462 30232 17467 30288
rect 15285 30230 17467 30232
rect 15285 30227 15351 30230
rect 17401 30227 17467 30230
rect 200 30018 800 30048
rect 1761 30018 1827 30021
rect 200 30016 1827 30018
rect 200 29960 1766 30016
rect 1822 29960 1827 30016
rect 200 29958 1827 29960
rect 200 29928 800 29958
rect 1761 29955 1827 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 17677 29882 17743 29885
rect 24761 29882 24827 29885
rect 17677 29880 24827 29882
rect 17677 29824 17682 29880
rect 17738 29824 24766 29880
rect 24822 29824 24827 29880
rect 17677 29822 24827 29824
rect 17677 29819 17743 29822
rect 24761 29819 24827 29822
rect 14549 29474 14615 29477
rect 17217 29474 17283 29477
rect 14549 29472 17283 29474
rect 14549 29416 14554 29472
rect 14610 29416 17222 29472
rect 17278 29416 17283 29472
rect 14549 29414 17283 29416
rect 14549 29411 14615 29414
rect 17217 29411 17283 29414
rect 20253 29474 20319 29477
rect 20478 29474 20484 29476
rect 20253 29472 20484 29474
rect 20253 29416 20258 29472
rect 20314 29416 20484 29472
rect 20253 29414 20484 29416
rect 20253 29411 20319 29414
rect 20478 29412 20484 29414
rect 20548 29412 20554 29476
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 19057 29338 19123 29341
rect 12390 29336 19123 29338
rect 12390 29280 19062 29336
rect 19118 29280 19123 29336
rect 12390 29278 19123 29280
rect 4061 29202 4127 29205
rect 12390 29202 12450 29278
rect 19057 29275 19123 29278
rect 19977 29338 20043 29341
rect 20345 29338 20411 29341
rect 19977 29336 20411 29338
rect 19977 29280 19982 29336
rect 20038 29280 20350 29336
rect 20406 29280 20411 29336
rect 19977 29278 20411 29280
rect 19977 29275 20043 29278
rect 20345 29275 20411 29278
rect 37457 29338 37523 29341
rect 39200 29338 39800 29368
rect 37457 29336 39800 29338
rect 37457 29280 37462 29336
rect 37518 29280 39800 29336
rect 37457 29278 39800 29280
rect 37457 29275 37523 29278
rect 39200 29248 39800 29278
rect 22461 29202 22527 29205
rect 4061 29200 12450 29202
rect 4061 29144 4066 29200
rect 4122 29144 12450 29200
rect 4061 29142 12450 29144
rect 17174 29200 22527 29202
rect 17174 29144 22466 29200
rect 22522 29144 22527 29200
rect 17174 29142 22527 29144
rect 4061 29139 4127 29142
rect 1577 29066 1643 29069
rect 1894 29066 1900 29068
rect 1577 29064 1900 29066
rect 1577 29008 1582 29064
rect 1638 29008 1900 29064
rect 1577 29006 1900 29008
rect 1577 29003 1643 29006
rect 1894 29004 1900 29006
rect 1964 29004 1970 29068
rect 12341 29066 12407 29069
rect 17174 29066 17234 29142
rect 22461 29139 22527 29142
rect 24853 29202 24919 29205
rect 26785 29202 26851 29205
rect 24853 29200 26851 29202
rect 24853 29144 24858 29200
rect 24914 29144 26790 29200
rect 26846 29144 26851 29200
rect 24853 29142 26851 29144
rect 24853 29139 24919 29142
rect 26785 29139 26851 29142
rect 12341 29064 17234 29066
rect 12341 29008 12346 29064
rect 12402 29008 17234 29064
rect 12341 29006 17234 29008
rect 18137 29066 18203 29069
rect 18965 29066 19031 29069
rect 18137 29064 19031 29066
rect 18137 29008 18142 29064
rect 18198 29008 18970 29064
rect 19026 29008 19031 29064
rect 18137 29006 19031 29008
rect 12341 29003 12407 29006
rect 18137 29003 18203 29006
rect 18965 29003 19031 29006
rect 19517 29066 19583 29069
rect 22185 29066 22251 29069
rect 19517 29064 22251 29066
rect 19517 29008 19522 29064
rect 19578 29008 22190 29064
rect 22246 29008 22251 29064
rect 19517 29006 22251 29008
rect 19517 29003 19583 29006
rect 22185 29003 22251 29006
rect 14089 28930 14155 28933
rect 21081 28930 21147 28933
rect 14089 28928 21147 28930
rect 14089 28872 14094 28928
rect 14150 28872 21086 28928
rect 21142 28872 21147 28928
rect 14089 28870 21147 28872
rect 14089 28867 14155 28870
rect 21081 28867 21147 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 14733 28794 14799 28797
rect 17309 28794 17375 28797
rect 14733 28792 17375 28794
rect 14733 28736 14738 28792
rect 14794 28736 17314 28792
rect 17370 28736 17375 28792
rect 14733 28734 17375 28736
rect 14733 28731 14799 28734
rect 17309 28731 17375 28734
rect 20069 28794 20135 28797
rect 26417 28794 26483 28797
rect 20069 28792 26483 28794
rect 20069 28736 20074 28792
rect 20130 28736 26422 28792
rect 26478 28736 26483 28792
rect 20069 28734 26483 28736
rect 20069 28731 20135 28734
rect 26417 28731 26483 28734
rect 200 28658 800 28688
rect 1761 28658 1827 28661
rect 200 28656 1827 28658
rect 200 28600 1766 28656
rect 1822 28600 1827 28656
rect 200 28598 1827 28600
rect 200 28568 800 28598
rect 1761 28595 1827 28598
rect 20529 28658 20595 28661
rect 21633 28658 21699 28661
rect 20529 28656 21699 28658
rect 20529 28600 20534 28656
rect 20590 28600 21638 28656
rect 21694 28600 21699 28656
rect 20529 28598 21699 28600
rect 20529 28595 20595 28598
rect 21633 28595 21699 28598
rect 21817 28658 21883 28661
rect 23565 28658 23631 28661
rect 21817 28656 23631 28658
rect 21817 28600 21822 28656
rect 21878 28600 23570 28656
rect 23626 28600 23631 28656
rect 21817 28598 23631 28600
rect 21817 28595 21883 28598
rect 23565 28595 23631 28598
rect 6453 28522 6519 28525
rect 20897 28522 20963 28525
rect 6453 28520 20963 28522
rect 6453 28464 6458 28520
rect 6514 28464 20902 28520
rect 20958 28464 20963 28520
rect 6453 28462 20963 28464
rect 6453 28459 6519 28462
rect 20897 28459 20963 28462
rect 16205 28386 16271 28389
rect 18229 28386 18295 28389
rect 16205 28384 18295 28386
rect 16205 28328 16210 28384
rect 16266 28328 18234 28384
rect 18290 28328 18295 28384
rect 16205 28326 18295 28328
rect 16205 28323 16271 28326
rect 18229 28323 18295 28326
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 21909 28250 21975 28253
rect 24945 28250 25011 28253
rect 21909 28248 25011 28250
rect 21909 28192 21914 28248
rect 21970 28192 24950 28248
rect 25006 28192 25011 28248
rect 21909 28190 25011 28192
rect 21909 28187 21975 28190
rect 24945 28187 25011 28190
rect 38285 27978 38351 27981
rect 39200 27978 39800 28008
rect 38285 27976 39800 27978
rect 38285 27920 38290 27976
rect 38346 27920 39800 27976
rect 38285 27918 39800 27920
rect 38285 27915 38351 27918
rect 39200 27888 39800 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 4981 27708 5047 27709
rect 4981 27704 5028 27708
rect 5092 27706 5098 27708
rect 13629 27706 13695 27709
rect 21449 27706 21515 27709
rect 4981 27648 4986 27704
rect 4981 27644 5028 27648
rect 5092 27646 5138 27706
rect 13629 27704 21515 27706
rect 13629 27648 13634 27704
rect 13690 27648 21454 27704
rect 21510 27648 21515 27704
rect 13629 27646 21515 27648
rect 5092 27644 5098 27646
rect 4981 27643 5047 27644
rect 13629 27643 13695 27646
rect 21449 27643 21515 27646
rect 15009 27570 15075 27573
rect 20897 27570 20963 27573
rect 15009 27568 20963 27570
rect 15009 27512 15014 27568
rect 15070 27512 20902 27568
rect 20958 27512 20963 27568
rect 15009 27510 20963 27512
rect 15009 27507 15075 27510
rect 20897 27507 20963 27510
rect 21909 27570 21975 27573
rect 22185 27570 22251 27573
rect 21909 27568 22251 27570
rect 21909 27512 21914 27568
rect 21970 27512 22190 27568
rect 22246 27512 22251 27568
rect 21909 27510 22251 27512
rect 21909 27507 21975 27510
rect 22185 27507 22251 27510
rect 19793 27434 19859 27437
rect 24301 27434 24367 27437
rect 19793 27432 24367 27434
rect 19793 27376 19798 27432
rect 19854 27376 24306 27432
rect 24362 27376 24367 27432
rect 19793 27374 24367 27376
rect 19793 27371 19859 27374
rect 24301 27371 24367 27374
rect 200 27298 800 27328
rect 1761 27298 1827 27301
rect 200 27296 1827 27298
rect 200 27240 1766 27296
rect 1822 27240 1827 27296
rect 200 27238 1827 27240
rect 200 27208 800 27238
rect 1761 27235 1827 27238
rect 38193 27298 38259 27301
rect 39200 27298 39800 27328
rect 38193 27296 39800 27298
rect 38193 27240 38198 27296
rect 38254 27240 39800 27296
rect 38193 27238 39800 27240
rect 38193 27235 38259 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 39200 27208 39800 27238
rect 19570 27167 19886 27168
rect 19425 27026 19491 27029
rect 26601 27026 26667 27029
rect 19425 27024 26667 27026
rect 19425 26968 19430 27024
rect 19486 26968 26606 27024
rect 26662 26968 26667 27024
rect 19425 26966 26667 26968
rect 19425 26963 19491 26966
rect 26601 26963 26667 26966
rect 19977 26890 20043 26893
rect 20662 26890 20668 26892
rect 19977 26888 20668 26890
rect 19977 26832 19982 26888
rect 20038 26832 20668 26888
rect 19977 26830 20668 26832
rect 19977 26827 20043 26830
rect 20662 26828 20668 26830
rect 20732 26828 20738 26892
rect 4210 26688 4526 26689
rect 200 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 1761 26618 1827 26621
rect 200 26616 1827 26618
rect 200 26560 1766 26616
rect 1822 26560 1827 26616
rect 200 26558 1827 26560
rect 200 26528 800 26558
rect 1761 26555 1827 26558
rect 17217 26482 17283 26485
rect 23105 26482 23171 26485
rect 17217 26480 23171 26482
rect 17217 26424 17222 26480
rect 17278 26424 23110 26480
rect 23166 26424 23171 26480
rect 17217 26422 23171 26424
rect 17217 26419 17283 26422
rect 23105 26419 23171 26422
rect 1577 26346 1643 26349
rect 2262 26346 2268 26348
rect 1577 26344 2268 26346
rect 1577 26288 1582 26344
rect 1638 26288 2268 26344
rect 1577 26286 2268 26288
rect 1577 26283 1643 26286
rect 2262 26284 2268 26286
rect 2332 26284 2338 26348
rect 5073 26346 5139 26349
rect 5206 26346 5212 26348
rect 5073 26344 5212 26346
rect 5073 26288 5078 26344
rect 5134 26288 5212 26344
rect 5073 26286 5212 26288
rect 5073 26283 5139 26286
rect 5206 26284 5212 26286
rect 5276 26284 5282 26348
rect 7005 26346 7071 26349
rect 15009 26346 15075 26349
rect 7005 26344 15075 26346
rect 7005 26288 7010 26344
rect 7066 26288 15014 26344
rect 15070 26288 15075 26344
rect 7005 26286 15075 26288
rect 7005 26283 7071 26286
rect 15009 26283 15075 26286
rect 17769 26346 17835 26349
rect 17902 26346 17908 26348
rect 17769 26344 17908 26346
rect 17769 26288 17774 26344
rect 17830 26288 17908 26344
rect 17769 26286 17908 26288
rect 17769 26283 17835 26286
rect 17902 26284 17908 26286
rect 17972 26284 17978 26348
rect 18965 26346 19031 26349
rect 21081 26346 21147 26349
rect 18965 26344 21147 26346
rect 18965 26288 18970 26344
rect 19026 26288 21086 26344
rect 21142 26288 21147 26344
rect 18965 26286 21147 26288
rect 18965 26283 19031 26286
rect 21081 26283 21147 26286
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 17401 25938 17467 25941
rect 21633 25938 21699 25941
rect 17401 25936 21699 25938
rect 17401 25880 17406 25936
rect 17462 25880 21638 25936
rect 21694 25880 21699 25936
rect 17401 25878 21699 25880
rect 17401 25875 17467 25878
rect 21633 25875 21699 25878
rect 38285 25938 38351 25941
rect 39200 25938 39800 25968
rect 38285 25936 39800 25938
rect 38285 25880 38290 25936
rect 38346 25880 39800 25936
rect 38285 25878 39800 25880
rect 38285 25875 38351 25878
rect 39200 25848 39800 25878
rect 11421 25802 11487 25805
rect 19149 25802 19215 25805
rect 11421 25800 19215 25802
rect 11421 25744 11426 25800
rect 11482 25744 19154 25800
rect 19210 25744 19215 25800
rect 11421 25742 19215 25744
rect 11421 25739 11487 25742
rect 19149 25739 19215 25742
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 200 25258 800 25288
rect 1669 25258 1735 25261
rect 200 25256 1735 25258
rect 200 25200 1674 25256
rect 1730 25200 1735 25256
rect 200 25198 1735 25200
rect 200 25168 800 25198
rect 1669 25195 1735 25198
rect 8661 25122 8727 25125
rect 9806 25122 9812 25124
rect 8661 25120 9812 25122
rect 8661 25064 8666 25120
rect 8722 25064 9812 25120
rect 8661 25062 9812 25064
rect 8661 25059 8727 25062
rect 9806 25060 9812 25062
rect 9876 25060 9882 25124
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 20621 24988 20687 24989
rect 20621 24986 20668 24988
rect 20576 24984 20668 24986
rect 20576 24928 20626 24984
rect 20576 24926 20668 24928
rect 20621 24924 20668 24926
rect 20732 24924 20738 24988
rect 20621 24923 20687 24924
rect 19977 24850 20043 24853
rect 21541 24850 21607 24853
rect 19977 24848 21607 24850
rect 19977 24792 19982 24848
rect 20038 24792 21546 24848
rect 21602 24792 21607 24848
rect 19977 24790 21607 24792
rect 19977 24787 20043 24790
rect 21541 24787 21607 24790
rect 15469 24714 15535 24717
rect 17401 24714 17467 24717
rect 15469 24712 17467 24714
rect 15469 24656 15474 24712
rect 15530 24656 17406 24712
rect 17462 24656 17467 24712
rect 15469 24654 17467 24656
rect 15469 24651 15535 24654
rect 17401 24651 17467 24654
rect 21725 24714 21791 24717
rect 24025 24714 24091 24717
rect 21725 24712 24091 24714
rect 21725 24656 21730 24712
rect 21786 24656 24030 24712
rect 24086 24656 24091 24712
rect 21725 24654 24091 24656
rect 21725 24651 21791 24654
rect 24025 24651 24091 24654
rect 17125 24578 17191 24581
rect 18045 24578 18111 24581
rect 20989 24578 21055 24581
rect 17125 24576 21055 24578
rect 17125 24520 17130 24576
rect 17186 24520 18050 24576
rect 18106 24520 20994 24576
rect 21050 24520 21055 24576
rect 17125 24518 21055 24520
rect 17125 24515 17191 24518
rect 18045 24515 18111 24518
rect 20989 24515 21055 24518
rect 38193 24578 38259 24581
rect 39200 24578 39800 24608
rect 38193 24576 39800 24578
rect 38193 24520 38198 24576
rect 38254 24520 39800 24576
rect 38193 24518 39800 24520
rect 38193 24515 38259 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 39200 24488 39800 24518
rect 34930 24447 35246 24448
rect 21725 24170 21791 24173
rect 21909 24170 21975 24173
rect 21725 24168 21975 24170
rect 21725 24112 21730 24168
rect 21786 24112 21914 24168
rect 21970 24112 21975 24168
rect 21725 24110 21975 24112
rect 21725 24107 21791 24110
rect 21909 24107 21975 24110
rect 19570 23968 19886 23969
rect 200 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 1761 23898 1827 23901
rect 200 23896 1827 23898
rect 200 23840 1766 23896
rect 1822 23840 1827 23896
rect 200 23838 1827 23840
rect 200 23808 800 23838
rect 1761 23835 1827 23838
rect 38193 23898 38259 23901
rect 39200 23898 39800 23928
rect 38193 23896 39800 23898
rect 38193 23840 38198 23896
rect 38254 23840 39800 23896
rect 38193 23838 39800 23840
rect 38193 23835 38259 23838
rect 39200 23808 39800 23838
rect 4521 23626 4587 23629
rect 4838 23626 4844 23628
rect 4521 23624 4844 23626
rect 4521 23568 4526 23624
rect 4582 23568 4844 23624
rect 4521 23566 4844 23568
rect 4521 23563 4587 23566
rect 4838 23564 4844 23566
rect 4908 23564 4914 23628
rect 16849 23626 16915 23629
rect 21817 23626 21883 23629
rect 22553 23626 22619 23629
rect 16849 23624 22619 23626
rect 16849 23568 16854 23624
rect 16910 23568 21822 23624
rect 21878 23568 22558 23624
rect 22614 23568 22619 23624
rect 16849 23566 22619 23568
rect 16849 23563 16915 23566
rect 21817 23563 21883 23566
rect 22553 23563 22619 23566
rect 22001 23490 22067 23493
rect 22277 23490 22343 23493
rect 22001 23488 22343 23490
rect 22001 23432 22006 23488
rect 22062 23432 22282 23488
rect 22338 23432 22343 23488
rect 22001 23430 22343 23432
rect 22001 23427 22067 23430
rect 22277 23427 22343 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 200 23218 800 23248
rect 2773 23218 2839 23221
rect 200 23216 2839 23218
rect 200 23160 2778 23216
rect 2834 23160 2839 23216
rect 200 23158 2839 23160
rect 200 23128 800 23158
rect 2773 23155 2839 23158
rect 12801 23082 12867 23085
rect 17401 23082 17467 23085
rect 12801 23080 17467 23082
rect 12801 23024 12806 23080
rect 12862 23024 17406 23080
rect 17462 23024 17467 23080
rect 12801 23022 17467 23024
rect 12801 23019 12867 23022
rect 17401 23019 17467 23022
rect 11053 22946 11119 22949
rect 11053 22944 12450 22946
rect 11053 22888 11058 22944
rect 11114 22888 12450 22944
rect 11053 22886 12450 22888
rect 11053 22883 11119 22886
rect 12390 22674 12450 22886
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 30925 22674 30991 22677
rect 12390 22672 30991 22674
rect 12390 22616 30930 22672
rect 30986 22616 30991 22672
rect 12390 22614 30991 22616
rect 30925 22611 30991 22614
rect 17769 22538 17835 22541
rect 17902 22538 17908 22540
rect 17769 22536 17908 22538
rect 17769 22480 17774 22536
rect 17830 22480 17908 22536
rect 17769 22478 17908 22480
rect 17769 22475 17835 22478
rect 17902 22476 17908 22478
rect 17972 22476 17978 22540
rect 38193 22538 38259 22541
rect 39200 22538 39800 22568
rect 38193 22536 39800 22538
rect 38193 22480 38198 22536
rect 38254 22480 39800 22536
rect 38193 22478 39800 22480
rect 38193 22475 38259 22478
rect 39200 22448 39800 22478
rect 5758 22340 5764 22404
rect 5828 22402 5834 22404
rect 5993 22402 6059 22405
rect 5828 22400 6059 22402
rect 5828 22344 5998 22400
rect 6054 22344 6059 22400
rect 5828 22342 6059 22344
rect 5828 22340 5834 22342
rect 5993 22339 6059 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 20529 22266 20595 22269
rect 20662 22266 20668 22268
rect 20529 22264 20668 22266
rect 20529 22208 20534 22264
rect 20590 22208 20668 22264
rect 20529 22206 20668 22208
rect 20529 22203 20595 22206
rect 20662 22204 20668 22206
rect 20732 22204 20738 22268
rect 5349 22132 5415 22133
rect 5349 22130 5396 22132
rect 5304 22128 5396 22130
rect 5304 22072 5354 22128
rect 5304 22070 5396 22072
rect 5349 22068 5396 22070
rect 5460 22068 5466 22132
rect 19149 22130 19215 22133
rect 21633 22130 21699 22133
rect 19149 22128 21699 22130
rect 19149 22072 19154 22128
rect 19210 22072 21638 22128
rect 21694 22072 21699 22128
rect 19149 22070 21699 22072
rect 5349 22067 5415 22068
rect 19149 22067 19215 22070
rect 21633 22067 21699 22070
rect 200 21858 800 21888
rect 1669 21858 1735 21861
rect 200 21856 1735 21858
rect 200 21800 1674 21856
rect 1730 21800 1735 21856
rect 200 21798 1735 21800
rect 200 21768 800 21798
rect 1669 21795 1735 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 38193 21178 38259 21181
rect 39200 21178 39800 21208
rect 38193 21176 39800 21178
rect 38193 21120 38198 21176
rect 38254 21120 39800 21176
rect 38193 21118 39800 21120
rect 38193 21115 38259 21118
rect 39200 21088 39800 21118
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 200 20498 800 20528
rect 1669 20498 1735 20501
rect 200 20496 1735 20498
rect 200 20440 1674 20496
rect 1730 20440 1735 20496
rect 200 20438 1735 20440
rect 200 20408 800 20438
rect 1669 20435 1735 20438
rect 19977 20498 20043 20501
rect 20478 20498 20484 20500
rect 19977 20496 20484 20498
rect 19977 20440 19982 20496
rect 20038 20440 20484 20496
rect 19977 20438 20484 20440
rect 19977 20435 20043 20438
rect 20478 20436 20484 20438
rect 20548 20436 20554 20500
rect 37181 20498 37247 20501
rect 39200 20498 39800 20528
rect 37181 20496 39800 20498
rect 37181 20440 37186 20496
rect 37242 20440 39800 20496
rect 37181 20438 39800 20440
rect 37181 20435 37247 20438
rect 39200 20408 39800 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 18822 19756 18828 19820
rect 18892 19818 18898 19820
rect 22093 19818 22159 19821
rect 18892 19816 22159 19818
rect 18892 19760 22098 19816
rect 22154 19760 22159 19816
rect 18892 19758 22159 19760
rect 18892 19756 18898 19758
rect 22093 19755 22159 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 3182 19348 3188 19412
rect 3252 19410 3258 19412
rect 3417 19410 3483 19413
rect 3252 19408 3483 19410
rect 3252 19352 3422 19408
rect 3478 19352 3483 19408
rect 3252 19350 3483 19352
rect 3252 19348 3258 19350
rect 3417 19347 3483 19350
rect 17902 19212 17908 19276
rect 17972 19274 17978 19276
rect 23565 19274 23631 19277
rect 17972 19272 23631 19274
rect 17972 19216 23570 19272
rect 23626 19216 23631 19272
rect 17972 19214 23631 19216
rect 17972 19212 17978 19214
rect 23565 19211 23631 19214
rect 200 19138 800 19168
rect 1761 19138 1827 19141
rect 200 19136 1827 19138
rect 200 19080 1766 19136
rect 1822 19080 1827 19136
rect 200 19078 1827 19080
rect 200 19048 800 19078
rect 1761 19075 1827 19078
rect 38285 19138 38351 19141
rect 39200 19138 39800 19168
rect 38285 19136 39800 19138
rect 38285 19080 38290 19136
rect 38346 19080 39800 19136
rect 38285 19078 39800 19080
rect 38285 19075 38351 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 39800 19078
rect 34930 19007 35246 19008
rect 5165 18866 5231 18869
rect 5574 18866 5580 18868
rect 5165 18864 5580 18866
rect 5165 18808 5170 18864
rect 5226 18808 5580 18864
rect 5165 18806 5580 18808
rect 5165 18803 5231 18806
rect 5574 18804 5580 18806
rect 5644 18804 5650 18868
rect 19570 18528 19886 18529
rect 200 18458 800 18488
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 1669 18458 1735 18461
rect 200 18456 1735 18458
rect 200 18400 1674 18456
rect 1730 18400 1735 18456
rect 200 18398 1735 18400
rect 200 18368 800 18398
rect 1669 18395 1735 18398
rect 15009 18322 15075 18325
rect 17769 18322 17835 18325
rect 15009 18320 17835 18322
rect 15009 18264 15014 18320
rect 15070 18264 17774 18320
rect 17830 18264 17835 18320
rect 15009 18262 17835 18264
rect 15009 18259 15075 18262
rect 17769 18259 17835 18262
rect 19885 18322 19951 18325
rect 28349 18322 28415 18325
rect 19885 18320 28415 18322
rect 19885 18264 19890 18320
rect 19946 18264 28354 18320
rect 28410 18264 28415 18320
rect 19885 18262 28415 18264
rect 19885 18259 19951 18262
rect 28349 18259 28415 18262
rect 3509 18186 3575 18189
rect 7414 18186 7420 18188
rect 3509 18184 7420 18186
rect 3509 18128 3514 18184
rect 3570 18128 7420 18184
rect 3509 18126 7420 18128
rect 3509 18123 3575 18126
rect 7414 18124 7420 18126
rect 7484 18186 7490 18188
rect 7833 18186 7899 18189
rect 7484 18184 7899 18186
rect 7484 18128 7838 18184
rect 7894 18128 7899 18184
rect 7484 18126 7899 18128
rect 7484 18124 7490 18126
rect 7833 18123 7899 18126
rect 19885 18186 19951 18189
rect 22921 18186 22987 18189
rect 19885 18184 22987 18186
rect 19885 18128 19890 18184
rect 19946 18128 22926 18184
rect 22982 18128 22987 18184
rect 19885 18126 22987 18128
rect 19885 18123 19951 18126
rect 22921 18123 22987 18126
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 7649 17914 7715 17917
rect 8150 17914 8156 17916
rect 7649 17912 8156 17914
rect 7649 17856 7654 17912
rect 7710 17856 8156 17912
rect 7649 17854 8156 17856
rect 7649 17851 7715 17854
rect 8150 17852 8156 17854
rect 8220 17852 8226 17916
rect 3601 17778 3667 17781
rect 6862 17778 6868 17780
rect 3601 17776 6868 17778
rect 3601 17720 3606 17776
rect 3662 17720 6868 17776
rect 3601 17718 6868 17720
rect 3601 17715 3667 17718
rect 6862 17716 6868 17718
rect 6932 17716 6938 17780
rect 19885 17778 19951 17781
rect 24577 17778 24643 17781
rect 19885 17776 24643 17778
rect 19885 17720 19890 17776
rect 19946 17720 24582 17776
rect 24638 17720 24643 17776
rect 19885 17718 24643 17720
rect 19885 17715 19951 17718
rect 24577 17715 24643 17718
rect 38193 17778 38259 17781
rect 39200 17778 39800 17808
rect 38193 17776 39800 17778
rect 38193 17720 38198 17776
rect 38254 17720 39800 17776
rect 38193 17718 39800 17720
rect 38193 17715 38259 17718
rect 39200 17688 39800 17718
rect 19609 17642 19675 17645
rect 21173 17642 21239 17645
rect 19609 17640 21239 17642
rect 19609 17584 19614 17640
rect 19670 17584 21178 17640
rect 21234 17584 21239 17640
rect 19609 17582 21239 17584
rect 19609 17579 19675 17582
rect 21173 17579 21239 17582
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 14181 17234 14247 17237
rect 17217 17234 17283 17237
rect 14181 17232 17283 17234
rect 14181 17176 14186 17232
rect 14242 17176 17222 17232
rect 17278 17176 17283 17232
rect 14181 17174 17283 17176
rect 14181 17171 14247 17174
rect 17217 17171 17283 17174
rect 200 17098 800 17128
rect 1669 17098 1735 17101
rect 200 17096 1735 17098
rect 200 17040 1674 17096
rect 1730 17040 1735 17096
rect 200 17038 1735 17040
rect 200 17008 800 17038
rect 1669 17035 1735 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 38193 16418 38259 16421
rect 39200 16418 39800 16448
rect 38193 16416 39800 16418
rect 38193 16360 38198 16416
rect 38254 16360 39800 16416
rect 38193 16358 39800 16360
rect 38193 16355 38259 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 39200 16328 39800 16358
rect 19570 16287 19886 16288
rect 4705 16146 4771 16149
rect 5533 16146 5599 16149
rect 4705 16144 5599 16146
rect 4705 16088 4710 16144
rect 4766 16088 5538 16144
rect 5594 16088 5599 16144
rect 4705 16086 5599 16088
rect 4705 16083 4771 16086
rect 5533 16083 5599 16086
rect 13077 16146 13143 16149
rect 18965 16146 19031 16149
rect 13077 16144 19031 16146
rect 13077 16088 13082 16144
rect 13138 16088 18970 16144
rect 19026 16088 19031 16144
rect 13077 16086 19031 16088
rect 13077 16083 13143 16086
rect 18965 16083 19031 16086
rect 2221 16010 2287 16013
rect 10409 16010 10475 16013
rect 2221 16008 10475 16010
rect 2221 15952 2226 16008
rect 2282 15952 10414 16008
rect 10470 15952 10475 16008
rect 2221 15950 10475 15952
rect 2221 15947 2287 15950
rect 10409 15947 10475 15950
rect 5257 15874 5323 15877
rect 9305 15874 9371 15877
rect 5257 15872 9371 15874
rect 5257 15816 5262 15872
rect 5318 15816 9310 15872
rect 9366 15816 9371 15872
rect 5257 15814 9371 15816
rect 5257 15811 5323 15814
rect 9305 15811 9371 15814
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1761 15738 1827 15741
rect 200 15736 1827 15738
rect 200 15680 1766 15736
rect 1822 15680 1827 15736
rect 200 15678 1827 15680
rect 200 15648 800 15678
rect 1761 15675 1827 15678
rect 38193 15738 38259 15741
rect 39200 15738 39800 15768
rect 38193 15736 39800 15738
rect 38193 15680 38198 15736
rect 38254 15680 39800 15736
rect 38193 15678 39800 15680
rect 38193 15675 38259 15678
rect 39200 15648 39800 15678
rect 5441 15466 5507 15469
rect 6913 15466 6979 15469
rect 5441 15464 6979 15466
rect 5441 15408 5446 15464
rect 5502 15408 6918 15464
rect 6974 15408 6979 15464
rect 5441 15406 6979 15408
rect 5441 15403 5507 15406
rect 6913 15403 6979 15406
rect 15469 15466 15535 15469
rect 17033 15466 17099 15469
rect 15469 15464 17099 15466
rect 15469 15408 15474 15464
rect 15530 15408 17038 15464
rect 17094 15408 17099 15464
rect 15469 15406 17099 15408
rect 15469 15403 15535 15406
rect 17033 15403 17099 15406
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 9765 15196 9831 15197
rect 9765 15192 9812 15196
rect 9876 15194 9882 15196
rect 9765 15136 9770 15192
rect 9765 15132 9812 15136
rect 9876 15134 9922 15194
rect 9876 15132 9882 15134
rect 9765 15131 9831 15132
rect 200 15058 800 15088
rect 2497 15058 2563 15061
rect 200 15056 2563 15058
rect 200 15000 2502 15056
rect 2558 15000 2563 15056
rect 200 14998 2563 15000
rect 200 14968 800 14998
rect 2497 14995 2563 14998
rect 2865 15058 2931 15061
rect 4889 15058 4955 15061
rect 2865 15056 4955 15058
rect 2865 15000 2870 15056
rect 2926 15000 4894 15056
rect 4950 15000 4955 15056
rect 2865 14998 4955 15000
rect 2865 14995 2931 14998
rect 4889 14995 4955 14998
rect 11697 14786 11763 14789
rect 12065 14786 12131 14789
rect 11697 14784 12131 14786
rect 11697 14728 11702 14784
rect 11758 14728 12070 14784
rect 12126 14728 12131 14784
rect 11697 14726 12131 14728
rect 11697 14723 11763 14726
rect 12065 14723 12131 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19241 14514 19307 14517
rect 21357 14514 21423 14517
rect 19241 14512 21423 14514
rect 19241 14456 19246 14512
rect 19302 14456 21362 14512
rect 21418 14456 21423 14512
rect 19241 14454 21423 14456
rect 19241 14451 19307 14454
rect 21357 14451 21423 14454
rect 2773 14378 2839 14381
rect 13629 14378 13695 14381
rect 2773 14376 13695 14378
rect 2773 14320 2778 14376
rect 2834 14320 13634 14376
rect 13690 14320 13695 14376
rect 2773 14318 13695 14320
rect 2773 14315 2839 14318
rect 13629 14315 13695 14318
rect 22737 14378 22803 14381
rect 25589 14378 25655 14381
rect 22737 14376 25655 14378
rect 22737 14320 22742 14376
rect 22798 14320 25594 14376
rect 25650 14320 25655 14376
rect 22737 14318 25655 14320
rect 22737 14315 22803 14318
rect 25589 14315 25655 14318
rect 38193 14378 38259 14381
rect 39200 14378 39800 14408
rect 38193 14376 39800 14378
rect 38193 14320 38198 14376
rect 38254 14320 39800 14376
rect 38193 14318 39800 14320
rect 38193 14315 38259 14318
rect 39200 14288 39800 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 2681 13834 2747 13837
rect 2814 13834 2820 13836
rect 2681 13832 2820 13834
rect 2681 13776 2686 13832
rect 2742 13776 2820 13832
rect 2681 13774 2820 13776
rect 2681 13771 2747 13774
rect 2814 13772 2820 13774
rect 2884 13772 2890 13836
rect 9765 13834 9831 13837
rect 11237 13834 11303 13837
rect 15193 13834 15259 13837
rect 9765 13832 15259 13834
rect 9765 13776 9770 13832
rect 9826 13776 11242 13832
rect 11298 13776 15198 13832
rect 15254 13776 15259 13832
rect 9765 13774 15259 13776
rect 9765 13771 9831 13774
rect 11237 13771 11303 13774
rect 15193 13771 15259 13774
rect 200 13698 800 13728
rect 1669 13698 1735 13701
rect 5441 13700 5507 13701
rect 5390 13698 5396 13700
rect 200 13696 1735 13698
rect 200 13640 1674 13696
rect 1730 13640 1735 13696
rect 200 13638 1735 13640
rect 5350 13638 5396 13698
rect 5460 13696 5507 13700
rect 5502 13640 5507 13696
rect 200 13608 800 13638
rect 1669 13635 1735 13638
rect 5390 13636 5396 13638
rect 5460 13636 5507 13640
rect 6862 13636 6868 13700
rect 6932 13698 6938 13700
rect 8109 13698 8175 13701
rect 6932 13696 8175 13698
rect 6932 13640 8114 13696
rect 8170 13640 8175 13696
rect 6932 13638 8175 13640
rect 6932 13636 6938 13638
rect 5441 13635 5507 13636
rect 8109 13635 8175 13638
rect 9489 13698 9555 13701
rect 12014 13698 12020 13700
rect 9489 13696 12020 13698
rect 9489 13640 9494 13696
rect 9550 13640 12020 13696
rect 9489 13638 12020 13640
rect 9489 13635 9555 13638
rect 12014 13636 12020 13638
rect 12084 13636 12090 13700
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 38193 13018 38259 13021
rect 39200 13018 39800 13048
rect 38193 13016 39800 13018
rect 38193 12960 38198 13016
rect 38254 12960 39800 13016
rect 38193 12958 39800 12960
rect 38193 12955 38259 12958
rect 39200 12928 39800 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 200 12338 800 12368
rect 1761 12338 1827 12341
rect 200 12336 1827 12338
rect 200 12280 1766 12336
rect 1822 12280 1827 12336
rect 200 12278 1827 12280
rect 200 12248 800 12278
rect 1761 12275 1827 12278
rect 5533 12340 5599 12341
rect 5533 12336 5580 12340
rect 5644 12338 5650 12340
rect 38285 12338 38351 12341
rect 39200 12338 39800 12368
rect 5533 12280 5538 12336
rect 5533 12276 5580 12280
rect 5644 12278 5690 12338
rect 38285 12336 39800 12338
rect 38285 12280 38290 12336
rect 38346 12280 39800 12336
rect 38285 12278 39800 12280
rect 5644 12276 5650 12278
rect 5533 12275 5599 12276
rect 38285 12275 38351 12278
rect 39200 12248 39800 12278
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 2313 11930 2379 11933
rect 5022 11930 5028 11932
rect 2313 11928 5028 11930
rect 2313 11872 2318 11928
rect 2374 11872 5028 11928
rect 2313 11870 5028 11872
rect 2313 11867 2379 11870
rect 5022 11868 5028 11870
rect 5092 11868 5098 11932
rect 8201 11796 8267 11797
rect 8150 11794 8156 11796
rect 8110 11734 8156 11794
rect 8220 11792 8267 11796
rect 8262 11736 8267 11792
rect 8150 11732 8156 11734
rect 8220 11732 8267 11736
rect 8201 11731 8267 11732
rect 200 11658 800 11688
rect 3601 11658 3667 11661
rect 200 11656 3667 11658
rect 200 11600 3606 11656
rect 3662 11600 3667 11656
rect 200 11598 3667 11600
rect 200 11568 800 11598
rect 3601 11595 3667 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 5625 10978 5691 10981
rect 5758 10978 5764 10980
rect 5625 10976 5764 10978
rect 5625 10920 5630 10976
rect 5686 10920 5764 10976
rect 5625 10918 5764 10920
rect 5625 10915 5691 10918
rect 5758 10916 5764 10918
rect 5828 10916 5834 10980
rect 38285 10978 38351 10981
rect 39200 10978 39800 11008
rect 38285 10976 39800 10978
rect 38285 10920 38290 10976
rect 38346 10920 39800 10976
rect 38285 10918 39800 10920
rect 38285 10915 38351 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 39200 10888 39800 10918
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 200 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 3417 10298 3483 10301
rect 200 10296 3483 10298
rect 200 10240 3422 10296
rect 3478 10240 3483 10296
rect 200 10238 3483 10240
rect 200 10208 800 10238
rect 3417 10235 3483 10238
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 3049 9618 3115 9621
rect 3182 9618 3188 9620
rect 3049 9616 3188 9618
rect 3049 9560 3054 9616
rect 3110 9560 3188 9616
rect 3049 9558 3188 9560
rect 3049 9555 3115 9558
rect 3182 9556 3188 9558
rect 3252 9556 3258 9620
rect 3601 9618 3667 9621
rect 5206 9618 5212 9620
rect 3601 9616 5212 9618
rect 3601 9560 3606 9616
rect 3662 9560 5212 9616
rect 3601 9558 5212 9560
rect 3601 9555 3667 9558
rect 5206 9556 5212 9558
rect 5276 9556 5282 9620
rect 19425 9618 19491 9621
rect 20161 9618 20227 9621
rect 20294 9618 20300 9620
rect 19425 9616 20300 9618
rect 19425 9560 19430 9616
rect 19486 9560 20166 9616
rect 20222 9560 20300 9616
rect 19425 9558 20300 9560
rect 19425 9555 19491 9558
rect 20161 9555 20227 9558
rect 20294 9556 20300 9558
rect 20364 9556 20370 9620
rect 37181 9618 37247 9621
rect 39200 9618 39800 9648
rect 37181 9616 39800 9618
rect 37181 9560 37186 9616
rect 37242 9560 39800 9616
rect 37181 9558 39800 9560
rect 37181 9555 37247 9558
rect 39200 9528 39800 9558
rect 2814 9420 2820 9484
rect 2884 9482 2890 9484
rect 3141 9482 3207 9485
rect 2884 9480 3207 9482
rect 2884 9424 3146 9480
rect 3202 9424 3207 9480
rect 2884 9422 3207 9424
rect 2884 9420 2890 9422
rect 3141 9419 3207 9422
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 2037 9212 2103 9213
rect 2037 9210 2084 9212
rect 1992 9208 2084 9210
rect 1992 9152 2042 9208
rect 1992 9150 2084 9152
rect 2037 9148 2084 9150
rect 2148 9148 2154 9212
rect 2037 9147 2103 9148
rect 200 8938 800 8968
rect 1761 8938 1827 8941
rect 200 8936 1827 8938
rect 200 8880 1766 8936
rect 1822 8880 1827 8936
rect 200 8878 1827 8880
rect 200 8848 800 8878
rect 1761 8875 1827 8878
rect 15929 8938 15995 8941
rect 20110 8938 20116 8940
rect 15929 8936 20116 8938
rect 15929 8880 15934 8936
rect 15990 8880 20116 8936
rect 15929 8878 20116 8880
rect 15929 8875 15995 8878
rect 20110 8876 20116 8878
rect 20180 8876 20186 8940
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 38285 8258 38351 8261
rect 39200 8258 39800 8288
rect 38285 8256 39800 8258
rect 38285 8200 38290 8256
rect 38346 8200 39800 8256
rect 38285 8198 39800 8200
rect 38285 8195 38351 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 39200 8168 39800 8198
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 200 7578 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 1761 7578 1827 7581
rect 200 7576 1827 7578
rect 200 7520 1766 7576
rect 1822 7520 1827 7576
rect 200 7518 1827 7520
rect 200 7488 800 7518
rect 1761 7515 1827 7518
rect 38285 7578 38351 7581
rect 39200 7578 39800 7608
rect 38285 7576 39800 7578
rect 38285 7520 38290 7576
rect 38346 7520 39800 7576
rect 38285 7518 39800 7520
rect 38285 7515 38351 7518
rect 39200 7488 39800 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 200 6898 800 6928
rect 1761 6898 1827 6901
rect 200 6896 1827 6898
rect 200 6840 1766 6896
rect 1822 6840 1827 6896
rect 200 6838 1827 6840
rect 200 6808 800 6838
rect 1761 6835 1827 6838
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 1945 6492 2011 6493
rect 1894 6490 1900 6492
rect 1854 6430 1900 6490
rect 1964 6488 2011 6492
rect 2006 6432 2011 6488
rect 1894 6428 1900 6430
rect 1964 6428 2011 6432
rect 1945 6427 2011 6428
rect 38285 6218 38351 6221
rect 39200 6218 39800 6248
rect 38285 6216 39800 6218
rect 38285 6160 38290 6216
rect 38346 6160 39800 6216
rect 38285 6158 39800 6160
rect 38285 6155 38351 6158
rect 39200 6128 39800 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 2037 5946 2103 5949
rect 2262 5946 2268 5948
rect 2037 5944 2268 5946
rect 2037 5888 2042 5944
rect 2098 5888 2268 5944
rect 2037 5886 2268 5888
rect 2037 5883 2103 5886
rect 2262 5884 2268 5886
rect 2332 5884 2338 5948
rect 200 5538 800 5568
rect 1761 5538 1827 5541
rect 200 5536 1827 5538
rect 200 5480 1766 5536
rect 1822 5480 1827 5536
rect 200 5478 1827 5480
rect 200 5448 800 5478
rect 1761 5475 1827 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 38193 4858 38259 4861
rect 39200 4858 39800 4888
rect 38193 4856 39800 4858
rect 38193 4800 38198 4856
rect 38254 4800 39800 4856
rect 38193 4798 39800 4800
rect 38193 4795 38259 4798
rect 39200 4768 39800 4798
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 200 4178 800 4208
rect 1761 4178 1827 4181
rect 200 4176 1827 4178
rect 200 4120 1766 4176
rect 1822 4120 1827 4176
rect 200 4118 1827 4120
rect 200 4088 800 4118
rect 1761 4115 1827 4118
rect 38285 4178 38351 4181
rect 39200 4178 39800 4208
rect 38285 4176 39800 4178
rect 38285 4120 38290 4176
rect 38346 4120 39800 4176
rect 38285 4118 39800 4120
rect 38285 4115 38351 4118
rect 39200 4088 39800 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 200 3498 800 3528
rect 1393 3498 1459 3501
rect 200 3496 1459 3498
rect 200 3440 1398 3496
rect 1454 3440 1459 3496
rect 200 3438 1459 3440
rect 200 3408 800 3438
rect 1393 3435 1459 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 3141 3226 3207 3229
rect 4838 3226 4844 3228
rect 3141 3224 4844 3226
rect 3141 3168 3146 3224
rect 3202 3168 4844 3224
rect 3141 3166 4844 3168
rect 3141 3163 3207 3166
rect 4838 3164 4844 3166
rect 4908 3164 4914 3228
rect 38193 2818 38259 2821
rect 39200 2818 39800 2848
rect 38193 2816 39800 2818
rect 38193 2760 38198 2816
rect 38254 2760 39800 2816
rect 38193 2758 39800 2760
rect 38193 2755 38259 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 39200 2728 39800 2758
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 200 2138 800 2168
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 1669 2138 1735 2141
rect 200 2136 1735 2138
rect 200 2080 1674 2136
rect 1730 2080 1735 2136
rect 200 2078 1735 2080
rect 200 2048 800 2078
rect 1669 2075 1735 2078
rect 37181 1458 37247 1461
rect 39200 1458 39800 1488
rect 37181 1456 39800 1458
rect 37181 1400 37186 1456
rect 37242 1400 39800 1456
rect 37181 1398 39800 1400
rect 37181 1395 37247 1398
rect 39200 1368 39800 1398
rect 200 778 800 808
rect 2773 778 2839 781
rect 200 776 2839 778
rect 200 720 2778 776
rect 2834 720 2839 776
rect 200 718 2839 720
rect 200 688 800 718
rect 2773 715 2839 718
rect 37273 778 37339 781
rect 39200 778 39800 808
rect 37273 776 39800 778
rect 37273 720 37278 776
rect 37334 720 39800 776
rect 37273 718 39800 720
rect 37273 715 37339 718
rect 39200 688 39800 718
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 12020 37360 12084 37364
rect 12020 37304 12034 37360
rect 12034 37304 12084 37360
rect 12020 37300 12084 37304
rect 20668 37300 20732 37364
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 2084 36348 2148 36412
rect 19380 36076 19444 36140
rect 7420 36000 7484 36004
rect 7420 35944 7434 36000
rect 7434 35944 7484 36000
rect 7420 35940 7484 35944
rect 20116 36000 20180 36004
rect 20116 35944 20130 36000
rect 20130 35944 20180 36000
rect 20116 35940 20180 35944
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 20668 32948 20732 33012
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 20300 32328 20364 32332
rect 20300 32272 20314 32328
rect 20314 32272 20364 32328
rect 20300 32268 20364 32272
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19380 31860 19444 31924
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 18828 31240 18892 31244
rect 18828 31184 18842 31240
rect 18842 31184 18892 31240
rect 18828 31180 18892 31184
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 20484 29412 20548 29476
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 1900 29004 1964 29068
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 5028 27704 5092 27708
rect 5028 27648 5042 27704
rect 5042 27648 5092 27704
rect 5028 27644 5092 27648
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 20668 26828 20732 26892
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 2268 26284 2332 26348
rect 5212 26284 5276 26348
rect 17908 26284 17972 26348
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 9812 25060 9876 25124
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 20668 24984 20732 24988
rect 20668 24928 20682 24984
rect 20682 24928 20732 24984
rect 20668 24924 20732 24928
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4844 23564 4908 23628
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 17908 22476 17972 22540
rect 5764 22340 5828 22404
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 20668 22204 20732 22268
rect 5396 22128 5460 22132
rect 5396 22072 5410 22128
rect 5410 22072 5460 22128
rect 5396 22068 5460 22072
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 20484 20436 20548 20500
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 18828 19756 18892 19820
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 3188 19348 3252 19412
rect 17908 19212 17972 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 5580 18804 5644 18868
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 7420 18124 7484 18188
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 8156 17852 8220 17916
rect 6868 17716 6932 17780
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 9812 15192 9876 15196
rect 9812 15136 9826 15192
rect 9826 15136 9876 15192
rect 9812 15132 9876 15136
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 2820 13772 2884 13836
rect 5396 13696 5460 13700
rect 5396 13640 5446 13696
rect 5446 13640 5460 13696
rect 5396 13636 5460 13640
rect 6868 13636 6932 13700
rect 12020 13636 12084 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 5580 12336 5644 12340
rect 5580 12280 5594 12336
rect 5594 12280 5644 12336
rect 5580 12276 5644 12280
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 5028 11868 5092 11932
rect 8156 11792 8220 11796
rect 8156 11736 8206 11792
rect 8206 11736 8220 11792
rect 8156 11732 8220 11736
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 5764 10916 5828 10980
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 3188 9556 3252 9620
rect 5212 9556 5276 9620
rect 20300 9556 20364 9620
rect 2820 9420 2884 9484
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 2084 9208 2148 9212
rect 2084 9152 2098 9208
rect 2098 9152 2148 9208
rect 2084 9148 2148 9152
rect 20116 8876 20180 8940
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 1900 6488 1964 6492
rect 1900 6432 1950 6488
rect 1950 6432 1964 6488
rect 1900 6428 1964 6432
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 2268 5884 2332 5948
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4844 3164 4908 3228
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 12019 37364 12085 37365
rect 12019 37300 12020 37364
rect 12084 37300 12085 37364
rect 12019 37299 12085 37300
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 2083 36412 2149 36413
rect 2083 36348 2084 36412
rect 2148 36348 2149 36412
rect 2083 36347 2149 36348
rect 1899 29068 1965 29069
rect 1899 29004 1900 29068
rect 1964 29004 1965 29068
rect 1899 29003 1965 29004
rect 1902 6493 1962 29003
rect 2086 9213 2146 36347
rect 4208 35392 4528 36416
rect 7419 36004 7485 36005
rect 7419 35940 7420 36004
rect 7484 35940 7485 36004
rect 7419 35939 7485 35940
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 5027 27708 5093 27709
rect 5027 27644 5028 27708
rect 5092 27644 5093 27708
rect 5027 27643 5093 27644
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 2267 26348 2333 26349
rect 2267 26284 2268 26348
rect 2332 26284 2333 26348
rect 2267 26283 2333 26284
rect 2083 9212 2149 9213
rect 2083 9148 2084 9212
rect 2148 9148 2149 9212
rect 2083 9147 2149 9148
rect 1899 6492 1965 6493
rect 1899 6428 1900 6492
rect 1964 6428 1965 6492
rect 1899 6427 1965 6428
rect 2270 5949 2330 26283
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4843 23628 4909 23629
rect 4843 23564 4844 23628
rect 4908 23564 4909 23628
rect 4843 23563 4909 23564
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 3187 19412 3253 19413
rect 3187 19348 3188 19412
rect 3252 19348 3253 19412
rect 3187 19347 3253 19348
rect 2819 13836 2885 13837
rect 2819 13772 2820 13836
rect 2884 13772 2885 13836
rect 2819 13771 2885 13772
rect 2822 9485 2882 13771
rect 3190 9621 3250 19347
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 3187 9620 3253 9621
rect 3187 9556 3188 9620
rect 3252 9556 3253 9620
rect 3187 9555 3253 9556
rect 2819 9484 2885 9485
rect 2819 9420 2820 9484
rect 2884 9420 2885 9484
rect 2819 9419 2885 9420
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 2267 5948 2333 5949
rect 2267 5884 2268 5948
rect 2332 5884 2333 5948
rect 2267 5883 2333 5884
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4846 3229 4906 23563
rect 5030 11933 5090 27643
rect 5211 26348 5277 26349
rect 5211 26284 5212 26348
rect 5276 26284 5277 26348
rect 5211 26283 5277 26284
rect 5027 11932 5093 11933
rect 5027 11868 5028 11932
rect 5092 11868 5093 11932
rect 5027 11867 5093 11868
rect 5214 9621 5274 26283
rect 5763 22404 5829 22405
rect 5763 22340 5764 22404
rect 5828 22340 5829 22404
rect 5763 22339 5829 22340
rect 5395 22132 5461 22133
rect 5395 22068 5396 22132
rect 5460 22068 5461 22132
rect 5395 22067 5461 22068
rect 5398 13701 5458 22067
rect 5579 18868 5645 18869
rect 5579 18804 5580 18868
rect 5644 18804 5645 18868
rect 5579 18803 5645 18804
rect 5395 13700 5461 13701
rect 5395 13636 5396 13700
rect 5460 13636 5461 13700
rect 5395 13635 5461 13636
rect 5582 12341 5642 18803
rect 5579 12340 5645 12341
rect 5579 12276 5580 12340
rect 5644 12276 5645 12340
rect 5579 12275 5645 12276
rect 5766 10981 5826 22339
rect 7422 18189 7482 35939
rect 9811 25124 9877 25125
rect 9811 25060 9812 25124
rect 9876 25060 9877 25124
rect 9811 25059 9877 25060
rect 7419 18188 7485 18189
rect 7419 18124 7420 18188
rect 7484 18124 7485 18188
rect 7419 18123 7485 18124
rect 8155 17916 8221 17917
rect 8155 17852 8156 17916
rect 8220 17852 8221 17916
rect 8155 17851 8221 17852
rect 6867 17780 6933 17781
rect 6867 17716 6868 17780
rect 6932 17716 6933 17780
rect 6867 17715 6933 17716
rect 6870 13701 6930 17715
rect 6867 13700 6933 13701
rect 6867 13636 6868 13700
rect 6932 13636 6933 13700
rect 6867 13635 6933 13636
rect 8158 11797 8218 17851
rect 9814 15197 9874 25059
rect 9811 15196 9877 15197
rect 9811 15132 9812 15196
rect 9876 15132 9877 15196
rect 9811 15131 9877 15132
rect 12022 13701 12082 37299
rect 19568 37024 19888 37584
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 20667 37364 20733 37365
rect 20667 37300 20668 37364
rect 20732 37300 20733 37364
rect 20667 37299 20733 37300
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19379 36140 19445 36141
rect 19379 36076 19380 36140
rect 19444 36076 19445 36140
rect 19379 36075 19445 36076
rect 19382 31925 19442 36075
rect 19568 35936 19888 36960
rect 20115 36004 20181 36005
rect 20115 35940 20116 36004
rect 20180 35940 20181 36004
rect 20115 35939 20181 35940
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19379 31924 19445 31925
rect 19379 31860 19380 31924
rect 19444 31860 19445 31924
rect 19379 31859 19445 31860
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 18827 31244 18893 31245
rect 18827 31180 18828 31244
rect 18892 31180 18893 31244
rect 18827 31179 18893 31180
rect 17907 26348 17973 26349
rect 17907 26284 17908 26348
rect 17972 26284 17973 26348
rect 17907 26283 17973 26284
rect 17910 22541 17970 26283
rect 17907 22540 17973 22541
rect 17907 22476 17908 22540
rect 17972 22476 17973 22540
rect 17907 22475 17973 22476
rect 17910 19277 17970 22475
rect 18830 19821 18890 31179
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 18827 19820 18893 19821
rect 18827 19756 18828 19820
rect 18892 19756 18893 19820
rect 18827 19755 18893 19756
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 17907 19276 17973 19277
rect 17907 19212 17908 19276
rect 17972 19212 17973 19276
rect 17907 19211 17973 19212
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 12019 13700 12085 13701
rect 12019 13636 12020 13700
rect 12084 13636 12085 13700
rect 12019 13635 12085 13636
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 8155 11796 8221 11797
rect 8155 11732 8156 11796
rect 8220 11732 8221 11796
rect 8155 11731 8221 11732
rect 5763 10980 5829 10981
rect 5763 10916 5764 10980
rect 5828 10916 5829 10980
rect 5763 10915 5829 10916
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 5211 9620 5277 9621
rect 5211 9556 5212 9620
rect 5276 9556 5277 9620
rect 5211 9555 5277 9556
rect 19568 8736 19888 9760
rect 20118 8941 20178 35939
rect 20670 33013 20730 37299
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 20667 33012 20733 33013
rect 20667 32948 20668 33012
rect 20732 32948 20733 33012
rect 20667 32947 20733 32948
rect 20299 32332 20365 32333
rect 20299 32268 20300 32332
rect 20364 32268 20365 32332
rect 20299 32267 20365 32268
rect 20302 9621 20362 32267
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 20483 29476 20549 29477
rect 20483 29412 20484 29476
rect 20548 29412 20549 29476
rect 20483 29411 20549 29412
rect 20486 20501 20546 29411
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 20667 26892 20733 26893
rect 20667 26828 20668 26892
rect 20732 26828 20733 26892
rect 20667 26827 20733 26828
rect 20670 24989 20730 26827
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 20667 24988 20733 24989
rect 20667 24924 20668 24988
rect 20732 24924 20733 24988
rect 20667 24923 20733 24924
rect 20670 22269 20730 24923
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 20667 22268 20733 22269
rect 20667 22204 20668 22268
rect 20732 22204 20733 22268
rect 20667 22203 20733 22204
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 20483 20500 20549 20501
rect 20483 20436 20484 20500
rect 20548 20436 20549 20500
rect 20483 20435 20549 20436
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 20299 9620 20365 9621
rect 20299 9556 20300 9620
rect 20364 9556 20365 9620
rect 20299 9555 20365 9556
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 20115 8940 20181 8941
rect 20115 8876 20116 8940
rect 20180 8876 20181 8940
rect 20115 8875 20181 8876
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 4843 3228 4909 3229
rect 4843 3164 4844 3228
rect 4908 3164 4909 3228
rect 4843 3163 4909 3164
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 13616 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform -1 0 2852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1667941163
transform -1 0 8280 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1667941163
transform -1 0 2944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1667941163
transform -1 0 2300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2392 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41
timestamp 1667941163
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49
timestamp 1667941163
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1667941163
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1667941163
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7544 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_105
timestamp 1667941163
transform 1 0 10764 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1667941163
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118
timestamp 1667941163
transform 1 0 11960 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_126 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12696 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132
timestamp 1667941163
transform 1 0 13248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149
timestamp 1667941163
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_154
timestamp 1667941163
transform 1 0 15272 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1667941163
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_174
timestamp 1667941163
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1667941163
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1667941163
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1667941163
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_202
timestamp 1667941163
transform 1 0 19688 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_210
timestamp 1667941163
transform 1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_216
timestamp 1667941163
transform 1 0 20976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1667941163
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_238
timestamp 1667941163
transform 1 0 23000 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1667941163
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_258
timestamp 1667941163
transform 1 0 24840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_266
timestamp 1667941163
transform 1 0 25576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_274
timestamp 1667941163
transform 1 0 26312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_286
timestamp 1667941163
transform 1 0 27416 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_294
timestamp 1667941163
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_300
timestamp 1667941163
transform 1 0 28704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_315
timestamp 1667941163
transform 1 0 30084 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_322
timestamp 1667941163
transform 1 0 30728 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1667941163
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_342
timestamp 1667941163
transform 1 0 32568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_350
timestamp 1667941163
transform 1 0 33304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_358
timestamp 1667941163
transform 1 0 34040 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_371
timestamp 1667941163
transform 1 0 35236 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_379
timestamp 1667941163
transform 1 0 35972 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1667941163
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1667941163
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_17
timestamp 1667941163
transform 1 0 2668 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_24
timestamp 1667941163
transform 1 0 3312 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_36
timestamp 1667941163
transform 1 0 4416 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_48
timestamp 1667941163
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_62
timestamp 1667941163
transform 1 0 6808 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_74
timestamp 1667941163
transform 1 0 7912 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_86
timestamp 1667941163
transform 1 0 9016 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_97
timestamp 1667941163
transform 1 0 10028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp 1667941163
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1667941163
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_132
timestamp 1667941163
transform 1 0 13248 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_140
timestamp 1667941163
transform 1 0 13984 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_147
timestamp 1667941163
transform 1 0 14628 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp 1667941163
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1667941163
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_176
timestamp 1667941163
transform 1 0 17296 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_188
timestamp 1667941163
transform 1 0 18400 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_200
timestamp 1667941163
transform 1 0 19504 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_212
timestamp 1667941163
transform 1 0 20608 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1667941163
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1667941163
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1667941163
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1667941163
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1667941163
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1667941163
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1667941163
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1667941163
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1667941163
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1667941163
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_385
timestamp 1667941163
transform 1 0 36524 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1667941163
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_9
timestamp 1667941163
transform 1 0 1932 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_13
timestamp 1667941163
transform 1 0 2300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_25
timestamp 1667941163
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1667941163
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1667941163
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1667941163
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1667941163
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1667941163
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1667941163
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_221
timestamp 1667941163
transform 1 0 21436 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_227
timestamp 1667941163
transform 1 0 21988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_239
timestamp 1667941163
transform 1 0 23092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1667941163
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1667941163
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1667941163
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_341
timestamp 1667941163
transform 1 0 32476 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_389
timestamp 1667941163
transform 1 0 36892 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_397
timestamp 1667941163
transform 1 0 37628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_8
timestamp 1667941163
transform 1 0 1840 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_20
timestamp 1667941163
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_32
timestamp 1667941163
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_44
timestamp 1667941163
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_61
timestamp 1667941163
transform 1 0 6716 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_65
timestamp 1667941163
transform 1 0 7084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_77
timestamp 1667941163
transform 1 0 8188 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_89
timestamp 1667941163
transform 1 0 9292 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_101
timestamp 1667941163
transform 1 0 10396 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_109
timestamp 1667941163
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1667941163
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1667941163
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1667941163
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1667941163
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1667941163
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_205
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_214
timestamp 1667941163
transform 1 0 20792 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1667941163
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1667941163
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1667941163
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_384
timestamp 1667941163
transform 1 0 36432 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_9
timestamp 1667941163
transform 1 0 1932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_21
timestamp 1667941163
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1667941163
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1667941163
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1667941163
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_401
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1667941163
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_8
timestamp 1667941163
transform 1 0 1840 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_20
timestamp 1667941163
transform 1 0 2944 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_32
timestamp 1667941163
transform 1 0 4048 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_44
timestamp 1667941163
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_177
timestamp 1667941163
transform 1 0 17388 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_192
timestamp 1667941163
transform 1 0 18768 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_204
timestamp 1667941163
transform 1 0 19872 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_216
timestamp 1667941163
transform 1 0 20976 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_316
timestamp 1667941163
transform 1 0 30176 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_328
timestamp 1667941163
transform 1 0 31280 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_11
timestamp 1667941163
transform 1 0 2116 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_18
timestamp 1667941163
transform 1 0 2760 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1667941163
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1667941163
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1667941163
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1667941163
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_146
timestamp 1667941163
transform 1 0 14536 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_158
timestamp 1667941163
transform 1 0 15640 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_170
timestamp 1667941163
transform 1 0 16744 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_182
timestamp 1667941163
transform 1 0 17848 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1667941163
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_268
timestamp 1667941163
transform 1 0 25760 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_280
timestamp 1667941163
transform 1 0 26864 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_291
timestamp 1667941163
transform 1 0 27876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_303
timestamp 1667941163
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1667941163
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_401
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_11
timestamp 1667941163
transform 1 0 2116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_23
timestamp 1667941163
transform 1 0 3220 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_35
timestamp 1667941163
transform 1 0 4324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1667941163
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_62
timestamp 1667941163
transform 1 0 6808 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_74
timestamp 1667941163
transform 1 0 7912 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_86
timestamp 1667941163
transform 1 0 9016 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_98
timestamp 1667941163
transform 1 0 10120 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1667941163
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_119
timestamp 1667941163
transform 1 0 12052 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_134
timestamp 1667941163
transform 1 0 13432 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_141
timestamp 1667941163
transform 1 0 14076 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_153
timestamp 1667941163
transform 1 0 15180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_160
timestamp 1667941163
transform 1 0 15824 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_177
timestamp 1667941163
transform 1 0 17388 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_187
timestamp 1667941163
transform 1 0 18308 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_191
timestamp 1667941163
transform 1 0 18676 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_203
timestamp 1667941163
transform 1 0 19780 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_215
timestamp 1667941163
transform 1 0 20884 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_261
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_265
timestamp 1667941163
transform 1 0 25484 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_272
timestamp 1667941163
transform 1 0 26128 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_401
timestamp 1667941163
transform 1 0 37996 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_8
timestamp 1667941163
transform 1 0 1840 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_20
timestamp 1667941163
transform 1 0 2944 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1667941163
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_59
timestamp 1667941163
transform 1 0 6532 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_63
timestamp 1667941163
transform 1 0 6900 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_75
timestamp 1667941163
transform 1 0 8004 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_116
timestamp 1667941163
transform 1 0 11776 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_125
timestamp 1667941163
transform 1 0 12604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1667941163
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_163
timestamp 1667941163
transform 1 0 16100 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_175
timestamp 1667941163
transform 1 0 17204 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_184
timestamp 1667941163
transform 1 0 18032 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_206
timestamp 1667941163
transform 1 0 20056 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_218
timestamp 1667941163
transform 1 0 21160 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_230
timestamp 1667941163
transform 1 0 22264 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_239
timestamp 1667941163
transform 1 0 23092 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_246
timestamp 1667941163
transform 1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1667941163
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1667941163
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1667941163
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_8
timestamp 1667941163
transform 1 0 1840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_15
timestamp 1667941163
transform 1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_32
timestamp 1667941163
transform 1 0 4048 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_44
timestamp 1667941163
transform 1 0 5152 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_62
timestamp 1667941163
transform 1 0 6808 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_74
timestamp 1667941163
transform 1 0 7912 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_86
timestamp 1667941163
transform 1 0 9016 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_98
timestamp 1667941163
transform 1 0 10120 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_106
timestamp 1667941163
transform 1 0 10856 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1667941163
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_124
timestamp 1667941163
transform 1 0 12512 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_136
timestamp 1667941163
transform 1 0 13616 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_144
timestamp 1667941163
transform 1 0 14352 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_150
timestamp 1667941163
transform 1 0 14904 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_162
timestamp 1667941163
transform 1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_180
timestamp 1667941163
transform 1 0 17664 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_184
timestamp 1667941163
transform 1 0 18032 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_198
timestamp 1667941163
transform 1 0 19320 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_211
timestamp 1667941163
transform 1 0 20516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1667941163
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_230
timestamp 1667941163
transform 1 0 22264 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_236
timestamp 1667941163
transform 1 0 22816 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_246
timestamp 1667941163
transform 1 0 23736 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_258
timestamp 1667941163
transform 1 0 24840 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_270
timestamp 1667941163
transform 1 0 25944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1667941163
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_9
timestamp 1667941163
transform 1 0 1932 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1667941163
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1667941163
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_34
timestamp 1667941163
transform 1 0 4232 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_46
timestamp 1667941163
transform 1 0 5336 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_58
timestamp 1667941163
transform 1 0 6440 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_70
timestamp 1667941163
transform 1 0 7544 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1667941163
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_102
timestamp 1667941163
transform 1 0 10488 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_114
timestamp 1667941163
transform 1 0 11592 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_125
timestamp 1667941163
transform 1 0 12604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_132
timestamp 1667941163
transform 1 0 13248 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_156
timestamp 1667941163
transform 1 0 15456 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_164
timestamp 1667941163
transform 1 0 16192 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_169
timestamp 1667941163
transform 1 0 16652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_181
timestamp 1667941163
transform 1 0 17756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1667941163
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_202
timestamp 1667941163
transform 1 0 19688 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_214
timestamp 1667941163
transform 1 0 20792 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_220
timestamp 1667941163
transform 1 0 21344 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_234
timestamp 1667941163
transform 1 0 22632 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_242
timestamp 1667941163
transform 1 0 23368 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_246
timestamp 1667941163
transform 1 0 23736 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_281
timestamp 1667941163
transform 1 0 26956 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_288
timestamp 1667941163
transform 1 0 27600 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_300
timestamp 1667941163
transform 1 0 28704 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_401
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1667941163
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_9
timestamp 1667941163
transform 1 0 1932 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_16
timestamp 1667941163
transform 1 0 2576 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_20
timestamp 1667941163
transform 1 0 2944 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_24
timestamp 1667941163
transform 1 0 3312 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_36
timestamp 1667941163
transform 1 0 4416 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_48
timestamp 1667941163
transform 1 0 5520 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1667941163
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1667941163
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_127
timestamp 1667941163
transform 1 0 12788 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_134
timestamp 1667941163
transform 1 0 13432 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_146
timestamp 1667941163
transform 1 0 14536 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_150
timestamp 1667941163
transform 1 0 14904 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_154
timestamp 1667941163
transform 1 0 15272 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_158
timestamp 1667941163
transform 1 0 15640 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp 1667941163
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_205
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_212
timestamp 1667941163
transform 1 0 20608 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1667941163
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_286
timestamp 1667941163
transform 1 0 27416 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_298
timestamp 1667941163
transform 1 0 28520 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_310
timestamp 1667941163
transform 1 0 29624 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_322
timestamp 1667941163
transform 1 0 30728 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1667941163
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_381
timestamp 1667941163
transform 1 0 36156 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_401
timestamp 1667941163
transform 1 0 37996 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_11
timestamp 1667941163
transform 1 0 2116 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_18
timestamp 1667941163
transform 1 0 2760 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 1667941163
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_122
timestamp 1667941163
transform 1 0 12328 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 1667941163
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_151
timestamp 1667941163
transform 1 0 14996 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_157
timestamp 1667941163
transform 1 0 15548 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_162
timestamp 1667941163
transform 1 0 16008 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_174
timestamp 1667941163
transform 1 0 17112 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_180
timestamp 1667941163
transform 1 0 17664 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_184
timestamp 1667941163
transform 1 0 18032 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_190
timestamp 1667941163
transform 1 0 18584 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1667941163
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_207
timestamp 1667941163
transform 1 0 20148 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_219
timestamp 1667941163
transform 1 0 21252 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_234
timestamp 1667941163
transform 1 0 22632 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_247
timestamp 1667941163
transform 1 0 23828 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_272
timestamp 1667941163
transform 1 0 26128 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_279
timestamp 1667941163
transform 1 0 26772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_291
timestamp 1667941163
transform 1 0 27876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_303
timestamp 1667941163
transform 1 0 28980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1667941163
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_382
timestamp 1667941163
transform 1 0 36248 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_394
timestamp 1667941163
transform 1 0 37352 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_406
timestamp 1667941163
transform 1 0 38456 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_9
timestamp 1667941163
transform 1 0 1932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_16
timestamp 1667941163
transform 1 0 2576 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_20
timestamp 1667941163
transform 1 0 2944 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_24
timestamp 1667941163
transform 1 0 3312 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_31
timestamp 1667941163
transform 1 0 3956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_43
timestamp 1667941163
transform 1 0 5060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_68
timestamp 1667941163
transform 1 0 7360 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_80
timestamp 1667941163
transform 1 0 8464 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_92
timestamp 1667941163
transform 1 0 9568 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_104
timestamp 1667941163
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_137
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_141
timestamp 1667941163
transform 1 0 14076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_145
timestamp 1667941163
transform 1 0 14444 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_153
timestamp 1667941163
transform 1 0 15180 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_162
timestamp 1667941163
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_189
timestamp 1667941163
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_193
timestamp 1667941163
transform 1 0 18860 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_197
timestamp 1667941163
transform 1 0 19228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_207
timestamp 1667941163
transform 1 0 20148 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1667941163
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_249
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_257
timestamp 1667941163
transform 1 0 24748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_263
timestamp 1667941163
transform 1 0 25300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_275
timestamp 1667941163
transform 1 0 26404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_291
timestamp 1667941163
transform 1 0 27876 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_303
timestamp 1667941163
transform 1 0 28980 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_315
timestamp 1667941163
transform 1 0 30084 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_319
timestamp 1667941163
transform 1 0 30452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_331
timestamp 1667941163
transform 1 0 31556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_9
timestamp 1667941163
transform 1 0 1932 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_13
timestamp 1667941163
transform 1 0 2300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1667941163
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_34
timestamp 1667941163
transform 1 0 4232 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_46
timestamp 1667941163
transform 1 0 5336 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_50
timestamp 1667941163
transform 1 0 5704 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_54
timestamp 1667941163
transform 1 0 6072 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_66
timestamp 1667941163
transform 1 0 7176 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_78
timestamp 1667941163
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1667941163
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_160
timestamp 1667941163
transform 1 0 15824 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_167
timestamp 1667941163
transform 1 0 16468 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_187
timestamp 1667941163
transform 1 0 18308 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1667941163
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_207
timestamp 1667941163
transform 1 0 20148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1667941163
transform 1 0 21252 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_223
timestamp 1667941163
transform 1 0 21620 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_240
timestamp 1667941163
transform 1 0 23184 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_244
timestamp 1667941163
transform 1 0 23552 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1667941163
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_261
timestamp 1667941163
transform 1 0 25116 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_272
timestamp 1667941163
transform 1 0 26128 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_284
timestamp 1667941163
transform 1 0 27232 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_296
timestamp 1667941163
transform 1 0 28336 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_405
timestamp 1667941163
transform 1 0 38364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_15
timestamp 1667941163
transform 1 0 2484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_22
timestamp 1667941163
transform 1 0 3128 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_29
timestamp 1667941163
transform 1 0 3772 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_38
timestamp 1667941163
transform 1 0 4600 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_45
timestamp 1667941163
transform 1 0 5244 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1667941163
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_62
timestamp 1667941163
transform 1 0 6808 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_74
timestamp 1667941163
transform 1 0 7912 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_86
timestamp 1667941163
transform 1 0 9016 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_98
timestamp 1667941163
transform 1 0 10120 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1667941163
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_118
timestamp 1667941163
transform 1 0 11960 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_130
timestamp 1667941163
transform 1 0 13064 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_142
timestamp 1667941163
transform 1 0 14168 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_149
timestamp 1667941163
transform 1 0 14812 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_156
timestamp 1667941163
transform 1 0 15456 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_177
timestamp 1667941163
transform 1 0 17388 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_182
timestamp 1667941163
transform 1 0 17848 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_189
timestamp 1667941163
transform 1 0 18492 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_193
timestamp 1667941163
transform 1 0 18860 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_203
timestamp 1667941163
transform 1 0 19780 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_211
timestamp 1667941163
transform 1 0 20516 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_216
timestamp 1667941163
transform 1 0 20976 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_230
timestamp 1667941163
transform 1 0 22264 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_237
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_244
timestamp 1667941163
transform 1 0 23552 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_251
timestamp 1667941163
transform 1 0 24196 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_258
timestamp 1667941163
transform 1 0 24840 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_265
timestamp 1667941163
transform 1 0 25484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1667941163
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_288
timestamp 1667941163
transform 1 0 27600 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_297
timestamp 1667941163
transform 1 0 28428 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_309
timestamp 1667941163
transform 1 0 29532 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_321
timestamp 1667941163
transform 1 0 30636 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_333
timestamp 1667941163
transform 1 0 31740 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_8
timestamp 1667941163
transform 1 0 1840 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_25
timestamp 1667941163
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_37
timestamp 1667941163
transform 1 0 4508 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_52
timestamp 1667941163
transform 1 0 5888 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_58
timestamp 1667941163
transform 1 0 6440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_62
timestamp 1667941163
transform 1 0 6808 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_69
timestamp 1667941163
transform 1 0 7452 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1667941163
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_92
timestamp 1667941163
transform 1 0 9568 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_99
timestamp 1667941163
transform 1 0 10212 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_112
timestamp 1667941163
transform 1 0 11408 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_119
timestamp 1667941163
transform 1 0 12052 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_131
timestamp 1667941163
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_152
timestamp 1667941163
transform 1 0 15088 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_162
timestamp 1667941163
transform 1 0 16008 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_187
timestamp 1667941163
transform 1 0 18308 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_209
timestamp 1667941163
transform 1 0 20332 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_223
timestamp 1667941163
transform 1 0 21620 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_235
timestamp 1667941163
transform 1 0 22724 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_247
timestamp 1667941163
transform 1 0 23828 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_264
timestamp 1667941163
transform 1 0 25392 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_276
timestamp 1667941163
transform 1 0 26496 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_284
timestamp 1667941163
transform 1 0 27232 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_288
timestamp 1667941163
transform 1 0 27600 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_297
timestamp 1667941163
transform 1 0 28428 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_305
timestamp 1667941163
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_401
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_405
timestamp 1667941163
transform 1 0 38364 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1667941163
transform 1 0 1748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_11
timestamp 1667941163
transform 1 0 2116 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_24
timestamp 1667941163
transform 1 0 3312 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_31
timestamp 1667941163
transform 1 0 3956 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_38
timestamp 1667941163
transform 1 0 4600 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_46
timestamp 1667941163
transform 1 0 5336 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_68
timestamp 1667941163
transform 1 0 7360 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_77
timestamp 1667941163
transform 1 0 8188 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_94
timestamp 1667941163
transform 1 0 9752 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_102
timestamp 1667941163
transform 1 0 10488 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1667941163
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1667941163
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_137
timestamp 1667941163
transform 1 0 13708 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_143
timestamp 1667941163
transform 1 0 14260 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_150
timestamp 1667941163
transform 1 0 14904 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_162
timestamp 1667941163
transform 1 0 16008 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_174
timestamp 1667941163
transform 1 0 17112 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_186
timestamp 1667941163
transform 1 0 18216 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_198
timestamp 1667941163
transform 1 0 19320 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_210
timestamp 1667941163
transform 1 0 20424 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1667941163
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_230
timestamp 1667941163
transform 1 0 22264 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_242
timestamp 1667941163
transform 1 0 23368 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_254
timestamp 1667941163
transform 1 0 24472 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1667941163
transform 1 0 25852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_277
timestamp 1667941163
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_285
timestamp 1667941163
transform 1 0 27324 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_289
timestamp 1667941163
transform 1 0 27692 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_302
timestamp 1667941163
transform 1 0 28888 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_314
timestamp 1667941163
transform 1 0 29992 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_326
timestamp 1667941163
transform 1 0 31096 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 1667941163
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_9
timestamp 1667941163
transform 1 0 1932 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_16
timestamp 1667941163
transform 1 0 2576 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1667941163
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_44
timestamp 1667941163
transform 1 0 5152 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_51
timestamp 1667941163
transform 1 0 5796 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_66
timestamp 1667941163
transform 1 0 7176 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_78
timestamp 1667941163
transform 1 0 8280 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_113
timestamp 1667941163
transform 1 0 11500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_117
timestamp 1667941163
transform 1 0 11868 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_126
timestamp 1667941163
transform 1 0 12696 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1667941163
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1667941163
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_152
timestamp 1667941163
transform 1 0 15088 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_160
timestamp 1667941163
transform 1 0 15824 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_164
timestamp 1667941163
transform 1 0 16192 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_176
timestamp 1667941163
transform 1 0 17296 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_188
timestamp 1667941163
transform 1 0 18400 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_203
timestamp 1667941163
transform 1 0 19780 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_217
timestamp 1667941163
transform 1 0 21068 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_229
timestamp 1667941163
transform 1 0 22172 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_242
timestamp 1667941163
transform 1 0 23368 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_249
timestamp 1667941163
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_264
timestamp 1667941163
transform 1 0 25392 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_272
timestamp 1667941163
transform 1 0 26128 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_284
timestamp 1667941163
transform 1 0 27232 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_296
timestamp 1667941163
transform 1 0 28336 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1667941163
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1667941163
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1667941163
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_14
timestamp 1667941163
transform 1 0 2392 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_21
timestamp 1667941163
transform 1 0 3036 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_28
timestamp 1667941163
transform 1 0 3680 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_35
timestamp 1667941163
transform 1 0 4324 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_41
timestamp 1667941163
transform 1 0 4876 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1667941163
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1667941163
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_63
timestamp 1667941163
transform 1 0 6900 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_73
timestamp 1667941163
transform 1 0 7820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_85
timestamp 1667941163
transform 1 0 8924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_97
timestamp 1667941163
transform 1 0 10028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 1667941163
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1667941163
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_152
timestamp 1667941163
transform 1 0 15088 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_159
timestamp 1667941163
transform 1 0 15732 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1667941163
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_174
timestamp 1667941163
transform 1 0 17112 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_178
timestamp 1667941163
transform 1 0 17480 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_188
timestamp 1667941163
transform 1 0 18400 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_195
timestamp 1667941163
transform 1 0 19044 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_207
timestamp 1667941163
transform 1 0 20148 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_212
timestamp 1667941163
transform 1 0 20608 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_231
timestamp 1667941163
transform 1 0 22356 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_238
timestamp 1667941163
transform 1 0 23000 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_253
timestamp 1667941163
transform 1 0 24380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_265
timestamp 1667941163
transform 1 0 25484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1667941163
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_301
timestamp 1667941163
transform 1 0 28796 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_307
timestamp 1667941163
transform 1 0 29348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_319
timestamp 1667941163
transform 1 0 30452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_331
timestamp 1667941163
transform 1 0 31556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1667941163
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_342
timestamp 1667941163
transform 1 0 32568 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_354
timestamp 1667941163
transform 1 0 33672 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_366
timestamp 1667941163
transform 1 0 34776 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_378
timestamp 1667941163
transform 1 0 35880 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_390
timestamp 1667941163
transform 1 0 36984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_401
timestamp 1667941163
transform 1 0 37996 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_9
timestamp 1667941163
transform 1 0 1932 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_18
timestamp 1667941163
transform 1 0 2760 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_22
timestamp 1667941163
transform 1 0 3128 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1667941163
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_34
timestamp 1667941163
transform 1 0 4232 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_52
timestamp 1667941163
transform 1 0 5888 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_64
timestamp 1667941163
transform 1 0 6992 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_68
timestamp 1667941163
transform 1 0 7360 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_72
timestamp 1667941163
transform 1 0 7728 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_79
timestamp 1667941163
transform 1 0 8372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_92
timestamp 1667941163
transform 1 0 9568 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_107
timestamp 1667941163
transform 1 0 10948 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_119
timestamp 1667941163
transform 1 0 12052 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_131
timestamp 1667941163
transform 1 0 13156 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1667941163
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_160
timestamp 1667941163
transform 1 0 15824 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_177
timestamp 1667941163
transform 1 0 17388 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1667941163
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_209
timestamp 1667941163
transform 1 0 20332 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_217
timestamp 1667941163
transform 1 0 21068 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_223
timestamp 1667941163
transform 1 0 21620 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_230
timestamp 1667941163
transform 1 0 22264 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1667941163
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1667941163
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_265
timestamp 1667941163
transform 1 0 25484 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_272
timestamp 1667941163
transform 1 0 26128 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_279
timestamp 1667941163
transform 1 0 26772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_291
timestamp 1667941163
transform 1 0 27876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1667941163
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_332
timestamp 1667941163
transform 1 0 31648 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_344
timestamp 1667941163
transform 1 0 32752 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_356
timestamp 1667941163
transform 1 0 33856 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_405
timestamp 1667941163
transform 1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1667941163
transform 1 0 1748 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_12
timestamp 1667941163
transform 1 0 2208 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_18
timestamp 1667941163
transform 1 0 2760 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_22
timestamp 1667941163
transform 1 0 3128 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_39
timestamp 1667941163
transform 1 0 4692 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_46
timestamp 1667941163
transform 1 0 5336 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1667941163
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_62
timestamp 1667941163
transform 1 0 6808 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_68
timestamp 1667941163
transform 1 0 7360 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_82
timestamp 1667941163
transform 1 0 8648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_95
timestamp 1667941163
transform 1 0 9844 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1667941163
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_124
timestamp 1667941163
transform 1 0 12512 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_136
timestamp 1667941163
transform 1 0 13616 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_146
timestamp 1667941163
transform 1 0 14536 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_158
timestamp 1667941163
transform 1 0 15640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1667941163
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_174
timestamp 1667941163
transform 1 0 17112 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_181
timestamp 1667941163
transform 1 0 17756 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_198
timestamp 1667941163
transform 1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_211
timestamp 1667941163
transform 1 0 20516 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_218
timestamp 1667941163
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_230
timestamp 1667941163
transform 1 0 22264 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_242
timestamp 1667941163
transform 1 0 23368 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_251
timestamp 1667941163
transform 1 0 24196 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_263
timestamp 1667941163
transform 1 0 25300 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_267
timestamp 1667941163
transform 1 0 25668 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_277
timestamp 1667941163
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_303
timestamp 1667941163
transform 1 0 28980 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_315
timestamp 1667941163
transform 1 0 30084 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_321
timestamp 1667941163
transform 1 0 30636 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_325
timestamp 1667941163
transform 1 0 31004 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_333
timestamp 1667941163
transform 1 0 31740 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_9
timestamp 1667941163
transform 1 0 1932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_19
timestamp 1667941163
transform 1 0 2852 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1667941163
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_34
timestamp 1667941163
transform 1 0 4232 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_40
timestamp 1667941163
transform 1 0 4784 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_49
timestamp 1667941163
transform 1 0 5612 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_66
timestamp 1667941163
transform 1 0 7176 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_70
timestamp 1667941163
transform 1 0 7544 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_74
timestamp 1667941163
transform 1 0 7912 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1667941163
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_91
timestamp 1667941163
transform 1 0 9476 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_104
timestamp 1667941163
transform 1 0 10672 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_129
timestamp 1667941163
transform 1 0 12972 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_133
timestamp 1667941163
transform 1 0 13340 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1667941163
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_154
timestamp 1667941163
transform 1 0 15272 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_160
timestamp 1667941163
transform 1 0 15824 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_174
timestamp 1667941163
transform 1 0 17112 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_186
timestamp 1667941163
transform 1 0 18216 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1667941163
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_208
timestamp 1667941163
transform 1 0 20240 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_220
timestamp 1667941163
transform 1 0 21344 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_232
timestamp 1667941163
transform 1 0 22448 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_240
timestamp 1667941163
transform 1 0 23184 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1667941163
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_268
timestamp 1667941163
transform 1 0 25760 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_280
timestamp 1667941163
transform 1 0 26864 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_292
timestamp 1667941163
transform 1 0 27968 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_300
timestamp 1667941163
transform 1 0 28704 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1667941163
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_315
timestamp 1667941163
transform 1 0 30084 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_329
timestamp 1667941163
transform 1 0 31372 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_336
timestamp 1667941163
transform 1 0 32016 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_348
timestamp 1667941163
transform 1 0 33120 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_360
timestamp 1667941163
transform 1 0 34224 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_405
timestamp 1667941163
transform 1 0 38364 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_16
timestamp 1667941163
transform 1 0 2576 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_28
timestamp 1667941163
transform 1 0 3680 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_35
timestamp 1667941163
transform 1 0 4324 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_42
timestamp 1667941163
transform 1 0 4968 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_49
timestamp 1667941163
transform 1 0 5612 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_72
timestamp 1667941163
transform 1 0 7728 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_79
timestamp 1667941163
transform 1 0 8372 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_86
timestamp 1667941163
transform 1 0 9016 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_97
timestamp 1667941163
transform 1 0 10028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1667941163
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_129
timestamp 1667941163
transform 1 0 12972 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_136
timestamp 1667941163
transform 1 0 13616 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_144
timestamp 1667941163
transform 1 0 14352 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_153
timestamp 1667941163
transform 1 0 15180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1667941163
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_176
timestamp 1667941163
transform 1 0 17296 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_188
timestamp 1667941163
transform 1 0 18400 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_195
timestamp 1667941163
transform 1 0 19044 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_207
timestamp 1667941163
transform 1 0 20148 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1667941163
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_237
timestamp 1667941163
transform 1 0 22908 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_250
timestamp 1667941163
transform 1 0 24104 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_260
timestamp 1667941163
transform 1 0 25024 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_272
timestamp 1667941163
transform 1 0 26128 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1667941163
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_291
timestamp 1667941163
transform 1 0 27876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_303
timestamp 1667941163
transform 1 0 28980 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_308
timestamp 1667941163
transform 1 0 29440 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_315
timestamp 1667941163
transform 1 0 30084 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_327
timestamp 1667941163
transform 1 0 31188 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1667941163
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_369
timestamp 1667941163
transform 1 0 35052 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_402
timestamp 1667941163
transform 1 0 38088 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_406
timestamp 1667941163
transform 1 0 38456 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_9
timestamp 1667941163
transform 1 0 1932 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_19
timestamp 1667941163
transform 1 0 2852 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1667941163
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_34
timestamp 1667941163
transform 1 0 4232 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_38
timestamp 1667941163
transform 1 0 4600 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_42
timestamp 1667941163
transform 1 0 4968 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_49
timestamp 1667941163
transform 1 0 5612 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_56
timestamp 1667941163
transform 1 0 6256 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_63
timestamp 1667941163
transform 1 0 6900 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_71
timestamp 1667941163
transform 1 0 7636 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_75
timestamp 1667941163
transform 1 0 8004 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1667941163
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_90
timestamp 1667941163
transform 1 0 9384 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_105
timestamp 1667941163
transform 1 0 10764 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_117
timestamp 1667941163
transform 1 0 11868 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_121
timestamp 1667941163
transform 1 0 12236 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1667941163
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_148
timestamp 1667941163
transform 1 0 14720 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_154
timestamp 1667941163
transform 1 0 15272 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_158
timestamp 1667941163
transform 1 0 15640 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_165
timestamp 1667941163
transform 1 0 16284 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_172
timestamp 1667941163
transform 1 0 16928 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_180
timestamp 1667941163
transform 1 0 17664 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_186
timestamp 1667941163
transform 1 0 18216 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1667941163
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_201
timestamp 1667941163
transform 1 0 19596 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_206
timestamp 1667941163
transform 1 0 20056 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_219
timestamp 1667941163
transform 1 0 21252 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_231
timestamp 1667941163
transform 1 0 22356 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_246
timestamp 1667941163
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1667941163
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_277
timestamp 1667941163
transform 1 0 26588 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_283
timestamp 1667941163
transform 1 0 27140 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_297
timestamp 1667941163
transform 1 0 28428 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_305
timestamp 1667941163
transform 1 0 29164 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1667941163
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1667941163
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1667941163
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1667941163
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_17
timestamp 1667941163
transform 1 0 2668 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_32
timestamp 1667941163
transform 1 0 4048 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_39
timestamp 1667941163
transform 1 0 4692 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_43
timestamp 1667941163
transform 1 0 5060 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_47
timestamp 1667941163
transform 1 0 5428 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1667941163
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_62
timestamp 1667941163
transform 1 0 6808 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_74
timestamp 1667941163
transform 1 0 7912 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_78
timestamp 1667941163
transform 1 0 8280 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_89
timestamp 1667941163
transform 1 0 9292 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_96
timestamp 1667941163
transform 1 0 9936 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_103
timestamp 1667941163
transform 1 0 10580 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1667941163
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1667941163
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1667941163
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1667941163
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1667941163
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1667941163
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_174
timestamp 1667941163
transform 1 0 17112 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_182
timestamp 1667941163
transform 1 0 17848 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_197
timestamp 1667941163
transform 1 0 19228 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_205
timestamp 1667941163
transform 1 0 19964 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_214
timestamp 1667941163
transform 1 0 20792 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1667941163
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_237
timestamp 1667941163
transform 1 0 22908 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_241
timestamp 1667941163
transform 1 0 23276 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_253
timestamp 1667941163
transform 1 0 24380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_265
timestamp 1667941163
transform 1 0 25484 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_269
timestamp 1667941163
transform 1 0 25852 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_277
timestamp 1667941163
transform 1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_292
timestamp 1667941163
transform 1 0 27968 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_300
timestamp 1667941163
transform 1 0 28704 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_304
timestamp 1667941163
transform 1 0 29072 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_312
timestamp 1667941163
transform 1 0 29808 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1667941163
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1667941163
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1667941163
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_15
timestamp 1667941163
transform 1 0 2484 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_22
timestamp 1667941163
transform 1 0 3128 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_34
timestamp 1667941163
transform 1 0 4232 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_46
timestamp 1667941163
transform 1 0 5336 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_51
timestamp 1667941163
transform 1 0 5796 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_59
timestamp 1667941163
transform 1 0 6532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_64
timestamp 1667941163
transform 1 0 6992 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_71
timestamp 1667941163
transform 1 0 7636 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_75
timestamp 1667941163
transform 1 0 8004 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_79
timestamp 1667941163
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_96
timestamp 1667941163
transform 1 0 9936 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_104
timestamp 1667941163
transform 1 0 10672 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_109
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_116
timestamp 1667941163
transform 1 0 11776 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_123
timestamp 1667941163
transform 1 0 12420 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1667941163
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_146
timestamp 1667941163
transform 1 0 14536 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_158
timestamp 1667941163
transform 1 0 15640 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_170
timestamp 1667941163
transform 1 0 16744 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_182
timestamp 1667941163
transform 1 0 17848 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1667941163
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_205
timestamp 1667941163
transform 1 0 19964 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_209
timestamp 1667941163
transform 1 0 20332 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_217
timestamp 1667941163
transform 1 0 21068 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_221
timestamp 1667941163
transform 1 0 21436 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_229
timestamp 1667941163
transform 1 0 22172 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_239
timestamp 1667941163
transform 1 0 23092 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_246
timestamp 1667941163
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_258
timestamp 1667941163
transform 1 0 24840 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_265
timestamp 1667941163
transform 1 0 25484 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_274
timestamp 1667941163
transform 1 0 26312 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_286
timestamp 1667941163
transform 1 0 27416 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_293
timestamp 1667941163
transform 1 0 28060 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1667941163
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_319
timestamp 1667941163
transform 1 0 30452 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_331
timestamp 1667941163
transform 1 0 31556 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_343
timestamp 1667941163
transform 1 0 32660 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_355
timestamp 1667941163
transform 1 0 33764 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_405
timestamp 1667941163
transform 1 0 38364 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_9
timestamp 1667941163
transform 1 0 1932 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_16
timestamp 1667941163
transform 1 0 2576 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_28
timestamp 1667941163
transform 1 0 3680 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_40
timestamp 1667941163
transform 1 0 4784 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1667941163
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1667941163
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_137
timestamp 1667941163
transform 1 0 13708 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_144
timestamp 1667941163
transform 1 0 14352 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_156
timestamp 1667941163
transform 1 0 15456 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_174
timestamp 1667941163
transform 1 0 17112 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_180
timestamp 1667941163
transform 1 0 17664 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_184
timestamp 1667941163
transform 1 0 18032 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_196
timestamp 1667941163
transform 1 0 19136 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_208
timestamp 1667941163
transform 1 0 20240 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_214
timestamp 1667941163
transform 1 0 20792 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_218
timestamp 1667941163
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1667941163
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_249
timestamp 1667941163
transform 1 0 24012 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_255
timestamp 1667941163
transform 1 0 24564 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_259
timestamp 1667941163
transform 1 0 24932 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_266
timestamp 1667941163
transform 1 0 25576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1667941163
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_286
timestamp 1667941163
transform 1 0 27416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_290
timestamp 1667941163
transform 1 0 27784 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_299
timestamp 1667941163
transform 1 0 28612 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_324
timestamp 1667941163
transform 1 0 30912 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_25
timestamp 1667941163
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_74
timestamp 1667941163
transform 1 0 7912 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1667941163
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_90
timestamp 1667941163
transform 1 0 9384 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_98
timestamp 1667941163
transform 1 0 10120 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_102
timestamp 1667941163
transform 1 0 10488 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_131
timestamp 1667941163
transform 1 0 13156 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1667941163
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_149
timestamp 1667941163
transform 1 0 14812 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_175
timestamp 1667941163
transform 1 0 17204 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_187
timestamp 1667941163
transform 1 0 18308 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1667941163
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_201
timestamp 1667941163
transform 1 0 19596 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_215
timestamp 1667941163
transform 1 0 20884 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_221
timestamp 1667941163
transform 1 0 21436 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_225
timestamp 1667941163
transform 1 0 21804 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_242
timestamp 1667941163
transform 1 0 23368 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1667941163
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_258
timestamp 1667941163
transform 1 0 24840 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_262
timestamp 1667941163
transform 1 0 25208 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_266
timestamp 1667941163
transform 1 0 25576 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_275
timestamp 1667941163
transform 1 0 26404 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_287
timestamp 1667941163
transform 1 0 27508 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_293
timestamp 1667941163
transform 1 0 28060 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_301
timestamp 1667941163
transform 1 0 28796 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 1667941163
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_319
timestamp 1667941163
transform 1 0 30452 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_331
timestamp 1667941163
transform 1 0 31556 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_343
timestamp 1667941163
transform 1 0 32660 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_355
timestamp 1667941163
transform 1 0 33764 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_9
timestamp 1667941163
transform 1 0 1932 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_15
timestamp 1667941163
transform 1 0 2484 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1667941163
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1667941163
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1667941163
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_97
timestamp 1667941163
transform 1 0 10028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1667941163
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_125
timestamp 1667941163
transform 1 0 12604 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_151
timestamp 1667941163
transform 1 0 14996 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1667941163
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1667941163
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_191
timestamp 1667941163
transform 1 0 18676 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_216
timestamp 1667941163
transform 1 0 20976 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_237
timestamp 1667941163
transform 1 0 22908 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_258
timestamp 1667941163
transform 1 0 24840 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_270
timestamp 1667941163
transform 1 0 25944 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1667941163
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_305
timestamp 1667941163
transform 1 0 29164 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_309
timestamp 1667941163
transform 1 0 29532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_313
timestamp 1667941163
transform 1 0 29900 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_325
timestamp 1667941163
transform 1 0 31004 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_333
timestamp 1667941163
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_345
timestamp 1667941163
transform 1 0 32844 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_351
timestamp 1667941163
transform 1 0 33396 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_363
timestamp 1667941163
transform 1 0 34500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_375
timestamp 1667941163
transform 1 0 35604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_387
timestamp 1667941163
transform 1 0 36708 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1667941163
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_35
timestamp 1667941163
transform 1 0 4324 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_56
timestamp 1667941163
transform 1 0 6256 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1667941163
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1667941163
transform 1 0 9476 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_113
timestamp 1667941163
transform 1 0 11500 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_117
timestamp 1667941163
transform 1 0 11868 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1667941163
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_153
timestamp 1667941163
transform 1 0 15180 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_178
timestamp 1667941163
transform 1 0 17480 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_190
timestamp 1667941163
transform 1 0 18584 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_212
timestamp 1667941163
transform 1 0 20608 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_220
timestamp 1667941163
transform 1 0 21344 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_228
timestamp 1667941163
transform 1 0 22080 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_232
timestamp 1667941163
transform 1 0 22448 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_236
timestamp 1667941163
transform 1 0 22816 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_240
timestamp 1667941163
transform 1 0 23184 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1667941163
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1667941163
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1667941163
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1667941163
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_320
timestamp 1667941163
transform 1 0 30544 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_332
timestamp 1667941163
transform 1 0 31648 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_344
timestamp 1667941163
transform 1 0 32752 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_356
timestamp 1667941163
transform 1 0 33856 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1667941163
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_25
timestamp 1667941163
transform 1 0 3404 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_33
timestamp 1667941163
transform 1 0 4140 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1667941163
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_79
timestamp 1667941163
transform 1 0 8372 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_87
timestamp 1667941163
transform 1 0 9108 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1667941163
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_118
timestamp 1667941163
transform 1 0 11960 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_130
timestamp 1667941163
transform 1 0 13064 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_142
timestamp 1667941163
transform 1 0 14168 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1667941163
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1667941163
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_193
timestamp 1667941163
transform 1 0 18860 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_201
timestamp 1667941163
transform 1 0 19596 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_207
timestamp 1667941163
transform 1 0 20148 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_219
timestamp 1667941163
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1667941163
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_240
timestamp 1667941163
transform 1 0 23184 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_247
timestamp 1667941163
transform 1 0 23828 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_259
timestamp 1667941163
transform 1 0 24932 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_271
timestamp 1667941163
transform 1 0 26036 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1667941163
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1667941163
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_317
timestamp 1667941163
transform 1 0 30268 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_326
timestamp 1667941163
transform 1 0 31096 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1667941163
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_341
timestamp 1667941163
transform 1 0 32476 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_345
timestamp 1667941163
transform 1 0 32844 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_357
timestamp 1667941163
transform 1 0 33948 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_369
timestamp 1667941163
transform 1 0 35052 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_381
timestamp 1667941163
transform 1 0 36156 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_389
timestamp 1667941163
transform 1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_401
timestamp 1667941163
transform 1 0 37996 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1667941163
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_49
timestamp 1667941163
transform 1 0 5612 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_72
timestamp 1667941163
transform 1 0 7728 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_110
timestamp 1667941163
transform 1 0 11224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_135
timestamp 1667941163
transform 1 0 13524 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1667941163
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_149
timestamp 1667941163
transform 1 0 14812 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_172
timestamp 1667941163
transform 1 0 16928 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_184
timestamp 1667941163
transform 1 0 18032 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_209
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_223
timestamp 1667941163
transform 1 0 21620 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_236
timestamp 1667941163
transform 1 0 22816 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1667941163
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1667941163
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_298
timestamp 1667941163
transform 1 0 28520 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1667941163
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_327
timestamp 1667941163
transform 1 0 31188 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_331
timestamp 1667941163
transform 1 0 31556 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_343
timestamp 1667941163
transform 1 0 32660 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_355
timestamp 1667941163
transform 1 0 33764 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_8
timestamp 1667941163
transform 1 0 1840 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_16
timestamp 1667941163
transform 1 0 2576 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_37
timestamp 1667941163
transform 1 0 4508 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_49
timestamp 1667941163
transform 1 0 5612 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1667941163
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_88
timestamp 1667941163
transform 1 0 9200 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_100
timestamp 1667941163
transform 1 0 10304 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_126
timestamp 1667941163
transform 1 0 12696 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_134
timestamp 1667941163
transform 1 0 13432 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_148
timestamp 1667941163
transform 1 0 14720 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_160
timestamp 1667941163
transform 1 0 15824 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1667941163
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1667941163
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_205
timestamp 1667941163
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_215
timestamp 1667941163
transform 1 0 20884 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1667941163
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_230
timestamp 1667941163
transform 1 0 22264 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_242
timestamp 1667941163
transform 1 0 23368 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_254
timestamp 1667941163
transform 1 0 24472 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_266
timestamp 1667941163
transform 1 0 25576 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_270
timestamp 1667941163
transform 1 0 25944 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1667941163
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_287
timestamp 1667941163
transform 1 0 27508 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_294
timestamp 1667941163
transform 1 0 28152 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_302
timestamp 1667941163
transform 1 0 28888 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_314
timestamp 1667941163
transform 1 0 29992 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_318
timestamp 1667941163
transform 1 0 30360 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_322
timestamp 1667941163
transform 1 0 30728 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1667941163
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_9
timestamp 1667941163
transform 1 0 1932 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_21
timestamp 1667941163
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1667941163
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_63
timestamp 1667941163
transform 1 0 6900 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_75
timestamp 1667941163
transform 1 0 8004 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1667941163
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_107
timestamp 1667941163
transform 1 0 10948 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_119
timestamp 1667941163
transform 1 0 12052 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_131
timestamp 1667941163
transform 1 0 13156 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1667941163
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_149
timestamp 1667941163
transform 1 0 14812 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_171
timestamp 1667941163
transform 1 0 16836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_183
timestamp 1667941163
transform 1 0 17940 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1667941163
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_214
timestamp 1667941163
transform 1 0 20792 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1667941163
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1667941163
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1667941163
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1667941163
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_281
timestamp 1667941163
transform 1 0 26956 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_293
timestamp 1667941163
transform 1 0 28060 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_298
timestamp 1667941163
transform 1 0 28520 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_302
timestamp 1667941163
transform 1 0 28888 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_306
timestamp 1667941163
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_320
timestamp 1667941163
transform 1 0 30544 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_327
timestamp 1667941163
transform 1 0 31188 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_334
timestamp 1667941163
transform 1 0 31832 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_346
timestamp 1667941163
transform 1 0 32936 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_358
timestamp 1667941163
transform 1 0 34040 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_405
timestamp 1667941163
transform 1 0 38364 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1667941163
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1667941163
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_39
timestamp 1667941163
transform 1 0 4692 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1667941163
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_89
timestamp 1667941163
transform 1 0 9292 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_101
timestamp 1667941163
transform 1 0 10396 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_109
timestamp 1667941163
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1667941163
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_137
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1667941163
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_181
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_190
timestamp 1667941163
transform 1 0 18584 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_200
timestamp 1667941163
transform 1 0 19504 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_215
timestamp 1667941163
transform 1 0 20884 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1667941163
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_233
timestamp 1667941163
transform 1 0 22540 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_244
timestamp 1667941163
transform 1 0 23552 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_251
timestamp 1667941163
transform 1 0 24196 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_258
timestamp 1667941163
transform 1 0 24840 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_270
timestamp 1667941163
transform 1 0 25944 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1667941163
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_301
timestamp 1667941163
transform 1 0 28796 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_308
timestamp 1667941163
transform 1 0 29440 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_320
timestamp 1667941163
transform 1 0 30544 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_328
timestamp 1667941163
transform 1 0 31280 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_333
timestamp 1667941163
transform 1 0 31740 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_9
timestamp 1667941163
transform 1 0 1932 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_21
timestamp 1667941163
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_63
timestamp 1667941163
transform 1 0 6900 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_75
timestamp 1667941163
transform 1 0 8004 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1667941163
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_107
timestamp 1667941163
transform 1 0 10948 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_115
timestamp 1667941163
transform 1 0 11684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1667941163
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1667941163
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1667941163
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_177
timestamp 1667941163
transform 1 0 17388 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_185
timestamp 1667941163
transform 1 0 18124 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1667941163
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_202
timestamp 1667941163
transform 1 0 19688 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_212
timestamp 1667941163
transform 1 0 20608 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_229
timestamp 1667941163
transform 1 0 22172 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_236
timestamp 1667941163
transform 1 0 22816 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_243
timestamp 1667941163
transform 1 0 23460 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1667941163
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_268
timestamp 1667941163
transform 1 0 25760 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_275
timestamp 1667941163
transform 1 0 26404 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_287
timestamp 1667941163
transform 1 0 27508 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_299
timestamp 1667941163
transform 1 0 28612 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_314
timestamp 1667941163
transform 1 0 29992 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_326
timestamp 1667941163
transform 1 0 31096 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_338
timestamp 1667941163
transform 1 0 32200 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_350
timestamp 1667941163
transform 1 0 33304 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1667941163
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_401
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_26
timestamp 1667941163
transform 1 0 3496 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1667941163
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1667941163
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_125
timestamp 1667941163
transform 1 0 12604 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_131
timestamp 1667941163
transform 1 0 13156 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_155
timestamp 1667941163
transform 1 0 15364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1667941163
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_181
timestamp 1667941163
transform 1 0 17756 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_185
timestamp 1667941163
transform 1 0 18124 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_195
timestamp 1667941163
transform 1 0 19044 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1667941163
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1667941163
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_236
timestamp 1667941163
transform 1 0 22816 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_248
timestamp 1667941163
transform 1 0 23920 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_260
timestamp 1667941163
transform 1 0 25024 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_271
timestamp 1667941163
transform 1 0 26036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1667941163
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_296
timestamp 1667941163
transform 1 0 28336 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_303
timestamp 1667941163
transform 1 0 28980 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_315
timestamp 1667941163
transform 1 0 30084 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_323
timestamp 1667941163
transform 1 0 30820 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1667941163
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_357
timestamp 1667941163
transform 1 0 33948 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_363
timestamp 1667941163
transform 1 0 34500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_375
timestamp 1667941163
transform 1 0 35604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_387
timestamp 1667941163
transform 1 0 36708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1667941163
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_49
timestamp 1667941163
transform 1 0 5612 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_70
timestamp 1667941163
transform 1 0 7544 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1667941163
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_101
timestamp 1667941163
transform 1 0 10396 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_123
timestamp 1667941163
transform 1 0 12420 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_135
timestamp 1667941163
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1667941163
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_153
timestamp 1667941163
transform 1 0 15180 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_179
timestamp 1667941163
transform 1 0 17572 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_191
timestamp 1667941163
transform 1 0 18676 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1667941163
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_205
timestamp 1667941163
transform 1 0 19964 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_213
timestamp 1667941163
transform 1 0 20700 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_219
timestamp 1667941163
transform 1 0 21252 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_231
timestamp 1667941163
transform 1 0 22356 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_243
timestamp 1667941163
transform 1 0 23460 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1667941163
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_269
timestamp 1667941163
transform 1 0 25852 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_278
timestamp 1667941163
transform 1 0 26680 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_290
timestamp 1667941163
transform 1 0 27784 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_302
timestamp 1667941163
transform 1 0 28888 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_324
timestamp 1667941163
transform 1 0 30912 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_336
timestamp 1667941163
transform 1 0 32016 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_348
timestamp 1667941163
transform 1 0 33120 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_360
timestamp 1667941163
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_10
timestamp 1667941163
transform 1 0 2024 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_17
timestamp 1667941163
transform 1 0 2668 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_29
timestamp 1667941163
transform 1 0 3772 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_33
timestamp 1667941163
transform 1 0 4140 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1667941163
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_73
timestamp 1667941163
transform 1 0 7820 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_95
timestamp 1667941163
transform 1 0 9844 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_107
timestamp 1667941163
transform 1 0 10948 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1667941163
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1667941163
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1667941163
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_149
timestamp 1667941163
transform 1 0 14812 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1667941163
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_174
timestamp 1667941163
transform 1 0 17112 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_182
timestamp 1667941163
transform 1 0 17848 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1667941163
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_205
timestamp 1667941163
transform 1 0 19964 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_214
timestamp 1667941163
transform 1 0 20792 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1667941163
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_230
timestamp 1667941163
transform 1 0 22264 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_237
timestamp 1667941163
transform 1 0 22908 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_243
timestamp 1667941163
transform 1 0 23460 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_247
timestamp 1667941163
transform 1 0 23828 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_255
timestamp 1667941163
transform 1 0 24564 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_263
timestamp 1667941163
transform 1 0 25300 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1667941163
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_287
timestamp 1667941163
transform 1 0 27508 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_301
timestamp 1667941163
transform 1 0 28796 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_310
timestamp 1667941163
transform 1 0 29624 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_322
timestamp 1667941163
transform 1 0 30728 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1667941163
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_357
timestamp 1667941163
transform 1 0 33948 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_363
timestamp 1667941163
transform 1 0 34500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_375
timestamp 1667941163
transform 1 0 35604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_387
timestamp 1667941163
transform 1 0 36708 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1667941163
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_54
timestamp 1667941163
transform 1 0 6072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_78
timestamp 1667941163
transform 1 0 8280 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1667941163
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1667941163
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1667941163
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_153
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_176
timestamp 1667941163
transform 1 0 17296 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_184
timestamp 1667941163
transform 1 0 18032 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1667941163
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1667941163
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_209
timestamp 1667941163
transform 1 0 20332 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_220
timestamp 1667941163
transform 1 0 21344 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_237
timestamp 1667941163
transform 1 0 22908 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_249
timestamp 1667941163
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_258
timestamp 1667941163
transform 1 0 24840 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_270
timestamp 1667941163
transform 1 0 25944 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_282
timestamp 1667941163
transform 1 0 27048 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_293
timestamp 1667941163
transform 1 0 28060 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1667941163
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1667941163
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1667941163
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_8
timestamp 1667941163
transform 1 0 1840 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_20
timestamp 1667941163
transform 1 0 2944 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_32
timestamp 1667941163
transform 1 0 4048 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_38
timestamp 1667941163
transform 1 0 4600 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_50
timestamp 1667941163
transform 1 0 5704 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_77
timestamp 1667941163
transform 1 0 8188 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_100
timestamp 1667941163
transform 1 0 10304 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_126
timestamp 1667941163
transform 1 0 12696 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_133
timestamp 1667941163
transform 1 0 13340 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_41_162
timestamp 1667941163
transform 1 0 16008 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_184
timestamp 1667941163
transform 1 0 18032 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_198
timestamp 1667941163
transform 1 0 19320 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_206
timestamp 1667941163
transform 1 0 20056 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_211
timestamp 1667941163
transform 1 0 20516 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_218
timestamp 1667941163
transform 1 0 21160 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_233
timestamp 1667941163
transform 1 0 22540 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_244
timestamp 1667941163
transform 1 0 23552 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_251
timestamp 1667941163
transform 1 0 24196 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_263
timestamp 1667941163
transform 1 0 25300 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_269
timestamp 1667941163
transform 1 0 25852 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_277
timestamp 1667941163
transform 1 0 26588 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_298
timestamp 1667941163
transform 1 0 28520 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_302
timestamp 1667941163
transform 1 0 28888 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_306
timestamp 1667941163
transform 1 0 29256 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_318
timestamp 1667941163
transform 1 0 30360 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_330
timestamp 1667941163
transform 1 0 31464 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_9
timestamp 1667941163
transform 1 0 1932 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_21
timestamp 1667941163
transform 1 0 3036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_81
timestamp 1667941163
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_107
timestamp 1667941163
transform 1 0 10948 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_115
timestamp 1667941163
transform 1 0 11684 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1667941163
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_153
timestamp 1667941163
transform 1 0 15180 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_182
timestamp 1667941163
transform 1 0 17848 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_190
timestamp 1667941163
transform 1 0 18584 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1667941163
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_205
timestamp 1667941163
transform 1 0 19964 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_211
timestamp 1667941163
transform 1 0 20516 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_215
timestamp 1667941163
transform 1 0 20884 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_227
timestamp 1667941163
transform 1 0 21988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_239
timestamp 1667941163
transform 1 0 23092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1667941163
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_286
timestamp 1667941163
transform 1 0 27416 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_294
timestamp 1667941163
transform 1 0 28152 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_299
timestamp 1667941163
transform 1 0 28612 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 1667941163
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_314
timestamp 1667941163
transform 1 0 29992 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_326
timestamp 1667941163
transform 1 0 31096 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_338
timestamp 1667941163
transform 1 0 32200 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_350
timestamp 1667941163
transform 1 0 33304 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp 1667941163
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_401
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_19
timestamp 1667941163
transform 1 0 2852 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_23
timestamp 1667941163
transform 1 0 3220 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_47
timestamp 1667941163
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_73
timestamp 1667941163
transform 1 0 7820 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_85
timestamp 1667941163
transform 1 0 8924 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1667941163
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_135
timestamp 1667941163
transform 1 0 13524 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_147
timestamp 1667941163
transform 1 0 14628 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_159
timestamp 1667941163
transform 1 0 15732 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1667941163
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_192
timestamp 1667941163
transform 1 0 18768 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_200
timestamp 1667941163
transform 1 0 19504 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_204
timestamp 1667941163
transform 1 0 19872 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_211
timestamp 1667941163
transform 1 0 20516 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1667941163
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_231
timestamp 1667941163
transform 1 0 22356 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_238
timestamp 1667941163
transform 1 0 23000 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_245
timestamp 1667941163
transform 1 0 23644 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_257
timestamp 1667941163
transform 1 0 24748 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_269
timestamp 1667941163
transform 1 0 25852 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_277
timestamp 1667941163
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_296
timestamp 1667941163
transform 1 0 28336 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_307
timestamp 1667941163
transform 1 0 29348 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_321
timestamp 1667941163
transform 1 0 30636 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_333
timestamp 1667941163
transform 1 0 31740 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_346
timestamp 1667941163
transform 1 0 32936 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_358
timestamp 1667941163
transform 1 0 34040 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_370
timestamp 1667941163
transform 1 0 35144 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_382
timestamp 1667941163
transform 1 0 36248 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_390
timestamp 1667941163
transform 1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_9
timestamp 1667941163
transform 1 0 1932 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_23
timestamp 1667941163
transform 1 0 3220 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1667941163
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_117
timestamp 1667941163
transform 1 0 11868 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1667941163
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_153
timestamp 1667941163
transform 1 0 15180 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_182
timestamp 1667941163
transform 1 0 17848 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_190
timestamp 1667941163
transform 1 0 18584 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1667941163
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_212
timestamp 1667941163
transform 1 0 20608 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_224
timestamp 1667941163
transform 1 0 21712 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_236
timestamp 1667941163
transform 1 0 22816 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_242
timestamp 1667941163
transform 1 0 23368 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_249
timestamp 1667941163
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_262
timestamp 1667941163
transform 1 0 25208 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_269
timestamp 1667941163
transform 1 0 25852 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_282
timestamp 1667941163
transform 1 0 27048 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_294
timestamp 1667941163
transform 1 0 28152 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1667941163
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_337
timestamp 1667941163
transform 1 0 32108 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_350
timestamp 1667941163
transform 1 0 33304 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_362
timestamp 1667941163
transform 1 0 34408 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_401
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_405
timestamp 1667941163
transform 1 0 38364 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_8
timestamp 1667941163
transform 1 0 1840 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_20
timestamp 1667941163
transform 1 0 2944 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_32
timestamp 1667941163
transform 1 0 4048 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1667941163
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_65
timestamp 1667941163
transform 1 0 7084 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_86
timestamp 1667941163
transform 1 0 9016 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1667941163
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1667941163
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1667941163
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1667941163
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_175
timestamp 1667941163
transform 1 0 17204 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_179
timestamp 1667941163
transform 1 0 17572 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_196
timestamp 1667941163
transform 1 0 19136 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_203
timestamp 1667941163
transform 1 0 19780 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_210
timestamp 1667941163
transform 1 0 20424 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1667941163
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_230
timestamp 1667941163
transform 1 0 22264 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_254
timestamp 1667941163
transform 1 0 24472 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_262
timestamp 1667941163
transform 1 0 25208 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_269
timestamp 1667941163
transform 1 0 25852 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_277
timestamp 1667941163
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_292
timestamp 1667941163
transform 1 0 27968 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_299
timestamp 1667941163
transform 1 0 28612 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_308
timestamp 1667941163
transform 1 0 29440 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_320
timestamp 1667941163
transform 1 0 30544 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_332
timestamp 1667941163
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_357
timestamp 1667941163
transform 1 0 33948 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_362
timestamp 1667941163
transform 1 0 34408 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_374
timestamp 1667941163
transform 1 0 35512 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_386
timestamp 1667941163
transform 1 0 36616 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_9
timestamp 1667941163
transform 1 0 1932 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_21
timestamp 1667941163
transform 1 0 3036 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_123
timestamp 1667941163
transform 1 0 12420 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_135
timestamp 1667941163
transform 1 0 13524 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1667941163
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1667941163
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1667941163
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_177
timestamp 1667941163
transform 1 0 17388 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_191
timestamp 1667941163
transform 1 0 18676 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_214
timestamp 1667941163
transform 1 0 20792 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_240
timestamp 1667941163
transform 1 0 23184 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_247
timestamp 1667941163
transform 1 0 23828 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_258
timestamp 1667941163
transform 1 0 24840 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_266
timestamp 1667941163
transform 1 0 25576 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_281
timestamp 1667941163
transform 1 0 26956 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_293
timestamp 1667941163
transform 1 0 28060 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_305
timestamp 1667941163
transform 1 0 29164 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_314
timestamp 1667941163
transform 1 0 29992 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_326
timestamp 1667941163
transform 1 0 31096 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_338
timestamp 1667941163
transform 1 0 32200 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_350
timestamp 1667941163
transform 1 0 33304 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_362
timestamp 1667941163
transform 1 0 34408 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_405
timestamp 1667941163
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_43
timestamp 1667941163
transform 1 0 5060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_109
timestamp 1667941163
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_133
timestamp 1667941163
transform 1 0 13340 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_136
timestamp 1667941163
transform 1 0 13616 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1667941163
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1667941163
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_193
timestamp 1667941163
transform 1 0 18860 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_200
timestamp 1667941163
transform 1 0 19504 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_207
timestamp 1667941163
transform 1 0 20148 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_214
timestamp 1667941163
transform 1 0 20792 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_221
timestamp 1667941163
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_237
timestamp 1667941163
transform 1 0 22908 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_244
timestamp 1667941163
transform 1 0 23552 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_250
timestamp 1667941163
transform 1 0 24104 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_254
timestamp 1667941163
transform 1 0 24472 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_261
timestamp 1667941163
transform 1 0 25116 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_268
timestamp 1667941163
transform 1 0 25760 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_275
timestamp 1667941163
transform 1 0 26404 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1667941163
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_292
timestamp 1667941163
transform 1 0 27968 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_304
timestamp 1667941163
transform 1 0 29072 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_316
timestamp 1667941163
transform 1 0 30176 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_328
timestamp 1667941163
transform 1 0 31280 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_401
timestamp 1667941163
transform 1 0 37996 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_7
timestamp 1667941163
transform 1 0 1748 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_11
timestamp 1667941163
transform 1 0 2116 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_23
timestamp 1667941163
transform 1 0 3220 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_64
timestamp 1667941163
transform 1 0 6992 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_76
timestamp 1667941163
transform 1 0 8096 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_113
timestamp 1667941163
transform 1 0 11500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_135
timestamp 1667941163
transform 1 0 13524 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_159
timestamp 1667941163
transform 1 0 15732 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_181
timestamp 1667941163
transform 1 0 17756 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_193
timestamp 1667941163
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_202
timestamp 1667941163
transform 1 0 19688 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_220
timestamp 1667941163
transform 1 0 21344 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_232
timestamp 1667941163
transform 1 0 22448 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_236
timestamp 1667941163
transform 1 0 22816 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1667941163
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_258
timestamp 1667941163
transform 1 0 24840 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_282
timestamp 1667941163
transform 1 0 27048 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_295
timestamp 1667941163
transform 1 0 28244 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_302
timestamp 1667941163
transform 1 0 28888 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_330
timestamp 1667941163
transform 1 0 31464 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_347
timestamp 1667941163
transform 1 0 33028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_359
timestamp 1667941163
transform 1 0 34132 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_8
timestamp 1667941163
transform 1 0 1840 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_37
timestamp 1667941163
transform 1 0 4508 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_41
timestamp 1667941163
transform 1 0 4876 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1667941163
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1667941163
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_135
timestamp 1667941163
transform 1 0 13524 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_143
timestamp 1667941163
transform 1 0 14260 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_165
timestamp 1667941163
transform 1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_196
timestamp 1667941163
transform 1 0 19136 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1667941163
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_233
timestamp 1667941163
transform 1 0 22540 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_245
timestamp 1667941163
transform 1 0 23644 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_259
timestamp 1667941163
transform 1 0 24932 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1667941163
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_286
timestamp 1667941163
transform 1 0 27416 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_298
timestamp 1667941163
transform 1 0 28520 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_310
timestamp 1667941163
transform 1 0 29624 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_322
timestamp 1667941163
transform 1 0 30728 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_334
timestamp 1667941163
transform 1 0 31832 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_37
timestamp 1667941163
transform 1 0 4508 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1667941163
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1667941163
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_107
timestamp 1667941163
transform 1 0 10948 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_122
timestamp 1667941163
transform 1 0 12328 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_134
timestamp 1667941163
transform 1 0 13432 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_161
timestamp 1667941163
transform 1 0 15916 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_183
timestamp 1667941163
transform 1 0 17940 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1667941163
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_202
timestamp 1667941163
transform 1 0 19688 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_215
timestamp 1667941163
transform 1 0 20884 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_219
timestamp 1667941163
transform 1 0 21252 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_226
timestamp 1667941163
transform 1 0 21896 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_233
timestamp 1667941163
transform 1 0 22540 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_240
timestamp 1667941163
transform 1 0 23184 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_247
timestamp 1667941163
transform 1 0 23828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1667941163
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_257
timestamp 1667941163
transform 1 0 24748 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_271
timestamp 1667941163
transform 1 0 26036 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_278
timestamp 1667941163
transform 1 0 26680 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_285
timestamp 1667941163
transform 1 0 27324 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_291
timestamp 1667941163
transform 1 0 27876 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_300
timestamp 1667941163
transform 1 0 28704 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_314
timestamp 1667941163
transform 1 0 29992 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_325
timestamp 1667941163
transform 1 0 31004 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_337
timestamp 1667941163
transform 1 0 32108 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_349
timestamp 1667941163
transform 1 0 33212 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_361
timestamp 1667941163
transform 1 0 34316 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_370
timestamp 1667941163
transform 1 0 35144 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_382
timestamp 1667941163
transform 1 0 36248 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_394
timestamp 1667941163
transform 1 0 37352 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_405
timestamp 1667941163
transform 1 0 38364 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_9
timestamp 1667941163
transform 1 0 1932 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_21
timestamp 1667941163
transform 1 0 3036 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_33
timestamp 1667941163
transform 1 0 4140 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_45
timestamp 1667941163
transform 1 0 5244 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_53
timestamp 1667941163
transform 1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_91
timestamp 1667941163
transform 1 0 9476 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_106
timestamp 1667941163
transform 1 0 10856 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_125
timestamp 1667941163
transform 1 0 12604 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_147
timestamp 1667941163
transform 1 0 14628 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1667941163
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_191
timestamp 1667941163
transform 1 0 18676 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_202
timestamp 1667941163
transform 1 0 19688 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_209
timestamp 1667941163
transform 1 0 20332 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_216
timestamp 1667941163
transform 1 0 20976 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_232
timestamp 1667941163
transform 1 0 22448 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_240
timestamp 1667941163
transform 1 0 23184 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_245
timestamp 1667941163
transform 1 0 23644 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_253
timestamp 1667941163
transform 1 0 24380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_270
timestamp 1667941163
transform 1 0 25944 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_277
timestamp 1667941163
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_286
timestamp 1667941163
transform 1 0 27416 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_298
timestamp 1667941163
transform 1 0 28520 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_302
timestamp 1667941163
transform 1 0 28888 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_309
timestamp 1667941163
transform 1 0 29532 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_321
timestamp 1667941163
transform 1 0 30636 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_333
timestamp 1667941163
transform 1 0 31740 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1667941163
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_51
timestamp 1667941163
transform 1 0 5796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_78
timestamp 1667941163
transform 1 0 8280 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_122
timestamp 1667941163
transform 1 0 12328 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_134
timestamp 1667941163
transform 1 0 13432 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_159
timestamp 1667941163
transform 1 0 15732 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_180
timestamp 1667941163
transform 1 0 17664 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_188
timestamp 1667941163
transform 1 0 18400 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1667941163
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_206
timestamp 1667941163
transform 1 0 20056 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_214
timestamp 1667941163
transform 1 0 20792 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_218
timestamp 1667941163
transform 1 0 21160 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_235
timestamp 1667941163
transform 1 0 22724 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_242
timestamp 1667941163
transform 1 0 23368 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_249
timestamp 1667941163
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_271
timestamp 1667941163
transform 1 0 26036 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_285
timestamp 1667941163
transform 1 0 27324 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_299
timestamp 1667941163
transform 1 0 28612 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_401
timestamp 1667941163
transform 1 0 37996 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_405
timestamp 1667941163
transform 1 0 38364 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_42
timestamp 1667941163
transform 1 0 4968 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1667941163
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_91
timestamp 1667941163
transform 1 0 9476 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_103
timestamp 1667941163
transform 1 0 10580 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_138
timestamp 1667941163
transform 1 0 13800 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_150
timestamp 1667941163
transform 1 0 14904 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_162
timestamp 1667941163
transform 1 0 16008 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_176
timestamp 1667941163
transform 1 0 17296 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_201
timestamp 1667941163
transform 1 0 19596 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_206
timestamp 1667941163
transform 1 0 20056 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_213
timestamp 1667941163
transform 1 0 20700 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1667941163
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_235
timestamp 1667941163
transform 1 0 22724 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_239
timestamp 1667941163
transform 1 0 23092 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_243
timestamp 1667941163
transform 1 0 23460 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_250
timestamp 1667941163
transform 1 0 24104 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_258
timestamp 1667941163
transform 1 0 24840 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_274
timestamp 1667941163
transform 1 0 26312 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_285
timestamp 1667941163
transform 1 0 27324 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_294
timestamp 1667941163
transform 1 0 28152 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_306
timestamp 1667941163
transform 1 0 29256 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_315
timestamp 1667941163
transform 1 0 30084 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_322
timestamp 1667941163
transform 1 0 30728 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_334
timestamp 1667941163
transform 1 0 31832 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_9
timestamp 1667941163
transform 1 0 1932 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_16
timestamp 1667941163
transform 1 0 2576 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_110
timestamp 1667941163
transform 1 0 11224 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1667941163
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_161
timestamp 1667941163
transform 1 0 15916 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_182
timestamp 1667941163
transform 1 0 17848 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_190
timestamp 1667941163
transform 1 0 18584 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1667941163
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_208
timestamp 1667941163
transform 1 0 20240 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_215
timestamp 1667941163
transform 1 0 20884 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_227
timestamp 1667941163
transform 1 0 21988 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_235
timestamp 1667941163
transform 1 0 22724 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_246
timestamp 1667941163
transform 1 0 23736 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_261
timestamp 1667941163
transform 1 0 25116 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_266
timestamp 1667941163
transform 1 0 25576 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_283
timestamp 1667941163
transform 1 0 27140 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_290
timestamp 1667941163
transform 1 0 27784 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_297
timestamp 1667941163
transform 1 0 28428 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_305
timestamp 1667941163
transform 1 0 29164 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_9
timestamp 1667941163
transform 1 0 1932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_21
timestamp 1667941163
transform 1 0 3036 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_33
timestamp 1667941163
transform 1 0 4140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1667941163
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1667941163
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_70
timestamp 1667941163
transform 1 0 7544 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_82
timestamp 1667941163
transform 1 0 8648 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_110
timestamp 1667941163
transform 1 0 11224 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_117
timestamp 1667941163
transform 1 0 11868 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_129
timestamp 1667941163
transform 1 0 12972 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_141
timestamp 1667941163
transform 1 0 14076 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_165
timestamp 1667941163
transform 1 0 16284 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_191
timestamp 1667941163
transform 1 0 18676 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_195
timestamp 1667941163
transform 1 0 19044 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_199
timestamp 1667941163
transform 1 0 19412 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_212
timestamp 1667941163
transform 1 0 20608 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_230
timestamp 1667941163
transform 1 0 22264 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_241
timestamp 1667941163
transform 1 0 23276 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_255
timestamp 1667941163
transform 1 0 24564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_268
timestamp 1667941163
transform 1 0 25760 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_272
timestamp 1667941163
transform 1 0 26128 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_276
timestamp 1667941163
transform 1 0 26496 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_286
timestamp 1667941163
transform 1 0 27416 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_298
timestamp 1667941163
transform 1 0 28520 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_7
timestamp 1667941163
transform 1 0 1748 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_12
timestamp 1667941163
transform 1 0 2208 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_24
timestamp 1667941163
transform 1 0 3312 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_81
timestamp 1667941163
transform 1 0 8556 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_105
timestamp 1667941163
transform 1 0 10764 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_130
timestamp 1667941163
transform 1 0 13064 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1667941163
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_156
timestamp 1667941163
transform 1 0 15456 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_180
timestamp 1667941163
transform 1 0 17664 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1667941163
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_206
timestamp 1667941163
transform 1 0 20056 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_213
timestamp 1667941163
transform 1 0 20700 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_217
timestamp 1667941163
transform 1 0 21068 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_231
timestamp 1667941163
transform 1 0 22356 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_239
timestamp 1667941163
transform 1 0 23092 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_244
timestamp 1667941163
transform 1 0 23552 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_258
timestamp 1667941163
transform 1 0 24840 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_284
timestamp 1667941163
transform 1 0 27232 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1667941163
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_405
timestamp 1667941163
transform 1 0 38364 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_9
timestamp 1667941163
transform 1 0 1932 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_30
timestamp 1667941163
transform 1 0 3864 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 1667941163
transform 1 0 6072 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_89
timestamp 1667941163
transform 1 0 9292 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_104
timestamp 1667941163
transform 1 0 10672 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_191
timestamp 1667941163
transform 1 0 18676 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_199
timestamp 1667941163
transform 1 0 19412 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_203
timestamp 1667941163
transform 1 0 19780 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_222
timestamp 1667941163
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_233
timestamp 1667941163
transform 1 0 22540 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_238
timestamp 1667941163
transform 1 0 23000 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_244
timestamp 1667941163
transform 1 0 23552 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_256
timestamp 1667941163
transform 1 0 24656 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_263
timestamp 1667941163
transform 1 0 25300 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_270
timestamp 1667941163
transform 1 0 25944 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1667941163
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_292
timestamp 1667941163
transform 1 0 27968 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_299
timestamp 1667941163
transform 1 0 28612 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_306
timestamp 1667941163
transform 1 0 29256 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_313
timestamp 1667941163
transform 1 0 29900 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_325
timestamp 1667941163
transform 1 0 31004 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_333
timestamp 1667941163
transform 1 0 31740 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_9
timestamp 1667941163
transform 1 0 1932 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_16
timestamp 1667941163
transform 1 0 2576 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_69
timestamp 1667941163
transform 1 0 7452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_81
timestamp 1667941163
transform 1 0 8556 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_89
timestamp 1667941163
transform 1 0 9292 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_110
timestamp 1667941163
transform 1 0 11224 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_116
timestamp 1667941163
transform 1 0 11776 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1667941163
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_183
timestamp 1667941163
transform 1 0 17940 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_187
timestamp 1667941163
transform 1 0 18308 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_194
timestamp 1667941163
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_203
timestamp 1667941163
transform 1 0 19780 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_210
timestamp 1667941163
transform 1 0 20424 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_217
timestamp 1667941163
transform 1 0 21068 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_225
timestamp 1667941163
transform 1 0 21804 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_230
timestamp 1667941163
transform 1 0 22264 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_243
timestamp 1667941163
transform 1 0 23460 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_261
timestamp 1667941163
transform 1 0 25116 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_292
timestamp 1667941163
transform 1 0 27968 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_299
timestamp 1667941163
transform 1 0 28612 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_385
timestamp 1667941163
transform 1 0 36524 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_8
timestamp 1667941163
transform 1 0 1840 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_20
timestamp 1667941163
transform 1 0 2944 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_43
timestamp 1667941163
transform 1 0 5060 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_47
timestamp 1667941163
transform 1 0 5428 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1667941163
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1667941163
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_89
timestamp 1667941163
transform 1 0 9292 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_95
timestamp 1667941163
transform 1 0 9844 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_107
timestamp 1667941163
transform 1 0 10948 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_138
timestamp 1667941163
transform 1 0 13800 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_150
timestamp 1667941163
transform 1 0 14904 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_162
timestamp 1667941163
transform 1 0 16008 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_175
timestamp 1667941163
transform 1 0 17204 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_179
timestamp 1667941163
transform 1 0 17572 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_186
timestamp 1667941163
transform 1 0 18216 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_200
timestamp 1667941163
transform 1 0 19504 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_209
timestamp 1667941163
transform 1 0 20332 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_216
timestamp 1667941163
transform 1 0 20976 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_244
timestamp 1667941163
transform 1 0 23552 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_251
timestamp 1667941163
transform 1 0 24196 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_264
timestamp 1667941163
transform 1 0 25392 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_272
timestamp 1667941163
transform 1 0 26128 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_278
timestamp 1667941163
transform 1 0 26680 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_292
timestamp 1667941163
transform 1 0 27968 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_299
timestamp 1667941163
transform 1 0 28612 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_311
timestamp 1667941163
transform 1 0 29716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_323
timestamp 1667941163
transform 1 0 30820 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_9
timestamp 1667941163
transform 1 0 1932 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_21
timestamp 1667941163
transform 1 0 3036 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_37
timestamp 1667941163
transform 1 0 4508 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_59
timestamp 1667941163
transform 1 0 6532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_71
timestamp 1667941163
transform 1 0 7636 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_82
timestamp 1667941163
transform 1 0 8648 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_96
timestamp 1667941163
transform 1 0 9936 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_108
timestamp 1667941163
transform 1 0 11040 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_114
timestamp 1667941163
transform 1 0 11592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1667941163
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_146
timestamp 1667941163
transform 1 0 14536 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_158
timestamp 1667941163
transform 1 0 15640 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_182
timestamp 1667941163
transform 1 0 17848 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_190
timestamp 1667941163
transform 1 0 18584 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_194
timestamp 1667941163
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_203
timestamp 1667941163
transform 1 0 19780 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_207
timestamp 1667941163
transform 1 0 20148 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_214
timestamp 1667941163
transform 1 0 20792 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_228
timestamp 1667941163
transform 1 0 22080 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_236
timestamp 1667941163
transform 1 0 22816 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1667941163
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_258
timestamp 1667941163
transform 1 0 24840 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_262
timestamp 1667941163
transform 1 0 25208 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_266
timestamp 1667941163
transform 1 0 25576 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_272
timestamp 1667941163
transform 1 0 26128 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_282
timestamp 1667941163
transform 1 0 27048 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_290
timestamp 1667941163
transform 1 0 27784 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_306
timestamp 1667941163
transform 1 0 29256 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_372
timestamp 1667941163
transform 1 0 35328 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_384
timestamp 1667941163
transform 1 0 36432 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_392
timestamp 1667941163
transform 1 0 37168 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_398
timestamp 1667941163
transform 1 0 37720 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_406
timestamp 1667941163
transform 1 0 38456 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_26
timestamp 1667941163
transform 1 0 3496 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_38
timestamp 1667941163
transform 1 0 4600 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_50
timestamp 1667941163
transform 1 0 5704 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1667941163
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_83
timestamp 1667941163
transform 1 0 8740 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1667941163
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_121
timestamp 1667941163
transform 1 0 12236 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_126
timestamp 1667941163
transform 1 0 12696 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_138
timestamp 1667941163
transform 1 0 13800 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_142
timestamp 1667941163
transform 1 0 14168 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_166
timestamp 1667941163
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_191
timestamp 1667941163
transform 1 0 18676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_200
timestamp 1667941163
transform 1 0 19504 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_207
timestamp 1667941163
transform 1 0 20148 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1667941163
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_231
timestamp 1667941163
transform 1 0 22356 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_235
timestamp 1667941163
transform 1 0 22724 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_248
timestamp 1667941163
transform 1 0 23920 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_255
timestamp 1667941163
transform 1 0 24564 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_271
timestamp 1667941163
transform 1 0 26036 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_278
timestamp 1667941163
transform 1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_286
timestamp 1667941163
transform 1 0 27416 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_292
timestamp 1667941163
transform 1 0 27968 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_296
timestamp 1667941163
transform 1 0 28336 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_303
timestamp 1667941163
transform 1 0 28980 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_315
timestamp 1667941163
transform 1 0 30084 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_327
timestamp 1667941163
transform 1 0 31188 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_8
timestamp 1667941163
transform 1 0 1840 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_16
timestamp 1667941163
transform 1 0 2576 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_20
timestamp 1667941163
transform 1 0 2944 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_34
timestamp 1667941163
transform 1 0 4232 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_38
timestamp 1667941163
transform 1 0 4600 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_52
timestamp 1667941163
transform 1 0 5888 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_69
timestamp 1667941163
transform 1 0 7452 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_76
timestamp 1667941163
transform 1 0 8096 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_90
timestamp 1667941163
transform 1 0 9384 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_102
timestamp 1667941163
transform 1 0 10488 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_114
timestamp 1667941163
transform 1 0 11592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_138
timestamp 1667941163
transform 1 0 13800 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_145
timestamp 1667941163
transform 1 0 14444 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_149
timestamp 1667941163
transform 1 0 14812 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_156
timestamp 1667941163
transform 1 0 15456 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_181
timestamp 1667941163
transform 1 0 17756 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1667941163
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_203
timestamp 1667941163
transform 1 0 19780 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_207
timestamp 1667941163
transform 1 0 20148 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_211
timestamp 1667941163
transform 1 0 20516 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_215
timestamp 1667941163
transform 1 0 20884 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_228
timestamp 1667941163
transform 1 0 22080 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_258
timestamp 1667941163
transform 1 0 24840 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_273
timestamp 1667941163
transform 1 0 26220 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_280
timestamp 1667941163
transform 1 0 26864 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_295
timestamp 1667941163
transform 1 0 28244 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_302
timestamp 1667941163
transform 1 0 28888 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_384
timestamp 1667941163
transform 1 0 36432 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_392
timestamp 1667941163
transform 1 0 37168 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_397
timestamp 1667941163
transform 1 0 37628 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_16
timestamp 1667941163
transform 1 0 2576 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_23
timestamp 1667941163
transform 1 0 3220 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_30
timestamp 1667941163
transform 1 0 3864 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_37
timestamp 1667941163
transform 1 0 4508 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_44
timestamp 1667941163
transform 1 0 5152 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_64
timestamp 1667941163
transform 1 0 6992 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_76
timestamp 1667941163
transform 1 0 8096 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_93
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_97
timestamp 1667941163
transform 1 0 10028 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_101
timestamp 1667941163
transform 1 0 10396 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1667941163
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_124
timestamp 1667941163
transform 1 0 12512 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_131
timestamp 1667941163
transform 1 0 13156 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_138
timestamp 1667941163
transform 1 0 13800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_145
timestamp 1667941163
transform 1 0 14444 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_152
timestamp 1667941163
transform 1 0 15088 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_159
timestamp 1667941163
transform 1 0 15732 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_166
timestamp 1667941163
transform 1 0 16376 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_191
timestamp 1667941163
transform 1 0 18676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_197
timestamp 1667941163
transform 1 0 19228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_201
timestamp 1667941163
transform 1 0 19596 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_212
timestamp 1667941163
transform 1 0 20608 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_219
timestamp 1667941163
transform 1 0 21252 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_231
timestamp 1667941163
transform 1 0 22356 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_238
timestamp 1667941163
transform 1 0 23000 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_245
timestamp 1667941163
transform 1 0 23644 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_252
timestamp 1667941163
transform 1 0 24288 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_258
timestamp 1667941163
transform 1 0 24840 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_268
timestamp 1667941163
transform 1 0 25760 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_275
timestamp 1667941163
transform 1 0 26404 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1667941163
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_298
timestamp 1667941163
transform 1 0 28520 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_305
timestamp 1667941163
transform 1 0 29164 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_312
timestamp 1667941163
transform 1 0 29808 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_324
timestamp 1667941163
transform 1 0 30912 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_372
timestamp 1667941163
transform 1 0 35328 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_379
timestamp 1667941163
transform 1 0 35972 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_385
timestamp 1667941163
transform 1 0 36524 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1667941163
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_15
timestamp 1667941163
transform 1 0 2484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1667941163
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1667941163
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_34
timestamp 1667941163
transform 1 0 4232 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_41
timestamp 1667941163
transform 1 0 4876 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_49
timestamp 1667941163
transform 1 0 5612 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_54
timestamp 1667941163
transform 1 0 6072 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_62
timestamp 1667941163
transform 1 0 6808 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_74
timestamp 1667941163
transform 1 0 7912 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1667941163
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_93
timestamp 1667941163
transform 1 0 9660 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_98
timestamp 1667941163
transform 1 0 10120 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_106
timestamp 1667941163
transform 1 0 10856 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_110
timestamp 1667941163
transform 1 0 11224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_119
timestamp 1667941163
transform 1 0 12052 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_127
timestamp 1667941163
transform 1 0 12788 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_131
timestamp 1667941163
transform 1 0 13156 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1667941163
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_147
timestamp 1667941163
transform 1 0 14628 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_158
timestamp 1667941163
transform 1 0 15640 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_166
timestamp 1667941163
transform 1 0 16376 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_174
timestamp 1667941163
transform 1 0 17112 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_182
timestamp 1667941163
transform 1 0 17848 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_190
timestamp 1667941163
transform 1 0 18584 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_194
timestamp 1667941163
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_202
timestamp 1667941163
transform 1 0 19688 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_210
timestamp 1667941163
transform 1 0 20424 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_221
timestamp 1667941163
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_237
timestamp 1667941163
transform 1 0 22908 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1667941163
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1667941163
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_259
timestamp 1667941163
transform 1 0 24932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_266
timestamp 1667941163
transform 1 0 25576 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_273
timestamp 1667941163
transform 1 0 26220 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_279
timestamp 1667941163
transform 1 0 26772 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_286
timestamp 1667941163
transform 1 0 27416 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_294
timestamp 1667941163
transform 1 0 28152 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1667941163
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1667941163
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_314
timestamp 1667941163
transform 1 0 29992 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_321
timestamp 1667941163
transform 1 0 30636 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_328
timestamp 1667941163
transform 1 0 31280 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_343
timestamp 1667941163
transform 1 0 32660 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_350
timestamp 1667941163
transform 1 0 33304 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_362
timestamp 1667941163
transform 1 0 34408 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_377
timestamp 1667941163
transform 1 0 35788 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_385
timestamp 1667941163
transform 1 0 36524 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_391
timestamp 1667941163
transform 1 0 37076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1667941163
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0383_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22632 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0384_
timestamp 1667941163
transform 1 0 20884 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0385_
timestamp 1667941163
transform 1 0 23460 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0386_
timestamp 1667941163
transform 1 0 17296 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0387_
timestamp 1667941163
transform 1 0 21988 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0388_
timestamp 1667941163
transform 1 0 18492 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0389_
timestamp 1667941163
transform 1 0 15548 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0390_
timestamp 1667941163
transform 1 0 11592 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0391_
timestamp 1667941163
transform 1 0 14628 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0392_
timestamp 1667941163
transform 1 0 11684 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0393_
timestamp 1667941163
transform 1 0 18400 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0394_
timestamp 1667941163
transform 1 0 17480 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0395_
timestamp 1667941163
transform 1 0 25300 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0396_
timestamp 1667941163
transform 1 0 24840 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0397_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 26128 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0398_
timestamp 1667941163
transform 1 0 25576 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0399_
timestamp 1667941163
transform 1 0 9568 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0400_
timestamp 1667941163
transform 1 0 8372 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0401_
timestamp 1667941163
transform 1 0 12420 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0402_
timestamp 1667941163
transform 1 0 20516 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0403_
timestamp 1667941163
transform 1 0 23736 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0404_
timestamp 1667941163
transform 1 0 23184 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0405_
timestamp 1667941163
transform 1 0 3956 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0406_
timestamp 1667941163
transform 1 0 3588 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0407_
timestamp 1667941163
transform 1 0 30912 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0408_
timestamp 1667941163
transform 1 0 25668 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0409_
timestamp 1667941163
transform 1 0 26128 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0410_
timestamp 1667941163
transform 1 0 25760 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0411_
timestamp 1667941163
transform 1 0 30452 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0412_
timestamp 1667941163
transform 1 0 31556 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0413_
timestamp 1667941163
transform 1 0 23736 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0414_
timestamp 1667941163
transform 1 0 21988 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0415_
timestamp 1667941163
transform 1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0416_
timestamp 1667941163
transform 1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0417_
timestamp 1667941163
transform 1 0 25208 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0418_
timestamp 1667941163
transform 1 0 25208 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0419_
timestamp 1667941163
transform 1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0420_
timestamp 1667941163
transform 1 0 25024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0421_
timestamp 1667941163
transform 1 0 26496 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0422_
timestamp 1667941163
transform 1 0 24656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0423_
timestamp 1667941163
transform 1 0 20700 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0424_
timestamp 1667941163
transform 1 0 18676 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0425_
timestamp 1667941163
transform 1 0 18216 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0426_
timestamp 1667941163
transform 1 0 26036 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0427_
timestamp 1667941163
transform 1 0 27140 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0428_
timestamp 1667941163
transform 1 0 21988 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0429_
timestamp 1667941163
transform 1 0 23644 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0430_
timestamp 1667941163
transform 1 0 24564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0431_
timestamp 1667941163
transform 1 0 24564 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0432_
timestamp 1667941163
transform 1 0 20884 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0433_
timestamp 1667941163
transform 1 0 15916 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0434_
timestamp 1667941163
transform 1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0435_
timestamp 1667941163
transform 1 0 25300 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0436_
timestamp 1667941163
transform 1 0 26128 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0437_
timestamp 1667941163
transform 1 0 23000 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0438_
timestamp 1667941163
transform 1 0 25208 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0439_
timestamp 1667941163
transform 1 0 25576 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0440_
timestamp 1667941163
transform 1 0 21344 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0441_
timestamp 1667941163
transform 1 0 18676 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0442_
timestamp 1667941163
transform 1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0443_
timestamp 1667941163
transform 1 0 15364 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0444_
timestamp 1667941163
transform 1 0 23276 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0445_
timestamp 1667941163
transform 1 0 23920 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0446_
timestamp 1667941163
transform 1 0 27784 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0447_
timestamp 1667941163
transform 1 0 27324 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0448_
timestamp 1667941163
transform 1 0 28152 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0449_
timestamp 1667941163
transform 1 0 28612 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0450_
timestamp 1667941163
transform 1 0 29716 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0451_
timestamp 1667941163
transform 1 0 27784 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0452_
timestamp 1667941163
transform 1 0 28704 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0453_
timestamp 1667941163
transform 1 0 29716 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0454_
timestamp 1667941163
transform 1 0 29256 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0455_
timestamp 1667941163
transform 1 0 28888 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0456_
timestamp 1667941163
transform 1 0 29808 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0457_
timestamp 1667941163
transform 1 0 30452 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0458_
timestamp 1667941163
transform 1 0 13156 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0459_
timestamp 1667941163
transform 1 0 22356 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0460_
timestamp 1667941163
transform 1 0 22816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0461_
timestamp 1667941163
transform 1 0 23460 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0462_
timestamp 1667941163
transform 1 0 10948 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0463_
timestamp 1667941163
transform 1 0 11500 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0464_
timestamp 1667941163
transform 1 0 14168 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0465_
timestamp 1667941163
transform 1 0 13800 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0466_
timestamp 1667941163
transform 1 0 13156 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0467_
timestamp 1667941163
transform 1 0 29072 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0468_
timestamp 1667941163
transform 1 0 28980 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0469_
timestamp 1667941163
transform 1 0 29164 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0470_
timestamp 1667941163
transform 1 0 28796 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0471_
timestamp 1667941163
transform 1 0 28980 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0472_
timestamp 1667941163
transform 1 0 29716 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0473_
timestamp 1667941163
transform 1 0 27508 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0474_
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0475_
timestamp 1667941163
transform 1 0 28336 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0476_
timestamp 1667941163
transform 1 0 11960 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0477_
timestamp 1667941163
transform 1 0 6900 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1667941163
transform 1 0 1564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1667941163
transform 1 0 2300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0480_
timestamp 1667941163
transform 1 0 23184 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0481_
timestamp 1667941163
transform 1 0 13340 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0482_
timestamp 1667941163
transform 1 0 5520 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0483_
timestamp 1667941163
transform 1 0 2668 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1667941163
transform 1 0 17940 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1667941163
transform 1 0 14628 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0486_
timestamp 1667941163
transform 1 0 7176 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0487_
timestamp 1667941163
transform 1 0 22632 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0488_
timestamp 1667941163
transform 1 0 20976 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0489_
timestamp 1667941163
transform 1 0 22172 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1667941163
transform 1 0 14536 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1667941163
transform 1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0492_
timestamp 1667941163
transform 1 0 23920 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0493_
timestamp 1667941163
transform 1 0 18676 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0494_
timestamp 1667941163
transform 1 0 5612 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0495_
timestamp 1667941163
transform 1 0 7820 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1667941163
transform 1 0 24564 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1667941163
transform 1 0 22724 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0498_
timestamp 1667941163
transform 1 0 7636 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0499_
timestamp 1667941163
transform 1 0 18768 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0500_
timestamp 1667941163
transform 1 0 4968 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0501_
timestamp 1667941163
transform 1 0 16008 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502_
timestamp 1667941163
transform 1 0 3496 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1667941163
transform 1 0 16836 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0504_
timestamp 1667941163
transform 1 0 2484 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0505_
timestamp 1667941163
transform 1 0 6716 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0506_
timestamp 1667941163
transform 1 0 4600 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0507_
timestamp 1667941163
transform 1 0 28336 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0508_
timestamp 1667941163
transform 1 0 6532 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0509_
timestamp 1667941163
transform 1 0 29624 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0510_
timestamp 1667941163
transform 1 0 24564 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0511_
timestamp 1667941163
transform 1 0 28336 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0512_
timestamp 1667941163
transform 1 0 7176 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0513_
timestamp 1667941163
transform 1 0 24564 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1667941163
transform 1 0 25024 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0515_
timestamp 1667941163
transform 1 0 28704 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0516_
timestamp 1667941163
transform 1 0 24288 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0517_
timestamp 1667941163
transform 1 0 25668 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0518_
timestamp 1667941163
transform 1 0 25208 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0519_
timestamp 1667941163
transform 1 0 28336 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp 1667941163
transform 1 0 23368 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0521_
timestamp 1667941163
transform 1 0 24932 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0522_
timestamp 1667941163
transform 1 0 23552 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0523_
timestamp 1667941163
transform 1 0 21988 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0524_
timestamp 1667941163
transform 1 0 20608 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0525_
timestamp 1667941163
transform 1 0 16836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0526_
timestamp 1667941163
transform 1 0 20424 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0527_
timestamp 1667941163
transform 1 0 21988 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0528_
timestamp 1667941163
transform 1 0 19596 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1667941163
transform 1 0 23368 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0530_
timestamp 1667941163
transform 1 0 6532 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0531_
timestamp 1667941163
transform 1 0 20700 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1667941163
transform 1 0 24196 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1667941163
transform 1 0 22632 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0534_
timestamp 1667941163
transform 1 0 28612 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0535_
timestamp 1667941163
transform 1 0 22908 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0536_
timestamp 1667941163
transform 1 0 23920 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0537_
timestamp 1667941163
transform 1 0 12880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1667941163
transform 1 0 27140 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0539_
timestamp 1667941163
transform 1 0 28612 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0540_
timestamp 1667941163
transform 1 0 4048 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0541_
timestamp 1667941163
transform 1 0 8096 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0542_
timestamp 1667941163
transform 1 0 9200 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0543_
timestamp 1667941163
transform 1 0 17756 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0544_
timestamp 1667941163
transform 1 0 5520 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0545_
timestamp 1667941163
transform 1 0 3036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0546_
timestamp 1667941163
transform 1 0 2024 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1667941163
transform 1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0548_
timestamp 1667941163
transform 1 0 23092 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0549_
timestamp 1667941163
transform 1 0 2944 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1667941163
transform 1 0 25484 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0551_
timestamp 1667941163
transform 1 0 3956 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0552_
timestamp 1667941163
transform 1 0 23552 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0553_
timestamp 1667941163
transform 1 0 18768 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0554_
timestamp 1667941163
transform 1 0 27232 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0555_
timestamp 1667941163
transform 1 0 18308 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1667941163
transform 1 0 26404 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0557_
timestamp 1667941163
transform 1 0 21988 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0558_
timestamp 1667941163
transform 1 0 10120 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0559_
timestamp 1667941163
transform 1 0 23276 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0560_
timestamp 1667941163
transform 1 0 20332 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0561_
timestamp 1667941163
transform 1 0 30268 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0562_
timestamp 1667941163
transform 1 0 26404 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0563_
timestamp 1667941163
transform 1 0 25208 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0564_
timestamp 1667941163
transform 1 0 17480 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1667941163
transform 1 0 23276 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0566_
timestamp 1667941163
transform 1 0 24564 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0567_
timestamp 1667941163
transform 1 0 15180 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0568_
timestamp 1667941163
transform 1 0 23368 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0569_
timestamp 1667941163
transform 1 0 12420 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0570_
timestamp 1667941163
transform 1 0 9936 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1667941163
transform 1 0 15456 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0572_
timestamp 1667941163
transform 1 0 22264 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0573_
timestamp 1667941163
transform 1 0 24104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0574_
timestamp 1667941163
transform 1 0 11776 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0575_
timestamp 1667941163
transform 1 0 23460 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0576_
timestamp 1667941163
transform 1 0 10672 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 1667941163
transform 1 0 27140 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0578_
timestamp 1667941163
transform 1 0 24564 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0579_
timestamp 1667941163
transform 1 0 21344 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0580_
timestamp 1667941163
transform 1 0 2484 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0581_
timestamp 1667941163
transform 1 0 9292 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0582_
timestamp 1667941163
transform 1 0 6532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1667941163
transform 1 0 9752 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0584_
timestamp 1667941163
transform 1 0 23828 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0585_
timestamp 1667941163
transform 1 0 23828 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0586_
timestamp 1667941163
transform 1 0 3956 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0587_
timestamp 1667941163
transform 1 0 4324 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1667941163
transform 1 0 13064 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0589_
timestamp 1667941163
transform 1 0 22724 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0590_
timestamp 1667941163
transform 1 0 22080 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1667941163
transform 1 0 27876 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0592_
timestamp 1667941163
transform 1 0 26496 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0593_
timestamp 1667941163
transform 1 0 5612 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0594_
timestamp 1667941163
transform 1 0 14076 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0595_
timestamp 1667941163
transform 1 0 16836 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1667941163
transform 1 0 21160 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0597_
timestamp 1667941163
transform 1 0 23920 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0598_
timestamp 1667941163
transform 1 0 27784 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0599_
timestamp 1667941163
transform 1 0 25576 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0600_
timestamp 1667941163
transform 1 0 13524 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1667941163
transform 1 0 23552 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0602_
timestamp 1667941163
transform 1 0 23736 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0603_
timestamp 1667941163
transform 1 0 25208 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0604_
timestamp 1667941163
transform 1 0 21068 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0605_
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0606_
timestamp 1667941163
transform 1 0 17848 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1667941163
transform 1 0 22540 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0608_
timestamp 1667941163
transform 1 0 25300 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 1667941163
transform 1 0 23092 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1667941163
transform 1 0 22080 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0611_
timestamp 1667941163
transform 1 0 34224 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0612_
timestamp 1667941163
transform 1 0 13524 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0613_
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 1667941163
transform 1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0615_
timestamp 1667941163
transform 1 0 27324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1667941163
transform 1 0 21988 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0617_
timestamp 1667941163
transform 1 0 14628 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0618_
timestamp 1667941163
transform 1 0 3680 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1667941163
transform 1 0 28980 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 1667941163
transform 1 0 20516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 1667941163
transform 1 0 24380 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1667941163
transform 1 0 6532 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 1667941163
transform 1 0 29808 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0624_
timestamp 1667941163
transform 1 0 10948 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1667941163
transform 1 0 29072 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 1667941163
transform 1 0 18584 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 1667941163
transform 1 0 27416 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1667941163
transform 1 0 23920 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 1667941163
transform 1 0 18584 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0630_
timestamp 1667941163
transform 1 0 35052 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1667941163
transform 1 0 30728 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1667941163
transform 1 0 27048 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1667941163
transform 1 0 22448 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 1667941163
transform 1 0 19412 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0635_
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0636_
timestamp 1667941163
transform 1 0 22908 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1667941163
transform 1 0 28244 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1667941163
transform 1 0 13984 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0639_
timestamp 1667941163
transform 1 0 2300 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1667941163
transform 1 0 1840 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0642_
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1667941163
transform 1 0 3128 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0644_
timestamp 1667941163
transform 1 0 27140 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1667941163
transform 1 0 19780 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1667941163
transform 1 0 17756 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1667941163
transform 1 0 10488 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0648_
timestamp 1667941163
transform 1 0 7452 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0649_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1840 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1667941163
transform 1 0 35972 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0651_
timestamp 1667941163
transform 1 0 12236 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1667941163
transform 1 0 13892 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0653_
timestamp 1667941163
transform 1 0 29532 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0654_
timestamp 1667941163
transform 1 0 27324 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1667941163
transform 1 0 2852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1667941163
transform 1 0 18676 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1667941163
transform 1 0 20792 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 1667941163
transform 1 0 24564 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1667941163
transform 1 0 31188 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0660_
timestamp 1667941163
transform 1 0 26404 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1667941163
transform 1 0 5520 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0662_
timestamp 1667941163
transform 1 0 26404 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0663_
timestamp 1667941163
transform 1 0 2208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1667941163
transform 1 0 28980 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1667941163
transform 1 0 2944 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0666_
timestamp 1667941163
transform 1 0 3956 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1667941163
transform 1 0 7084 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1667941163
transform 1 0 24564 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 1667941163
transform 1 0 21160 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0671_
timestamp 1667941163
transform 1 0 4232 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1667941163
transform 1 0 21988 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1667941163
transform 1 0 14168 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1667941163
transform 1 0 2944 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1667941163
transform 1 0 30176 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1667941163
transform 1 0 26404 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1667941163
transform 1 0 29716 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0678_
timestamp 1667941163
transform 1 0 2300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1667941163
transform 1 0 3220 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0680_
timestamp 1667941163
transform 1 0 31832 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1667941163
transform 1 0 27140 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1667941163
transform 1 0 4600 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1667941163
transform 1 0 10212 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1667941163
transform 1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1667941163
transform 1 0 19872 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1667941163
transform 1 0 30728 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1667941163
transform 1 0 28888 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1667941163
transform 1 0 25208 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1667941163
transform 1 0 29624 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1667941163
transform 1 0 31372 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1667941163
transform 1 0 21988 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1667941163
transform 1 0 30820 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1667941163
transform 1 0 5796 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1667941163
transform 1 0 17572 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1667941163
transform 1 0 29900 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1667941163
transform 1 0 4968 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1667941163
transform 1 0 27600 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1667941163
transform 1 0 32568 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1667941163
transform 1 0 25576 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0700_
timestamp 1667941163
transform 1 0 1840 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1667941163
transform 1 0 26312 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1667941163
transform 1 0 5796 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1667941163
transform 1 0 23276 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform 1 0 6532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1667941163
transform 1 0 11776 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1667941163
transform 1 0 23460 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0707_
timestamp 1667941163
transform 1 0 12328 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1667941163
transform 1 0 24564 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 1667941163
transform 1 0 27140 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1667941163
transform 1 0 29992 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1667941163
transform 1 0 14260 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0712_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27324 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0713_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 18400 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0714_
timestamp 1667941163
transform 1 0 20056 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1667941163
transform 1 0 20056 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1667941163
transform 1 0 19872 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1667941163
transform 1 0 18676 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1667941163
transform 1 0 18676 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1667941163
transform 1 0 20700 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1667941163
transform 1 0 14536 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1667941163
transform 1 0 19872 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1667941163
transform 1 0 4416 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1667941163
transform 1 0 5152 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0725_
timestamp 1667941163
transform 1 0 21988 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1667941163
transform 1 0 5796 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1667941163
transform 1 0 6624 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1667941163
transform 1 0 21160 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1667941163
transform 1 0 20240 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1667941163
transform 1 0 20148 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1667941163
transform 1 0 20056 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1667941163
transform 1 0 5336 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1667941163
transform 1 0 5520 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1667941163
transform 1 0 8096 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1667941163
transform 1 0 19872 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0736_
timestamp 1667941163
transform 1 0 20332 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1667941163
transform 1 0 21988 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1667941163
transform 1 0 3220 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1667941163
transform 1 0 7728 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1667941163
transform 1 0 22632 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1667941163
transform 1 0 5336 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1667941163
transform 1 0 4692 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1667941163
transform 1 0 8740 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1667941163
transform 1 0 21160 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1667941163
transform 1 0 20608 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1667941163
transform 1 0 12144 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0747_
timestamp 1667941163
transform 1 0 18768 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1667941163
transform 1 0 21252 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform 1 0 20976 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1667941163
transform 1 0 20516 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1667941163
transform 1 0 21160 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1667941163
transform 1 0 21804 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1667941163
transform 1 0 19780 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1667941163
transform 1 0 19412 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1667941163
transform 1 0 20056 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1667941163
transform 1 0 21068 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1667941163
transform 1 0 19412 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0758_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19872 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1667941163
transform 1 0 3404 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1667941163
transform 1 0 2300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1667941163
transform 1 0 5060 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1667941163
transform 1 0 1840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1667941163
transform 1 0 18676 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1667941163
transform 1 0 21252 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1667941163
transform 1 0 20792 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1667941163
transform 1 0 19228 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1667941163
transform 1 0 18676 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1667941163
transform 1 0 19136 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0769_
timestamp 1667941163
transform 1 0 19412 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1667941163
transform 1 0 20332 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1667941163
transform 1 0 20608 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1667941163
transform 1 0 19412 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1667941163
transform 1 0 23368 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1667941163
transform 1 0 20884 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1667941163
transform 1 0 16100 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1667941163
transform 1 0 15456 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1667941163
transform 1 0 20976 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0780_
timestamp 1667941163
transform 1 0 19412 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1667941163
transform 1 0 19504 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1667941163
transform 1 0 19412 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1667941163
transform 1 0 11684 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1667941163
transform 1 0 8372 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1667941163
transform 1 0 22172 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1667941163
transform 1 0 17940 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1667941163
transform 1 0 17296 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1667941163
transform 1 0 18032 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1667941163
transform 1 0 7636 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0791_
timestamp 1667941163
transform 1 0 19412 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1667941163
transform 1 0 7360 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1667941163
transform 1 0 6716 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1667941163
transform 1 0 9108 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1667941163
transform 1 0 9108 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1667941163
transform 1 0 14812 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1667941163
transform 1 0 19228 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1667941163
transform 1 0 19872 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1667941163
transform 1 0 15364 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1667941163
transform 1 0 18584 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0802_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21988 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1667941163
transform 1 0 20516 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1667941163
transform 1 0 13064 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1667941163
transform 1 0 2852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0806_
timestamp 1667941163
transform 1 0 4048 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 3956 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1667941163
transform 1 0 21068 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1667941163
transform 1 0 16836 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1667941163
transform 1 0 2760 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1667941163
transform 1 0 3220 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0813_
timestamp 1667941163
transform 1 0 18952 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1667941163
transform 1 0 8096 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1667941163
transform 1 0 18676 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1667941163
transform 1 0 19688 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1667941163
transform 1 0 19320 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1667941163
transform 1 0 10212 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1667941163
transform 1 0 20240 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1667941163
transform 1 0 19504 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1667941163
transform 1 0 18676 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1667941163
transform 1 0 14260 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1667941163
transform 1 0 19412 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0824_
timestamp 1667941163
transform 1 0 18492 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1667941163
transform 1 0 23552 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1667941163
transform 1 0 15364 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1667941163
transform 1 0 17020 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1667941163
transform 1 0 20056 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1667941163
transform 1 0 16652 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1667941163
transform 1 0 21528 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1667941163
transform 1 0 19228 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1667941163
transform 1 0 14444 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1667941163
transform 1 0 19780 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1667941163
transform 1 0 21620 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1667941163
transform 1 0 19780 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1667941163
transform 1 0 20424 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1667941163
transform 1 0 18676 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1667941163
transform 1 0 20884 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1667941163
transform 1 0 10304 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1667941163
transform 1 0 10856 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1667941163
transform 1 0 11500 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1667941163
transform 1 0 19504 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _0843_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12788 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0844_
timestamp 1667941163
transform 1 0 16008 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0845_
timestamp 1667941163
transform 1 0 16836 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0846_
timestamp 1667941163
transform 1 0 15824 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0847_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11868 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0848_
timestamp 1667941163
transform 1 0 15824 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0849_
timestamp 1667941163
transform 1 0 10396 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0850_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3956 0 1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0851_
timestamp 1667941163
transform 1 0 4232 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0852_
timestamp 1667941163
transform 1 0 5060 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0853_
timestamp 1667941163
transform 1 0 6532 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0854_
timestamp 1667941163
transform 1 0 5704 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0855_
timestamp 1667941163
transform 1 0 14444 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0856_
timestamp 1667941163
transform 1 0 15364 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0857_
timestamp 1667941163
transform 1 0 15916 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0858_
timestamp 1667941163
transform 1 0 16836 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0859_
timestamp 1667941163
transform 1 0 5888 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0860_
timestamp 1667941163
transform 1 0 1656 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0861_
timestamp 1667941163
transform 1 0 6716 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0862_
timestamp 1667941163
transform 1 0 7636 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0863_
timestamp 1667941163
transform 1 0 7544 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0864_
timestamp 1667941163
transform 1 0 2576 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0865_
timestamp 1667941163
transform 1 0 7912 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0866_
timestamp 1667941163
transform 1 0 8372 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0867_
timestamp 1667941163
transform 1 0 9384 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0868_
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0869_
timestamp 1667941163
transform 1 0 9108 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0870_
timestamp 1667941163
transform 1 0 11960 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0871_
timestamp 1667941163
transform 1 0 10488 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0872_
timestamp 1667941163
transform 1 0 11224 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0873_
timestamp 1667941163
transform 1 0 14076 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0874_
timestamp 1667941163
transform 1 0 14904 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0875_
timestamp 1667941163
transform 1 0 9384 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0876_
timestamp 1667941163
transform 1 0 6716 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0877_
timestamp 1667941163
transform 1 0 16836 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0878_
timestamp 1667941163
transform 1 0 14444 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0879_
timestamp 1667941163
transform 1 0 15824 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0880_
timestamp 1667941163
transform 1 0 11592 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0881_
timestamp 1667941163
transform 1 0 9292 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0882_
timestamp 1667941163
transform 1 0 9292 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0883_
timestamp 1667941163
transform 1 0 1656 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0884_
timestamp 1667941163
transform 1 0 1656 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0885_
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0886_
timestamp 1667941163
transform 1 0 3220 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0887_
timestamp 1667941163
transform 1 0 6716 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0888_
timestamp 1667941163
transform 1 0 2392 0 -1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0889_
timestamp 1667941163
transform 1 0 3036 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0890_
timestamp 1667941163
transform 1 0 11684 0 1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0891_
timestamp 1667941163
transform 1 0 15824 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0892_
timestamp 1667941163
transform 1 0 16836 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0893_
timestamp 1667941163
transform 1 0 14444 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0894_
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0895_
timestamp 1667941163
transform 1 0 4600 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0896_
timestamp 1667941163
transform 1 0 15272 0 1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0897_
timestamp 1667941163
transform 1 0 12696 0 -1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0898_
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0899_
timestamp 1667941163
transform 1 0 16836 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0900_
timestamp 1667941163
transform 1 0 16836 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0901_
timestamp 1667941163
transform 1 0 14536 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0902_
timestamp 1667941163
transform 1 0 11684 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0903_
timestamp 1667941163
transform 1 0 9108 0 1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0904_
timestamp 1667941163
transform 1 0 10304 0 1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0905_
timestamp 1667941163
transform 1 0 4232 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0906_
timestamp 1667941163
transform 1 0 4232 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0907_
timestamp 1667941163
transform 1 0 3956 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0908_
timestamp 1667941163
transform 1 0 10948 0 1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0909_
timestamp 1667941163
transform 1 0 9108 0 -1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0910_
timestamp 1667941163
transform 1 0 11684 0 1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0911_
timestamp 1667941163
transform 1 0 1564 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0912_
timestamp 1667941163
transform 1 0 1564 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0913_
timestamp 1667941163
transform 1 0 2668 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0914_
timestamp 1667941163
transform 1 0 1564 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0915_
timestamp 1667941163
transform 1 0 5060 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0916_
timestamp 1667941163
transform 1 0 6440 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0917_
timestamp 1667941163
transform 1 0 9384 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0918_
timestamp 1667941163
transform 1 0 5612 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0919_
timestamp 1667941163
transform 1 0 4232 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0920_
timestamp 1667941163
transform 1 0 2024 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0921_
timestamp 1667941163
transform 1 0 3220 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0922_
timestamp 1667941163
transform 1 0 9108 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0923_
timestamp 1667941163
transform 1 0 9292 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0924_
timestamp 1667941163
transform 1 0 5244 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0925_
timestamp 1667941163
transform 1 0 6808 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0926_
timestamp 1667941163
transform 1 0 8188 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0927_
timestamp 1667941163
transform 1 0 9568 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0928_
timestamp 1667941163
transform 1 0 6072 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0929_
timestamp 1667941163
transform 1 0 11684 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0930_
timestamp 1667941163
transform 1 0 7176 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0931_
timestamp 1667941163
transform 1 0 1564 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0932_
timestamp 1667941163
transform 1 0 4416 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0933_
timestamp 1667941163
transform 1 0 4232 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0934_
timestamp 1667941163
transform 1 0 6348 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0935_
timestamp 1667941163
transform 1 0 11776 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0936_
timestamp 1667941163
transform 1 0 15732 0 1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0937_
timestamp 1667941163
transform 1 0 9108 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0938_
timestamp 1667941163
transform 1 0 15456 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0939_
timestamp 1667941163
transform 1 0 11960 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0940_
timestamp 1667941163
transform 1 0 11684 0 -1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0941_
timestamp 1667941163
transform 1 0 11960 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0942_
timestamp 1667941163
transform -1 0 15916 0 -1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0943_
timestamp 1667941163
transform 1 0 15088 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0944_
timestamp 1667941163
transform 1 0 12880 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0945_
timestamp 1667941163
transform 1 0 14536 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0946_
timestamp 1667941163
transform 1 0 15088 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0947_
timestamp 1667941163
transform 1 0 16836 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0948_
timestamp 1667941163
transform 1 0 15364 0 1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0949_
timestamp 1667941163
transform 1 0 9292 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0950_
timestamp 1667941163
transform 1 0 11592 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0951_
timestamp 1667941163
transform 1 0 5244 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0952_
timestamp 1667941163
transform 1 0 9292 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0953_
timestamp 1667941163
transform 1 0 6900 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0954_
timestamp 1667941163
transform 1 0 1564 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0955_
timestamp 1667941163
transform 1 0 16008 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0956_
timestamp 1667941163
transform 1 0 11684 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0957_
timestamp 1667941163
transform 1 0 9108 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0958_
timestamp 1667941163
transform 1 0 11868 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0959_
timestamp 1667941163
transform 1 0 13248 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0960_
timestamp 1667941163
transform 1 0 15732 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_1  _0985_
timestamp 1667941163
transform 1 0 28796 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0986_
timestamp 1667941163
transform 1 0 36156 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0987_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15640 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0988_
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0989_
timestamp 1667941163
transform 1 0 12972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0990_
timestamp 1667941163
transform 1 0 32568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0991_
timestamp 1667941163
transform 1 0 31464 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0992_
timestamp 1667941163
transform 1 0 32292 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0993_
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1667941163
transform 1 0 34868 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0995_
timestamp 1667941163
transform 1 0 2668 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0996_
timestamp 1667941163
transform 1 0 2300 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0997_
timestamp 1667941163
transform 1 0 33120 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1667941163
transform 1 0 6624 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0999_
timestamp 1667941163
transform 1 0 34132 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1667941163
transform 1 0 25300 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1001_
timestamp 1667941163
transform 1 0 31096 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1002_
timestamp 1667941163
transform 1 0 22724 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 1667941163
transform 1 0 3956 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1667941163
transform 1 0 21160 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1005_
timestamp 1667941163
transform 1 0 17020 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1667941163
transform 1 0 6532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1667941163
transform 1 0 22632 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1008_
timestamp 1667941163
transform 1 0 19688 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1667941163
transform 1 0 26128 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1667941163
transform 1 0 36248 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1011_
timestamp 1667941163
transform 1 0 22724 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1012_
timestamp 1667941163
transform 1 0 13432 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1013_
timestamp 1667941163
transform 1 0 28520 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1014_
timestamp 1667941163
transform 1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1667941163
transform 1 0 35144 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1667941163
transform 1 0 37812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1017_
timestamp 1667941163
transform 1 0 24840 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1667941163
transform 1 0 35696 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1019_
timestamp 1667941163
transform 1 0 31740 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1020_
timestamp 1667941163
transform 1 0 15640 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1021_
timestamp 1667941163
transform 1 0 25116 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1667941163
transform 1 0 21712 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1023_
timestamp 1667941163
transform 1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 1667941163
transform 1 0 20332 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1667941163
transform 1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1667941163
transform 1 0 7912 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1027_
timestamp 1667941163
transform 1 0 30084 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1028_
timestamp 1667941163
transform 1 0 23644 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1667941163
transform 1 0 35052 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1030_
timestamp 1667941163
transform 1 0 24196 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1667941163
transform 1 0 36616 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1032_
timestamp 1667941163
transform 1 0 27140 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1667941163
transform 1 0 16376 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1667941163
transform 1 0 20056 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1035_
timestamp 1667941163
transform 1 0 1748 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1036_
timestamp 1667941163
transform 1 0 9292 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1037_
timestamp 1667941163
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1038_
timestamp 1667941163
transform 1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1039_
timestamp 1667941163
transform 1 0 24656 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1040_
timestamp 1667941163
transform 1 0 20976 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1667941163
transform 1 0 34224 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1042_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27416 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1043_
timestamp 1667941163
transform 1 0 26220 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1044_
timestamp 1667941163
transform 1 0 32476 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1044__142 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 32660 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1045_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1046_
timestamp 1667941163
transform 1 0 19596 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1047_
timestamp 1667941163
transform 1 0 19412 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1048_
timestamp 1667941163
transform 1 0 27140 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1049_
timestamp 1667941163
transform 1 0 19504 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1050_
timestamp 1667941163
transform 1 0 27140 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1051_
timestamp 1667941163
transform 1 0 27140 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1052_
timestamp 1667941163
transform 1 0 12604 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1053_
timestamp 1667941163
transform 1 0 27140 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1054_
timestamp 1667941163
transform 1 0 20424 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1055_
timestamp 1667941163
transform 1 0 22172 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1056__143
timestamp 1667941163
transform 1 0 3036 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1056_
timestamp 1667941163
transform 1 0 2852 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1057_
timestamp 1667941163
transform 1 0 25760 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1058_
timestamp 1667941163
transform 1 0 27232 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1059_
timestamp 1667941163
transform 1 0 25484 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1060_
timestamp 1667941163
transform 1 0 25760 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1061_
timestamp 1667941163
transform 1 0 25760 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1062_
timestamp 1667941163
transform 1 0 20424 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1063_
timestamp 1667941163
transform 1 0 17112 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1064_
timestamp 1667941163
transform 1 0 20332 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1065_
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1066_
timestamp 1667941163
transform 1 0 9844 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1067_
timestamp 1667941163
transform 1 0 14260 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1068__144
timestamp 1667941163
transform 1 0 10672 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1068_
timestamp 1667941163
transform 1 0 10580 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1069_
timestamp 1667941163
transform 1 0 4692 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1070_
timestamp 1667941163
transform 1 0 3496 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1071_
timestamp 1667941163
transform 1 0 21160 0 1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1072_
timestamp 1667941163
transform 1 0 3956 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1073_
timestamp 1667941163
transform 1 0 24564 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1074_
timestamp 1667941163
transform 1 0 24748 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1075_
timestamp 1667941163
transform 1 0 11684 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1076_
timestamp 1667941163
transform 1 0 24564 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1077_
timestamp 1667941163
transform 1 0 27600 0 1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1078_
timestamp 1667941163
transform 1 0 14628 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1079_
timestamp 1667941163
transform 1 0 17572 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1080__145
timestamp 1667941163
transform 1 0 16192 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1080_
timestamp 1667941163
transform 1 0 14628 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1081_
timestamp 1667941163
transform 1 0 23644 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1082_
timestamp 1667941163
transform 1 0 8556 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1083_
timestamp 1667941163
transform 1 0 23368 0 -1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1084_
timestamp 1667941163
transform 1 0 23552 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1085_
timestamp 1667941163
transform 1 0 18952 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1086_
timestamp 1667941163
transform 1 0 23276 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1087_
timestamp 1667941163
transform 1 0 18124 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1088_
timestamp 1667941163
transform 1 0 21528 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1089_
timestamp 1667941163
transform 1 0 20700 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1090_
timestamp 1667941163
transform 1 0 25944 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1091_
timestamp 1667941163
transform 1 0 22448 0 1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1092__146
timestamp 1667941163
transform 1 0 28336 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1092_
timestamp 1667941163
transform 1 0 28060 0 1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1093_
timestamp 1667941163
transform 1 0 22908 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1094_
timestamp 1667941163
transform 1 0 25852 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1095_
timestamp 1667941163
transform 1 0 30176 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1096_
timestamp 1667941163
transform 1 0 27140 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1097_
timestamp 1667941163
transform 1 0 19688 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1098_
timestamp 1667941163
transform 1 0 27324 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1099_
timestamp 1667941163
transform 1 0 21988 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1100_
timestamp 1667941163
transform 1 0 19872 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1101_
timestamp 1667941163
transform 1 0 16192 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1102_
timestamp 1667941163
transform 1 0 1656 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1103_
timestamp 1667941163
transform 1 0 2024 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1104__147
timestamp 1667941163
transform 1 0 3680 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1104_
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1105_
timestamp 1667941163
transform 1 0 2024 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1106_
timestamp 1667941163
transform 1 0 25484 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1107_
timestamp 1667941163
transform 1 0 2024 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1108_
timestamp 1667941163
transform 1 0 10396 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1109_
timestamp 1667941163
transform 1 0 17572 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1110_
timestamp 1667941163
transform 1 0 14444 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1111_
timestamp 1667941163
transform 1 0 1748 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1112_
timestamp 1667941163
transform 1 0 26128 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1113_
timestamp 1667941163
transform 1 0 9016 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1114_
timestamp 1667941163
transform 1 0 23736 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1115_
timestamp 1667941163
transform 1 0 31832 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1116__148
timestamp 1667941163
transform 1 0 29348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1116_
timestamp 1667941163
transform 1 0 29716 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1117_
timestamp 1667941163
transform 1 0 27416 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1118_
timestamp 1667941163
transform 1 0 24932 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1119_
timestamp 1667941163
transform 1 0 25208 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1120_
timestamp 1667941163
transform 1 0 19596 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1121_
timestamp 1667941163
transform 1 0 16836 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1122_
timestamp 1667941163
transform 1 0 6532 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1123_
timestamp 1667941163
transform 1 0 17940 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1124_
timestamp 1667941163
transform 1 0 22724 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1125_
timestamp 1667941163
transform 1 0 19412 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1126_
timestamp 1667941163
transform 1 0 19412 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1127_
timestamp 1667941163
transform 1 0 22908 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1128_
timestamp 1667941163
transform 1 0 19688 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1129_
timestamp 1667941163
transform 1 0 18032 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1129__149
timestamp 1667941163
transform 1 0 18216 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1130_
timestamp 1667941163
transform 1 0 19320 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1131_
timestamp 1667941163
transform 1 0 19780 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1132_
timestamp 1667941163
transform 1 0 27140 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1133_
timestamp 1667941163
transform 1 0 22632 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1134_
timestamp 1667941163
transform 1 0 24564 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1135_
timestamp 1667941163
transform 1 0 23644 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1136_
timestamp 1667941163
transform 1 0 16928 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1137_
timestamp 1667941163
transform 1 0 26220 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1138_
timestamp 1667941163
transform -1 0 9292 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1139_
timestamp 1667941163
transform 1 0 9108 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1140_
timestamp 1667941163
transform 1 0 26036 0 1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1141__150
timestamp 1667941163
transform 1 0 20148 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1141_
timestamp 1667941163
transform 1 0 20332 0 -1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1142_
timestamp 1667941163
transform 1 0 27324 0 -1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1143_
timestamp 1667941163
transform 1 0 22356 0 -1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1144_
timestamp 1667941163
transform 1 0 27600 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1145_
timestamp 1667941163
transform 1 0 2852 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1146_
timestamp 1667941163
transform -1 0 2484 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1147_
timestamp 1667941163
transform 1 0 24840 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1148_
timestamp 1667941163
transform 1 0 21712 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1149_
timestamp 1667941163
transform 1 0 6256 0 1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1150_
timestamp 1667941163
transform 1 0 15916 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1151_
timestamp 1667941163
transform 1 0 2208 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1151__151
timestamp 1667941163
transform 1 0 2852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1152_
timestamp 1667941163
transform 1 0 20424 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1153_
timestamp 1667941163
transform 1 0 6532 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1154_
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1155_
timestamp 1667941163
transform 1 0 19412 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1156_
timestamp 1667941163
transform 1 0 20700 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1157__152
timestamp 1667941163
transform 1 0 25944 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1157_
timestamp 1667941163
transform 1 0 25392 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1158_
timestamp 1667941163
transform 1 0 8464 0 -1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1159_
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1160_
timestamp 1667941163
transform 1 0 21252 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1161_
timestamp 1667941163
transform 1 0 17940 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1162_
timestamp 1667941163
transform 1 0 25760 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1163_
timestamp 1667941163
transform 1 0 21988 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1164__153
timestamp 1667941163
transform 1 0 17020 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1164_
timestamp 1667941163
transform 1 0 17664 0 -1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1165_
timestamp 1667941163
transform 1 0 22356 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1166_
timestamp 1667941163
transform 1 0 7820 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1167_
timestamp 1667941163
transform 1 0 13708 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1168_
timestamp 1667941163
transform 1 0 18032 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1169_
timestamp 1667941163
transform 1 0 14260 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1170_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2944 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1171_
timestamp 1667941163
transform 1 0 11776 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1172_
timestamp 1667941163
transform 1 0 20976 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1172__154
timestamp 1667941163
transform 1 0 21252 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1173_
timestamp 1667941163
transform 1 0 1564 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1174_
timestamp 1667941163
transform 1 0 2024 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1175_
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1176_
timestamp 1667941163
transform 1 0 11776 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1177_
timestamp 1667941163
transform 1 0 6992 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1178_
timestamp 1667941163
transform 1 0 29900 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1179__155
timestamp 1667941163
transform 1 0 28980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1179_
timestamp 1667941163
transform 1 0 28428 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1180_
timestamp 1667941163
transform 1 0 28244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1181_
timestamp 1667941163
transform 1 0 31004 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1182_
timestamp 1667941163
transform 1 0 24932 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1183_
timestamp 1667941163
transform 1 0 29716 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1184_
timestamp 1667941163
transform 1 0 11868 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1185__156
timestamp 1667941163
transform 1 0 12972 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1185_
timestamp 1667941163
transform 1 0 12880 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1186_
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1187_
timestamp 1667941163
transform 1 0 12052 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1188_
timestamp 1667941163
transform 1 0 14260 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1189_
timestamp 1667941163
transform 1 0 23000 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1190_
timestamp 1667941163
transform 1 0 27876 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1191__157
timestamp 1667941163
transform 1 0 28152 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1191_
timestamp 1667941163
transform 1 0 27416 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1192_
timestamp 1667941163
transform 1 0 28152 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1193_
timestamp 1667941163
transform 1 0 27968 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1194_
timestamp 1667941163
transform 1 0 27784 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1195_
timestamp 1667941163
transform 1 0 27784 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1196_
timestamp 1667941163
transform 1 0 24564 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1197_
timestamp 1667941163
transform 1 0 28152 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1197__158
timestamp 1667941163
transform 1 0 28152 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1198_
timestamp 1667941163
transform 1 0 15272 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1199_
timestamp 1667941163
transform 1 0 20516 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1200_
timestamp 1667941163
transform 1 0 27876 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1201_
timestamp 1667941163
transform 1 0 19412 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1202_
timestamp 1667941163
transform 1 0 27140 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1203_
timestamp 1667941163
transform 1 0 25944 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1203__159
timestamp 1667941163
transform 1 0 25300 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1204_
timestamp 1667941163
transform 1 0 14444 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1205_
timestamp 1667941163
transform 1 0 23276 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1206_
timestamp 1667941163
transform 1 0 22356 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1207_
timestamp 1667941163
transform 1 0 20056 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1208_
timestamp 1667941163
transform 1 0 26404 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1209__160
timestamp 1667941163
transform 1 0 25576 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1209_
timestamp 1667941163
transform 1 0 25760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1210_
timestamp 1667941163
transform 1 0 17572 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1211_
timestamp 1667941163
transform 1 0 24564 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1212_
timestamp 1667941163
transform 1 0 21988 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1213_
timestamp 1667941163
transform 1 0 19412 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1214_
timestamp 1667941163
transform 1 0 25852 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1215_
timestamp 1667941163
transform 1 0 25668 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1215__161
timestamp 1667941163
transform 1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1216_
timestamp 1667941163
transform 1 0 18124 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1217_
timestamp 1667941163
transform 1 0 22540 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1218_
timestamp 1667941163
transform 1 0 27140 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1219_
timestamp 1667941163
transform 1 0 21988 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1220_
timestamp 1667941163
transform 1 0 31096 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1220__162
timestamp 1667941163
transform 1 0 31280 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1221_
timestamp 1667941163
transform 1 0 25944 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1222_
timestamp 1667941163
transform 1 0 29808 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1223_
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1224__163
timestamp 1667941163
transform 1 0 4876 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1224_
timestamp 1667941163
transform 1 0 4692 0 1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _1225_
timestamp 1667941163
transform 1 0 21988 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1226_
timestamp 1667941163
transform 1 0 22908 0 1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _1227_
timestamp 1667941163
transform 1 0 21252 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1228__164
timestamp 1667941163
transform 1 0 9108 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1228_
timestamp 1667941163
transform 1 0 9108 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1229_
timestamp 1667941163
transform 1 0 22172 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1230_
timestamp 1667941163
transform 1 0 23092 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1231_
timestamp 1667941163
transform 1 0 21712 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1232__165
timestamp 1667941163
transform 1 0 17388 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1232_
timestamp 1667941163
transform 1 0 17296 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1233_
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1234_
timestamp 1667941163
transform 1 0 18124 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1235_
timestamp 1667941163
transform 1 0 19688 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1236_
timestamp 1667941163
transform 1 0 11684 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1237_
timestamp 1667941163
transform 1 0 27324 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1238_
timestamp 1667941163
transform 1 0 17480 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _1239_
timestamp 1667941163
transform 1 0 15364 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1240_
timestamp 1667941163
transform 1 0 19780 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1241_
timestamp 1667941163
transform 1 0 14628 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1242_
timestamp 1667941163
transform 1 0 29716 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9384 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk
timestamp 1667941163
transform 1 0 5060 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1667941163
transform 1 0 8188 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1667941163
transform 1 0 4692 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1667941163
transform 1 0 7912 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1667941163
transform 1 0 11684 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1667941163
transform 1 0 11684 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1667941163
transform 1 0 15364 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1667941163
transform 1 0 4968 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1667941163
transform 1 0 9844 0 -1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1667941163
transform 1 0 6532 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1667941163
transform 1 0 11316 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1667941163
transform 1 0 15364 0 -1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1667941163
transform 1 0 11960 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1667941163
transform 1 0 14444 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 1564 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 5796 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 12972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1667941163
transform 1 0 1564 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1667941163
transform 1 0 1564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1667941163
transform 1 0 38088 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1667941163
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1667941163
transform 1 0 28520 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1667941163
transform 1 0 38088 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1667941163
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1667941163
transform 1 0 1564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1667941163
transform 1 0 28888 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1667941163
transform 1 0 2392 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1667941163
transform 1 0 10948 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1667941163
transform 1 0 38088 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1667941163
transform 1 0 28428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1667941163
transform 1 0 4600 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1667941163
transform 1 0 36156 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1667941163
transform 1 0 37444 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1667941163
transform 1 0 1564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1667941163
transform 1 0 20700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1667941163
transform 1 0 38088 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1667941163
transform 1 0 38088 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1667941163
transform 1 0 12880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37444 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1667941163
transform 1 0 33028 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1667941163
transform 1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1667941163
transform 1 0 3956 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1667941163
transform 1 0 10948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1667941163
transform 1 0 37996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1667941163
transform 1 0 13524 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1667941163
transform 1 0 31004 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1667941163
transform 1 0 37996 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1667941163
transform 1 0 23276 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1667941163
transform 1 0 9752 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1667941163
transform 1 0 1564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1667941163
transform 1 0 1564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1667941163
transform 1 0 32292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1667941163
transform 1 0 36616 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1667941163
transform 1 0 2300 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1667941163
transform 1 0 38088 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1667941163
transform 1 0 11684 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1667941163
transform 1 0 1564 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1667941163
transform 1 0 1564 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1667941163
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1667941163
transform 1 0 1564 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1667941163
transform 1 0 34868 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1667941163
transform 1 0 37444 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1667941163
transform 1 0 1564 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1667941163
transform 1 0 2300 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1667941163
transform 1 0 37996 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1667941163
transform 1 0 9108 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1667941163
transform 1 0 1564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1667941163
transform 1 0 37260 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1667941163
transform 1 0 14260 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1667941163
transform 1 0 30452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input60
timestamp 1667941163
transform 1 0 3956 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1667941163
transform 1 0 1564 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1667941163
transform 1 0 38088 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 1667941163
transform 1 0 37444 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1667941163
transform 1 0 37444 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1667941163
transform 1 0 32936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1667941163
transform 1 0 1564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1667941163
transform 1 0 37444 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1667941163
transform 1 0 1564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1667941163
transform 1 0 38088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1667941163
transform 1 0 4324 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1667941163
transform 1 0 7268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp 1667941163
transform 1 0 14260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1667941163
transform 1 0 1564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1667941163
transform 1 0 38088 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1667941163
transform 1 0 30360 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1667941163
transform 1 0 1564 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1667941163
transform 1 0 6532 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1667941163
transform 1 0 3956 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1667941163
transform 1 0 1564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1667941163
transform 1 0 38088 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output84 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37996 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 1564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1667941163
transform 1 0 33672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1667941163
transform 1 0 7544 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1667941163
transform 1 0 37996 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1667941163
transform 1 0 16008 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1667941163
transform 1 0 1564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1667941163
transform 1 0 37996 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1667941163
transform 1 0 1564 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1667941163
transform 1 0 1564 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1667941163
transform 1 0 37996 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1667941163
transform 1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1667941163
transform 1 0 37996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1667941163
transform 1 0 37996 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1667941163
transform 1 0 27784 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1667941163
transform 1 0 37260 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1667941163
transform 1 0 17480 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1667941163
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1667941163
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1667941163
transform 1 0 14260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1667941163
transform 1 0 8280 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1667941163
transform 1 0 37996 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1667941163
transform 1 0 36616 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1667941163
transform -1 0 3496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1667941163
transform 1 0 37996 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1667941163
transform 1 0 1564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1667941163
transform 1 0 2852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1667941163
transform 1 0 37996 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1667941163
transform 1 0 37996 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1667941163
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1667941163
transform 1 0 1564 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1667941163
transform -1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1667941163
transform 1 0 1564 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1667941163
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1667941163
transform 1 0 25944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1667941163
transform 1 0 9752 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1667941163
transform 1 0 1564 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1667941163
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1667941163
transform 1 0 2024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1667941163
transform 1 0 1564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1667941163
transform 1 0 21988 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1667941163
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1667941163
transform 1 0 36156 0 1 36992
box -38 -48 406 592
<< labels >>
flabel metal3 s 200 28568 800 28688 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 0 nsew signal input
flabel metal2 s 5814 39200 5870 39800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 1 nsew signal input
flabel metal2 s 12898 200 12954 800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 2 nsew signal input
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 3 nsew signal input
flabel metal3 s 200 26528 800 26648 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
port 4 nsew signal input
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
port 5 nsew signal input
flabel metal3 s 39200 30608 39800 30728 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
port 6 nsew signal input
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
port 7 nsew signal input
flabel metal2 s 25134 39200 25190 39800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 8 nsew signal input
flabel metal3 s 39200 8168 39800 8288 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 9 nsew signal input
flabel metal3 s 200 688 800 808 0 FreeSans 480 0 0 0 ccff_head
port 10 nsew signal input
flabel metal3 s 39200 35368 39800 35488 0 FreeSans 480 0 0 0 ccff_tail
port 11 nsew signal tristate
flabel metal3 s 200 19048 800 19168 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 12 nsew signal input
flabel metal2 s 26422 39200 26478 39800 0 FreeSans 224 90 0 0 chanx_right_in[10]
port 13 nsew signal input
flabel metal3 s 200 23128 800 23248 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 14 nsew signal input
flabel metal2 s 12254 39200 12310 39800 0 FreeSans 224 90 0 0 chanx_right_in[12]
port 15 nsew signal input
flabel metal3 s 39200 10888 39800 11008 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 16 nsew signal input
flabel metal2 s 28354 200 28410 800 0 FreeSans 224 90 0 0 chanx_right_in[14]
port 17 nsew signal input
flabel metal2 s 4526 39200 4582 39800 0 FreeSans 224 90 0 0 chanx_right_in[15]
port 18 nsew signal input
flabel metal2 s 36082 39200 36138 39800 0 FreeSans 224 90 0 0 chanx_right_in[16]
port 19 nsew signal input
flabel metal2 s 37370 39200 37426 39800 0 FreeSans 224 90 0 0 chanx_right_in[17]
port 20 nsew signal input
flabel metal3 s 200 5448 800 5568 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 21 nsew signal input
flabel metal2 s 20626 200 20682 800 0 FreeSans 224 90 0 0 chanx_right_in[1]
port 22 nsew signal input
flabel metal3 s 39200 27888 39800 28008 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 23 nsew signal input
flabel metal3 s 39200 12248 39800 12368 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 24 nsew signal input
flabel metal2 s 15474 39200 15530 39800 0 FreeSans 224 90 0 0 chanx_right_in[4]
port 25 nsew signal input
flabel metal2 s 39302 200 39358 800 0 FreeSans 224 90 0 0 chanx_right_in[5]
port 26 nsew signal input
flabel metal2 s 32862 39200 32918 39800 0 FreeSans 224 90 0 0 chanx_right_in[6]
port 27 nsew signal input
flabel metal2 s 17406 200 17462 800 0 FreeSans 224 90 0 0 chanx_right_in[7]
port 28 nsew signal input
flabel metal2 s 3238 39200 3294 39800 0 FreeSans 224 90 0 0 chanx_right_in[8]
port 29 nsew signal input
flabel metal2 s 10966 200 11022 800 0 FreeSans 224 90 0 0 chanx_right_in[9]
port 30 nsew signal input
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 31 nsew signal tristate
flabel metal2 s 25134 200 25190 800 0 FreeSans 224 90 0 0 chanx_right_out[10]
port 32 nsew signal tristate
flabel metal3 s 39200 12928 39800 13048 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 33 nsew signal tristate
flabel metal3 s 39200 27208 39800 27328 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 34 nsew signal tristate
flabel metal2 s 34794 200 34850 800 0 FreeSans 224 90 0 0 chanx_right_out[13]
port 35 nsew signal tristate
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chanx_right_out[14]
port 36 nsew signal tristate
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 chanx_right_out[15]
port 37 nsew signal tristate
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chanx_right_out[16]
port 38 nsew signal tristate
flabel metal2 s 33506 200 33562 800 0 FreeSans 224 90 0 0 chanx_right_out[17]
port 39 nsew signal tristate
flabel metal3 s 39200 16328 39800 16448 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 40 nsew signal tristate
flabel metal2 s 7746 39200 7802 39800 0 FreeSans 224 90 0 0 chanx_right_out[1]
port 41 nsew signal tristate
flabel metal3 s 39200 23808 39800 23928 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 42 nsew signal tristate
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 chanx_right_out[3]
port 43 nsew signal tristate
flabel metal3 s 39200 32648 39800 32768 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 44 nsew signal tristate
flabel metal3 s 200 4088 800 4208 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 45 nsew signal tristate
flabel metal3 s 39200 17688 39800 17808 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 46 nsew signal tristate
flabel metal3 s 200 31288 800 31408 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 47 nsew signal tristate
flabel metal3 s 200 35368 800 35488 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 48 nsew signal tristate
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 49 nsew signal tristate
flabel metal3 s 39200 1368 39800 1488 0 FreeSans 480 0 0 0 chany_bottom_in[0]
port 50 nsew signal input
flabel metal2 s 21270 39200 21326 39800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 51 nsew signal input
flabel metal2 s 18694 39200 18750 39800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 52 nsew signal input
flabel metal2 s 30930 39200 30986 39800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 53 nsew signal input
flabel metal3 s 39200 37408 39800 37528 0 FreeSans 480 0 0 0 chany_bottom_in[13]
port 54 nsew signal input
flabel metal2 s 23202 39200 23258 39800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 55 nsew signal input
flabel metal2 s 9678 200 9734 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 56 nsew signal input
flabel metal3 s 200 17008 800 17128 0 FreeSans 480 0 0 0 chany_bottom_in[16]
port 57 nsew signal input
flabel metal3 s 200 7488 800 7608 0 FreeSans 480 0 0 0 chany_bottom_in[17]
port 58 nsew signal input
flabel metal2 s 31574 200 31630 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 59 nsew signal input
flabel metal3 s 39200 688 39800 808 0 FreeSans 480 0 0 0 chany_bottom_in[1]
port 60 nsew signal input
flabel metal3 s 200 14968 800 15088 0 FreeSans 480 0 0 0 chany_bottom_in[2]
port 61 nsew signal input
flabel metal3 s 39200 7488 39800 7608 0 FreeSans 480 0 0 0 chany_bottom_in[3]
port 62 nsew signal input
flabel metal2 s 10966 39200 11022 39800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 63 nsew signal input
flabel metal3 s 200 38768 800 38888 0 FreeSans 480 0 0 0 chany_bottom_in[5]
port 64 nsew signal input
flabel metal3 s 200 21768 800 21888 0 FreeSans 480 0 0 0 chany_bottom_in[6]
port 65 nsew signal input
flabel metal2 s 16118 200 16174 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 66 nsew signal input
flabel metal3 s 200 25168 800 25288 0 FreeSans 480 0 0 0 chany_bottom_in[8]
port 67 nsew signal input
flabel metal2 s 34150 39200 34206 39800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 68 nsew signal input
flabel metal2 s 22558 200 22614 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 69 nsew signal tristate
flabel metal2 s 29642 200 29698 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 70 nsew signal tristate
flabel metal3 s 39200 24488 39800 24608 0 FreeSans 480 0 0 0 chany_bottom_out[11]
port 71 nsew signal tristate
flabel metal3 s 39200 4768 39800 4888 0 FreeSans 480 0 0 0 chany_bottom_out[12]
port 72 nsew signal tristate
flabel metal2 s 27710 39200 27766 39800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 73 nsew signal tristate
flabel metal3 s 39200 38768 39800 38888 0 FreeSans 480 0 0 0 chany_bottom_out[14]
port 74 nsew signal tristate
flabel metal2 s 17406 39200 17462 39800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 75 nsew signal tristate
flabel metal2 s 662 200 718 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 76 nsew signal tristate
flabel metal2 s 5170 200 5226 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 77 nsew signal tristate
flabel metal2 s 13542 39200 13598 39800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 78 nsew signal tristate
flabel metal2 s 9034 39200 9090 39800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 79 nsew signal tristate
flabel metal3 s 39200 21088 39800 21208 0 FreeSans 480 0 0 0 chany_bottom_out[2]
port 80 nsew signal tristate
flabel metal3 s 39200 14288 39800 14408 0 FreeSans 480 0 0 0 chany_bottom_out[3]
port 81 nsew signal tristate
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 82 nsew signal tristate
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 83 nsew signal tristate
flabel metal3 s 39200 2728 39800 2848 0 FreeSans 480 0 0 0 chany_bottom_out[6]
port 84 nsew signal tristate
flabel metal3 s 39200 15648 39800 15768 0 FreeSans 480 0 0 0 chany_bottom_out[7]
port 85 nsew signal tristate
flabel metal3 s 200 27208 800 27328 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 86 nsew signal tristate
flabel metal2 s 2594 39200 2650 39800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 87 nsew signal tristate
flabel metal2 s 36726 200 36782 800 0 FreeSans 224 90 0 0 chany_top_in[0]
port 88 nsew signal input
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 chany_top_in[10]
port 89 nsew signal input
flabel metal2 s 18 39200 74 39800 0 FreeSans 224 90 0 0 chany_top_in[11]
port 90 nsew signal input
flabel metal2 s 38658 39200 38714 39800 0 FreeSans 224 90 0 0 chany_top_in[12]
port 91 nsew signal input
flabel metal2 s 8390 200 8446 800 0 FreeSans 224 90 0 0 chany_top_in[13]
port 92 nsew signal input
flabel metal3 s 200 18368 800 18488 0 FreeSans 480 0 0 0 chany_top_in[14]
port 93 nsew signal input
flabel metal2 s 23846 200 23902 800 0 FreeSans 224 90 0 0 chany_top_in[15]
port 94 nsew signal input
flabel metal2 s 38014 200 38070 800 0 FreeSans 224 90 0 0 chany_top_in[16]
port 95 nsew signal input
flabel metal2 s 14186 39200 14242 39800 0 FreeSans 224 90 0 0 chany_top_in[17]
port 96 nsew signal input
flabel metal2 s 30286 200 30342 800 0 FreeSans 224 90 0 0 chany_top_in[18]
port 97 nsew signal input
flabel metal2 s 3882 200 3938 800 0 FreeSans 224 90 0 0 chany_top_in[1]
port 98 nsew signal input
flabel metal3 s 200 13608 800 13728 0 FreeSans 480 0 0 0 chany_top_in[2]
port 99 nsew signal input
flabel metal3 s 39200 4088 39800 4208 0 FreeSans 480 0 0 0 chany_top_in[3]
port 100 nsew signal input
flabel metal3 s 39200 29248 39800 29368 0 FreeSans 480 0 0 0 chany_top_in[4]
port 101 nsew signal input
flabel metal3 s 39200 20408 39800 20528 0 FreeSans 480 0 0 0 chany_top_in[5]
port 102 nsew signal input
flabel metal2 s 32862 200 32918 800 0 FreeSans 224 90 0 0 chany_top_in[6]
port 103 nsew signal input
flabel metal3 s 200 23808 800 23928 0 FreeSans 480 0 0 0 chany_top_in[7]
port 104 nsew signal input
flabel metal3 s 39200 9528 39800 9648 0 FreeSans 480 0 0 0 chany_top_in[8]
port 105 nsew signal input
flabel metal3 s 200 31968 800 32088 0 FreeSans 480 0 0 0 chany_top_in[9]
port 106 nsew signal input
flabel metal3 s 39200 22448 39800 22568 0 FreeSans 480 0 0 0 chany_top_out[0]
port 107 nsew signal tristate
flabel metal3 s 39200 34008 39800 34128 0 FreeSans 480 0 0 0 chany_top_out[10]
port 108 nsew signal tristate
flabel metal2 s 36082 200 36138 800 0 FreeSans 224 90 0 0 chany_top_out[11]
port 109 nsew signal tristate
flabel metal3 s 39200 36048 39800 36168 0 FreeSans 480 0 0 0 chany_top_out[12]
port 110 nsew signal tristate
flabel metal3 s 200 33328 800 33448 0 FreeSans 480 0 0 0 chany_top_out[13]
port 111 nsew signal tristate
flabel metal3 s 200 2048 800 2168 0 FreeSans 480 0 0 0 chany_top_out[14]
port 112 nsew signal tristate
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 chany_top_out[15]
port 113 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_top_out[16]
port 114 nsew signal tristate
flabel metal2 s 25778 200 25834 800 0 FreeSans 224 90 0 0 chany_top_out[17]
port 115 nsew signal tristate
flabel metal3 s 200 38088 800 38208 0 FreeSans 480 0 0 0 chany_top_out[18]
port 116 nsew signal tristate
flabel metal2 s 9678 39200 9734 39800 0 FreeSans 224 90 0 0 chany_top_out[1]
port 117 nsew signal tristate
flabel metal2 s 24490 39200 24546 39800 0 FreeSans 224 90 0 0 chany_top_out[2]
port 118 nsew signal tristate
flabel metal3 s 200 29928 800 30048 0 FreeSans 480 0 0 0 chany_top_out[3]
port 119 nsew signal tristate
flabel metal2 s 6458 200 6514 800 0 FreeSans 224 90 0 0 chany_top_out[4]
port 120 nsew signal tristate
flabel metal2 s 1950 200 2006 800 0 FreeSans 224 90 0 0 chany_top_out[5]
port 121 nsew signal tristate
flabel metal3 s 200 8848 800 8968 0 FreeSans 480 0 0 0 chany_top_out[6]
port 122 nsew signal tristate
flabel metal2 s 21914 39200 21970 39800 0 FreeSans 224 90 0 0 chany_top_out[7]
port 123 nsew signal tristate
flabel metal2 s 18050 200 18106 800 0 FreeSans 224 90 0 0 chany_top_out[8]
port 124 nsew signal tristate
flabel metal2 s 35438 39200 35494 39800 0 FreeSans 224 90 0 0 chany_top_out[9]
port 125 nsew signal tristate
flabel metal3 s 39200 6128 39800 6248 0 FreeSans 480 0 0 0 pReset
port 126 nsew signal input
flabel metal3 s 200 36728 800 36848 0 FreeSans 480 0 0 0 prog_clk
port 127 nsew signal input
flabel metal3 s 200 11568 800 11688 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 128 nsew signal input
flabel metal2 s 7102 200 7158 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 129 nsew signal input
flabel metal2 s 14186 200 14242 800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 130 nsew signal input
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 131 nsew signal input
flabel metal3 s 39200 25848 39800 25968 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 132 nsew signal input
flabel metal2 s 21914 200 21970 800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 133 nsew signal input
flabel metal2 s 29642 39200 29698 39800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 134 nsew signal input
flabel metal2 s 28354 39200 28410 39800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 135 nsew signal input
flabel metal2 s 1306 39200 1362 39800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
port 136 nsew signal input
flabel metal2 s 6458 39200 6514 39800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
port 137 nsew signal input
flabel metal2 s 27066 200 27122 800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
port 138 nsew signal input
flabel metal3 s 200 10208 800 10328 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
port 139 nsew signal input
flabel metal3 s 200 34688 800 34808 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 140 nsew signal input
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 141 nsew signal input
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 142 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 142 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 143 nsew ground bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel via2 5382 31365 5382 31365 0 _0000_
rlabel metal1 16468 34714 16468 34714 0 _0001_
rlabel metal1 17671 30634 17671 30634 0 _0002_
rlabel metal1 18821 30294 18821 30294 0 _0003_
rlabel metal2 20470 36380 20470 36380 0 _0004_
rlabel metal2 20746 35309 20746 35309 0 _0005_
rlabel metal2 19366 36244 19366 36244 0 _0006_
rlabel metal1 16889 33898 16889 33898 0 _0007_
rlabel metal2 17434 33796 17434 33796 0 _0008_
rlabel metal1 6447 28458 6447 28458 0 _0009_
rlabel metal1 17519 35734 17519 35734 0 _0010_
rlabel metal1 16599 36822 16599 36822 0 _0011_
rlabel metal2 20930 36108 20930 36108 0 _0012_
rlabel metal1 21068 36550 21068 36550 0 _0013_
rlabel metal2 10534 32164 10534 32164 0 _0014_
rlabel metal1 11730 27513 11730 27513 0 _0015_
rlabel metal1 9752 24310 9752 24310 0 _0016_
rlabel metal1 5750 26928 5750 26928 0 _0017_
rlabel via2 5382 30685 5382 30685 0 _0018_
rlabel metal1 12565 32810 12565 32810 0 _0019_
rlabel metal2 17434 34918 17434 34918 0 _0020_
rlabel metal2 18170 34170 18170 34170 0 _0021_
rlabel metal1 8832 15878 8832 15878 0 _0022_
rlabel metal2 7774 17986 7774 17986 0 _0023_
rlabel metal2 7498 18496 7498 18496 0 _0024_
rlabel metal1 6762 16490 6762 16490 0 _0025_
rlabel metal1 9154 15674 9154 15674 0 _0026_
rlabel metal1 8609 24106 8609 24106 0 _0027_
rlabel metal2 13846 32198 13846 32198 0 _0028_
rlabel metal2 14950 35292 14950 35292 0 _0029_
rlabel metal2 19366 35105 19366 35105 0 _0030_
rlabel metal2 18906 34221 18906 34221 0 _0031_
rlabel via1 15134 35717 15134 35717 0 _0032_
rlabel metal1 11277 29546 11277 29546 0 _0033_
rlabel metal2 10718 27846 10718 27846 0 _0034_
rlabel metal1 6838 27370 6838 27370 0 _0035_
rlabel metal1 3220 14042 3220 14042 0 _0036_
rlabel metal1 5382 15062 5382 15062 0 _0037_
rlabel metal1 7498 15538 7498 15538 0 _0038_
rlabel metal1 5566 14450 5566 14450 0 _0039_
rlabel metal1 20792 28730 20792 28730 0 _0040_
rlabel metal1 16744 23834 16744 23834 0 _0041_
rlabel metal1 3135 22678 3135 22678 0 _0042_
rlabel metal1 4554 14518 4554 14518 0 _0043_
rlabel metal2 8234 17986 8234 17986 0 _0044_
rlabel metal1 9253 30634 9253 30634 0 _0045_
rlabel metal1 14267 25262 14267 25262 0 _0046_
rlabel metal1 17487 34986 17487 34986 0 _0047_
rlabel metal1 10396 17850 10396 17850 0 _0048_
rlabel metal1 17579 23086 17579 23086 0 _0049_
rlabel metal2 19366 32640 19366 32640 0 _0050_
rlabel metal1 18676 34170 18676 34170 0 _0051_
rlabel metal2 14398 17612 14398 17612 0 _0052_
rlabel metal1 16935 28118 16935 28118 0 _0053_
rlabel metal1 16705 19754 16705 19754 0 _0054_
rlabel metal2 15502 17000 15502 17000 0 _0055_
rlabel metal1 16836 15130 16836 15130 0 _0056_
rlabel metal1 18630 16490 18630 16490 0 _0057_
rlabel metal2 16790 17000 16790 17000 0 _0058_
rlabel metal2 21666 18224 21666 18224 0 _0059_
rlabel metal1 12374 25976 12374 25976 0 _0060_
rlabel metal2 14582 17816 14582 17816 0 _0061_
rlabel metal1 16882 30906 16882 30906 0 _0062_
rlabel metal2 11546 29342 11546 29342 0 _0063_
rlabel via1 19918 32997 19918 32997 0 _0064_
rlabel via2 20562 32963 20562 32963 0 _0065_
rlabel metal1 17763 29614 17763 29614 0 _0066_
rlabel metal2 21022 25262 21022 25262 0 _0067_
rlabel metal1 10488 16218 10488 16218 0 _0068_
rlabel metal2 12650 19074 12650 19074 0 _0069_
rlabel metal2 14674 19550 14674 19550 0 _0070_
rlabel metal2 17158 26554 17158 26554 0 _0071_
rlabel metal1 19596 34646 19596 34646 0 _0072_
rlabel metal1 17579 31790 17579 31790 0 _0073_
rlabel metal2 18814 35394 18814 35394 0 _0074_
rlabel metal1 17671 32810 17671 32810 0 _0075_
rlabel metal2 19366 34204 19366 34204 0 _0076_
rlabel metal1 15134 36074 15134 36074 0 _0077_
rlabel metal1 20194 35462 20194 35462 0 _0078_
rlabel metal1 4876 15130 4876 15130 0 _0079_
rlabel metal1 5014 16150 5014 16150 0 _0080_
rlabel metal2 5290 19074 5290 19074 0 _0081_
rlabel metal1 6670 16218 6670 16218 0 _0082_
rlabel metal2 6762 19346 6762 19346 0 _0083_
rlabel metal1 18584 21114 18584 21114 0 _0084_
rlabel metal1 18131 24174 18131 24174 0 _0085_
rlabel metal1 18499 25194 18499 25194 0 _0086_
rlabel metal1 19688 28390 19688 28390 0 _0087_
rlabel metal1 6210 15606 6210 15606 0 _0088_
rlabel metal1 5612 16422 5612 16422 0 _0089_
rlabel metal1 8142 15062 8142 15062 0 _0090_
rlabel metal2 12098 31314 12098 31314 0 _0091_
rlabel metal2 12374 29631 12374 29631 0 _0092_
rlabel metal2 3358 17000 3358 17000 0 _0093_
rlabel metal1 8280 15674 8280 15674 0 _0094_
rlabel metal2 9798 24582 9798 24582 0 _0095_
rlabel metal1 7498 14790 7498 14790 0 _0096_
rlabel metal1 5336 15674 5336 15674 0 _0097_
rlabel metal1 9292 15062 9292 15062 0 _0098_
rlabel metal1 13386 26391 13386 26391 0 _0099_
rlabel metal1 11914 23127 11914 23127 0 _0100_
rlabel metal2 12558 17068 12558 17068 0 _0101_
rlabel metal2 21390 25160 21390 25160 0 _0102_
rlabel metal1 17073 20842 17073 20842 0 _0103_
rlabel metal2 20654 34510 20654 34510 0 _0104_
rlabel metal2 21298 34697 21298 34697 0 _0105_
rlabel metal1 18998 32368 18998 32368 0 _0106_
rlabel metal1 18216 31110 18216 31110 0 _0107_
rlabel metal1 18131 28458 18131 28458 0 _0108_
rlabel metal1 14589 28458 14589 28458 0 _0109_
rlabel metal1 10718 22569 10718 22569 0 _0110_
rlabel metal2 17986 21216 17986 21216 0 _0111_
rlabel metal1 3503 23018 3503 23018 0 _0112_
rlabel metal2 2484 19652 2484 19652 0 _0113_
rlabel metal1 5106 14042 5106 14042 0 _0114_
rlabel metal1 2162 11798 2162 11798 0 _0115_
rlabel metal1 9897 26350 9897 26350 0 _0116_
rlabel via2 4094 29189 4094 29189 0 _0117_
rlabel metal1 21344 25874 21344 25874 0 _0118_
rlabel metal2 19320 18428 19320 18428 0 _0119_
rlabel metal1 20884 36142 20884 36142 0 _0120_
rlabel metal1 18078 34578 18078 34578 0 _0121_
rlabel metal1 15548 36142 15548 36142 0 _0122_
rlabel metal2 16882 23647 16882 23647 0 _0123_
rlabel metal1 19136 21454 19136 21454 0 _0124_
rlabel metal2 21574 18309 21574 18309 0 _0125_
rlabel metal2 25806 27404 25806 27404 0 _0126_
rlabel metal1 9108 34714 9108 34714 0 _0127_
rlabel metal2 23782 31110 23782 31110 0 _0128_
rlabel metal2 4002 36550 4002 36550 0 _0129_
rlabel metal1 26082 22202 26082 22202 0 _0130_
rlabel metal2 31786 20740 31786 20740 0 _0131_
rlabel metal1 16974 11866 16974 11866 0 _0132_
rlabel metal2 25438 10234 25438 10234 0 _0133_
rlabel metal2 26266 9146 26266 9146 0 _0134_
rlabel metal2 18722 10268 18722 10268 0 _0135_
rlabel metal1 26726 16422 26726 16422 0 _0136_
rlabel metal1 24242 10234 24242 10234 0 _0137_
rlabel metal1 15686 12410 15686 12410 0 _0138_
rlabel metal1 26358 17612 26358 17612 0 _0139_
rlabel metal2 25806 16252 25806 16252 0 _0140_
rlabel metal1 15824 8466 15824 8466 0 _0141_
rlabel metal1 24150 10676 24150 10676 0 _0142_
rlabel metal1 28382 10676 28382 10676 0 _0143_
rlabel metal2 28934 23324 28934 23324 0 _0144_
rlabel metal2 29762 30022 29762 30022 0 _0145_
rlabel metal1 30682 31348 30682 31348 0 _0146_
rlabel metal1 23276 6630 23276 6630 0 _0147_
rlabel metal2 11730 6970 11730 6970 0 _0148_
rlabel metal1 13616 6290 13616 6290 0 _0149_
rlabel metal2 29026 14586 29026 14586 0 _0150_
rlabel metal1 29946 25228 29946 25228 0 _0151_
rlabel metal2 28566 25466 28566 25466 0 _0152_
rlabel metal2 20378 20060 20378 20060 0 _0153_
rlabel metal1 18308 21930 18308 21930 0 _0154_
rlabel metal1 20332 21930 20332 21930 0 _0155_
rlabel metal1 18354 17544 18354 17544 0 _0156_
rlabel metal2 20654 18496 20654 18496 0 _0157_
rlabel metal2 27646 28730 27646 28730 0 _0158_
rlabel metal1 24334 26010 24334 26010 0 _0159_
rlabel metal1 32430 26248 32430 26248 0 _0160_
rlabel metal2 25346 31518 25346 31518 0 _0161_
rlabel metal2 20654 21352 20654 21352 0 _0162_
rlabel metal1 19504 18598 19504 18598 0 _0163_
rlabel metal2 27370 35054 27370 35054 0 _0164_
rlabel metal1 20930 22678 20930 22678 0 _0165_
rlabel metal1 26358 33082 26358 33082 0 _0166_
rlabel metal1 27370 28152 27370 28152 0 _0167_
rlabel metal1 13248 15402 13248 15402 0 _0168_
rlabel metal1 24150 26350 24150 26350 0 _0169_
rlabel metal1 17480 17306 17480 17306 0 _0170_
rlabel metal2 22402 17408 22402 17408 0 _0171_
rlabel metal1 3174 7446 3174 7446 0 _0172_
rlabel metal1 25852 26554 25852 26554 0 _0173_
rlabel metal2 27462 15912 27462 15912 0 _0174_
rlabel metal1 24886 23834 24886 23834 0 _0175_
rlabel metal1 26036 7786 26036 7786 0 _0176_
rlabel metal1 27416 20570 27416 20570 0 _0177_
rlabel metal1 20746 11050 20746 11050 0 _0178_
rlabel metal2 17342 11560 17342 11560 0 _0179_
rlabel metal2 21298 28696 21298 28696 0 _0180_
rlabel metal2 21666 10234 21666 10234 0 _0181_
rlabel metal2 10074 14552 10074 14552 0 _0182_
rlabel metal1 11454 11152 11454 11152 0 _0183_
rlabel metal1 10120 11050 10120 11050 0 _0184_
rlabel metal1 4692 10778 4692 10778 0 _0185_
rlabel metal1 3910 13498 3910 13498 0 _0186_
rlabel metal1 21390 32776 21390 32776 0 _0187_
rlabel metal2 4646 10642 4646 10642 0 _0188_
rlabel metal2 23322 13804 23322 13804 0 _0189_
rlabel metal1 24840 28526 24840 28526 0 _0190_
rlabel metal1 11362 13498 11362 13498 0 _0191_
rlabel metal1 24794 21896 24794 21896 0 _0192_
rlabel metal1 27600 32810 27600 32810 0 _0193_
rlabel metal2 15594 13090 15594 13090 0 _0194_
rlabel metal1 16928 5270 16928 5270 0 _0195_
rlabel metal1 14352 9962 14352 9962 0 _0196_
rlabel metal1 23736 15674 23736 15674 0 _0197_
rlabel metal1 11224 11322 11224 11322 0 _0198_
rlabel metal1 23920 30294 23920 30294 0 _0199_
rlabel metal2 23782 13022 23782 13022 0 _0200_
rlabel metal1 17250 10710 17250 10710 0 _0201_
rlabel metal1 23598 14314 23598 14314 0 _0202_
rlabel metal1 17986 13974 17986 13974 0 _0203_
rlabel metal2 21758 30226 21758 30226 0 _0204_
rlabel metal2 20930 18190 20930 18190 0 _0205_
rlabel metal1 24748 32742 24748 32742 0 _0206_
rlabel metal2 13386 36873 13386 36873 0 _0207_
rlabel metal1 25208 34170 25208 34170 0 _0208_
rlabel metal1 23552 28458 23552 28458 0 _0209_
rlabel metal1 26312 28458 26312 28458 0 _0210_
rlabel metal2 30406 16456 30406 16456 0 _0211_
rlabel metal1 26956 22678 26956 22678 0 _0212_
rlabel metal2 18446 19414 18446 19414 0 _0213_
rlabel metal2 27554 19992 27554 19992 0 _0214_
rlabel viali 22214 27370 22214 27370 0 _0215_
rlabel metal1 20286 12614 20286 12614 0 _0216_
rlabel metal1 18078 12954 18078 12954 0 _0217_
rlabel metal1 1840 9690 1840 9690 0 _0218_
rlabel metal1 2208 10234 2208 10234 0 _0219_
rlabel metal1 3036 9622 3036 9622 0 _0220_
rlabel metal1 2254 7752 2254 7752 0 _0221_
rlabel metal2 25622 28696 25622 28696 0 _0222_
rlabel metal1 2668 26282 2668 26282 0 _0223_
rlabel metal1 8142 12342 8142 12342 0 _0224_
rlabel metal1 17848 12886 17848 12886 0 _0225_
rlabel metal2 12466 14382 12466 14382 0 _0226_
rlabel metal1 1978 15096 1978 15096 0 _0227_
rlabel metal1 26358 30600 26358 30600 0 _0228_
rlabel metal1 8740 13498 8740 13498 0 _0229_
rlabel metal1 23506 29206 23506 29206 0 _0230_
rlabel metal1 32062 28424 32062 28424 0 _0231_
rlabel metal2 29946 23290 29946 23290 0 _0232_
rlabel metal1 27784 36074 27784 36074 0 _0233_
rlabel metal2 27278 36176 27278 36176 0 _0234_
rlabel metal2 13018 36125 13018 36125 0 _0235_
rlabel via2 19826 27387 19826 27387 0 _0236_
rlabel metal1 17434 24854 17434 24854 0 _0237_
rlabel metal1 6716 15062 6716 15062 0 _0238_
rlabel metal1 18952 26010 18952 26010 0 _0239_
rlabel metal1 23230 24854 23230 24854 0 _0240_
rlabel metal2 20838 26078 20838 26078 0 _0241_
rlabel metal1 20194 31722 20194 31722 0 _0242_
rlabel metal1 23368 30158 23368 30158 0 _0243_
rlabel metal2 19918 13872 19918 13872 0 _0244_
rlabel metal1 18354 23800 18354 23800 0 _0245_
rlabel metal1 20056 9622 20056 9622 0 _0246_
rlabel metal1 20286 31450 20286 31450 0 _0247_
rlabel metal1 28106 33626 28106 33626 0 _0248_
rlabel metal1 23460 33898 23460 33898 0 _0249_
rlabel metal2 24794 35054 24794 35054 0 _0250_
rlabel metal1 24472 26554 24472 26554 0 _0251_
rlabel metal1 17066 13838 17066 13838 0 _0252_
rlabel metal1 26128 33626 26128 33626 0 _0253_
rlabel metal1 8188 16150 8188 16150 0 _0254_
rlabel metal1 8096 14042 8096 14042 0 _0255_
rlabel metal1 26266 32776 26266 32776 0 _0256_
rlabel metal1 20562 33592 20562 33592 0 _0257_
rlabel metal2 28842 36312 28842 36312 0 _0258_
rlabel metal2 25162 34170 25162 34170 0 _0259_
rlabel metal1 27876 23766 27876 23766 0 _0260_
rlabel metal2 4738 14756 4738 14756 0 _0261_
rlabel metal2 2622 14994 2622 14994 0 _0262_
rlabel metal1 29486 33286 29486 33286 0 _0263_
rlabel metal1 21942 24072 21942 24072 0 _0264_
rlabel metal2 6486 36312 6486 36312 0 _0265_
rlabel metal1 16284 14314 16284 14314 0 _0266_
rlabel metal2 2438 10880 2438 10880 0 _0267_
rlabel metal1 20378 15402 20378 15402 0 _0268_
rlabel metal1 5934 10778 5934 10778 0 _0269_
rlabel metal2 7682 14110 7682 14110 0 _0270_
rlabel metal2 19642 14586 19642 14586 0 _0271_
rlabel metal1 22540 33558 22540 33558 0 _0272_
rlabel metal1 25162 35258 25162 35258 0 _0273_
rlabel metal2 7958 36584 7958 36584 0 _0274_
rlabel metal1 5980 13498 5980 13498 0 _0275_
rlabel metal1 21206 36108 21206 36108 0 _0276_
rlabel metal2 18170 29121 18170 29121 0 _0277_
rlabel metal2 25990 13736 25990 13736 0 _0278_
rlabel metal1 22264 18938 22264 18938 0 _0279_
rlabel metal1 20884 29682 20884 29682 0 _0280_
rlabel metal2 22586 10200 22586 10200 0 _0281_
rlabel metal1 8050 11016 8050 11016 0 _0282_
rlabel metal1 14306 10778 14306 10778 0 _0283_
rlabel metal1 18032 15674 18032 15674 0 _0284_
rlabel metal2 14766 12002 14766 12002 0 _0285_
rlabel metal1 2990 10234 2990 10234 0 _0286_
rlabel metal1 12742 15062 12742 15062 0 _0287_
rlabel metal1 22264 21930 22264 21930 0 _0288_
rlabel metal1 2300 9622 2300 9622 0 _0289_
rlabel metal1 1794 11322 1794 11322 0 _0290_
rlabel metal1 5382 14382 5382 14382 0 _0291_
rlabel metal2 12006 14824 12006 14824 0 _0292_
rlabel metal1 7130 12410 7130 12410 0 _0293_
rlabel metal1 29946 25466 29946 25466 0 _0294_
rlabel metal2 28658 24616 28658 24616 0 _0295_
rlabel metal2 28474 14076 28474 14076 0 _0296_
rlabel metal1 30222 25874 30222 25874 0 _0297_
rlabel metal1 26404 31994 26404 31994 0 _0298_
rlabel metal2 29946 17068 29946 17068 0 _0299_
rlabel metal1 11822 6970 11822 6970 0 _0300_
rlabel metal1 13156 6426 13156 6426 0 _0301_
rlabel metal2 23506 7208 23506 7208 0 _0302_
rlabel metal1 12788 8398 12788 8398 0 _0303_
rlabel metal2 14490 9146 14490 9146 0 _0304_
rlabel metal1 23230 8840 23230 8840 0 _0305_
rlabel metal2 29302 30532 29302 30532 0 _0306_
rlabel metal1 29072 31246 29072 31246 0 _0307_
rlabel metal2 28750 22916 28750 22916 0 _0308_
rlabel metal2 28198 29852 28198 29852 0 _0309_
rlabel metal2 29026 32164 29026 32164 0 _0310_
rlabel metal1 28934 27574 28934 27574 0 _0311_
rlabel metal1 24380 10778 24380 10778 0 _0312_
rlabel metal1 28290 10778 28290 10778 0 _0313_
rlabel metal2 15410 9044 15410 9044 0 _0314_
rlabel metal2 20746 9758 20746 9758 0 _0315_
rlabel metal2 28106 17340 28106 17340 0 _0316_
rlabel metal1 19228 9010 19228 9010 0 _0317_
rlabel metal1 27324 16150 27324 16150 0 _0318_
rlabel metal1 25898 16218 25898 16218 0 _0319_
rlabel metal1 14766 12954 14766 12954 0 _0320_
rlabel metal2 23506 16286 23506 16286 0 _0321_
rlabel metal1 22862 16218 22862 16218 0 _0322_
rlabel metal2 21022 15028 21022 15028 0 _0323_
rlabel metal1 26818 12138 26818 12138 0 _0324_
rlabel metal1 25070 10506 25070 10506 0 _0325_
rlabel metal2 17802 10268 17802 10268 0 _0326_
rlabel metal2 24794 14552 24794 14552 0 _0327_
rlabel metal2 22218 11356 22218 11356 0 _0328_
rlabel metal1 20240 10098 20240 10098 0 _0329_
rlabel metal2 25254 10472 25254 10472 0 _0330_
rlabel metal2 26542 9316 26542 9316 0 _0331_
rlabel metal2 16882 13056 16882 13056 0 _0332_
rlabel metal1 22770 12104 22770 12104 0 _0333_
rlabel metal2 25990 9282 25990 9282 0 _0334_
rlabel metal1 22172 20570 22172 20570 0 _0335_
rlabel metal1 31464 20434 31464 20434 0 _0336_
rlabel metal1 25990 22746 25990 22746 0 _0337_
rlabel metal1 30544 20978 30544 20978 0 _0338_
rlabel metal1 26036 20570 26036 20570 0 _0339_
rlabel metal2 4922 36312 4922 36312 0 _0340_
rlabel metal1 22724 31246 22724 31246 0 _0341_
rlabel metal1 18262 34952 18262 34952 0 _0342_
rlabel metal1 21068 23766 21068 23766 0 _0343_
rlabel via2 9338 35003 9338 35003 0 _0344_
rlabel metal1 25208 26826 25208 26826 0 _0345_
rlabel metal1 25300 35190 25300 35190 0 _0346_
rlabel via2 24978 28203 24978 28203 0 _0347_
rlabel metal2 17618 6596 17618 6596 0 _0348_
rlabel metal2 11362 10472 11362 10472 0 _0349_
rlabel metal1 18492 20774 18492 20774 0 _0350_
rlabel metal1 18998 6426 18998 6426 0 _0351_
rlabel metal2 11914 8942 11914 8942 0 _0352_
rlabel metal1 24288 23630 24288 23630 0 _0353_
rlabel metal1 17572 27098 17572 27098 0 _0354_
rlabel metal2 15686 6596 15686 6596 0 _0355_
rlabel metal2 21022 17816 21022 17816 0 _0356_
rlabel metal1 14812 7514 14812 7514 0 _0357_
rlabel metal2 23598 16286 23598 16286 0 _0358_
rlabel metal3 1234 28628 1234 28628 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 5934 37230 5934 37230 0 bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 12926 1588 12926 1588 0 bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 19366 1588 19366 1588 0 bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal3 1234 26588 1234 26588 0 bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal3 1234 6868 1234 6868 0 bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
rlabel via2 38318 30685 38318 30685 0 bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal2 11638 1588 11638 1588 0 bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal1 28336 37230 28336 37230 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 38318 8347 38318 8347 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
rlabel metal3 1740 748 1740 748 0 ccff_head
rlabel via2 38226 35445 38226 35445 0 ccff_tail
rlabel metal3 1234 19108 1234 19108 0 chanx_right_in[0]
rlabel metal1 28888 36754 28888 36754 0 chanx_right_in[10]
rlabel metal3 1740 23188 1740 23188 0 chanx_right_in[11]
rlabel metal1 11730 37230 11730 37230 0 chanx_right_in[12]
rlabel metal2 38318 11033 38318 11033 0 chanx_right_in[13]
rlabel metal2 28382 1588 28382 1588 0 chanx_right_in[14]
rlabel metal1 4738 37230 4738 37230 0 chanx_right_in[15]
rlabel metal1 36248 36142 36248 36142 0 chanx_right_in[16]
rlabel metal1 37536 35054 37536 35054 0 chanx_right_in[17]
rlabel metal3 1234 5508 1234 5508 0 chanx_right_in[18]
rlabel metal2 20654 1588 20654 1588 0 chanx_right_in[1]
rlabel metal2 38318 27999 38318 27999 0 chanx_right_in[2]
rlabel metal2 38318 12563 38318 12563 0 chanx_right_in[3]
rlabel metal1 13110 37196 13110 37196 0 chanx_right_in[4]
rlabel metal2 39330 1894 39330 1894 0 chanx_right_in[5]
rlabel metal1 33074 37230 33074 37230 0 chanx_right_in[6]
rlabel metal2 17434 1588 17434 1588 0 chanx_right_in[7]
rlabel metal1 3726 37230 3726 37230 0 chanx_right_in[8]
rlabel metal2 10994 1588 10994 1588 0 chanx_right_in[9]
rlabel metal3 1234 15708 1234 15708 0 chanx_right_out[0]
rlabel metal2 25162 1520 25162 1520 0 chanx_right_out[10]
rlabel metal2 38226 13073 38226 13073 0 chanx_right_out[11]
rlabel via2 38226 27285 38226 27285 0 chanx_right_out[12]
rlabel metal2 34822 1520 34822 1520 0 chanx_right_out[13]
rlabel metal2 14858 1520 14858 1520 0 chanx_right_out[14]
rlabel metal1 32384 37094 32384 37094 0 chanx_right_out[15]
rlabel metal1 20148 37094 20148 37094 0 chanx_right_out[16]
rlabel metal2 33534 1520 33534 1520 0 chanx_right_out[17]
rlabel via2 38226 16405 38226 16405 0 chanx_right_out[18]
rlabel metal2 7774 38158 7774 38158 0 chanx_right_out[1]
rlabel metal2 38226 23953 38226 23953 0 chanx_right_out[2]
rlabel metal1 16514 37094 16514 37094 0 chanx_right_out[3]
rlabel via2 38226 32725 38226 32725 0 chanx_right_out[4]
rlabel metal3 1234 4148 1234 4148 0 chanx_right_out[5]
rlabel metal2 38226 17901 38226 17901 0 chanx_right_out[6]
rlabel metal3 1234 31348 1234 31348 0 chanx_right_out[7]
rlabel metal2 1794 35343 1794 35343 0 chanx_right_out[8]
rlabel metal2 38226 32113 38226 32113 0 chanx_right_out[9]
rlabel metal1 37674 4182 37674 4182 0 chany_bottom_in[0]
rlabel metal1 21666 37298 21666 37298 0 chany_bottom_in[10]
rlabel metal1 13938 37230 13938 37230 0 chany_bottom_in[11]
rlabel metal1 31096 37230 31096 37230 0 chany_bottom_in[12]
rlabel metal2 38134 37349 38134 37349 0 chany_bottom_in[13]
rlabel metal1 23322 37230 23322 37230 0 chany_bottom_in[14]
rlabel metal1 9844 3026 9844 3026 0 chany_bottom_in[15]
rlabel metal3 1188 17068 1188 17068 0 chany_bottom_in[16]
rlabel metal3 1234 7548 1234 7548 0 chany_bottom_in[17]
rlabel metal2 31602 1588 31602 1588 0 chany_bottom_in[18]
rlabel metal1 37030 3026 37030 3026 0 chany_bottom_in[1]
rlabel metal3 1602 15028 1602 15028 0 chany_bottom_in[2]
rlabel metal2 38318 7701 38318 7701 0 chany_bottom_in[3]
rlabel metal1 11454 37162 11454 37162 0 chany_bottom_in[4]
rlabel metal3 1142 38828 1142 38828 0 chany_bottom_in[5]
rlabel metal3 1188 21828 1188 21828 0 chany_bottom_in[6]
rlabel metal2 16146 1588 16146 1588 0 chany_bottom_in[7]
rlabel metal3 1188 25228 1188 25228 0 chany_bottom_in[8]
rlabel metal1 34546 37298 34546 37298 0 chany_bottom_in[9]
rlabel metal2 22586 1520 22586 1520 0 chany_bottom_out[0]
rlabel metal2 29670 1520 29670 1520 0 chany_bottom_out[10]
rlabel via2 38226 24565 38226 24565 0 chany_bottom_out[11]
rlabel metal2 38226 4913 38226 4913 0 chany_bottom_out[12]
rlabel metal1 27876 37094 27876 37094 0 chany_bottom_out[13]
rlabel metal1 37352 36346 37352 36346 0 chany_bottom_out[14]
rlabel metal1 17572 37094 17572 37094 0 chany_bottom_out[15]
rlabel metal2 690 1792 690 1792 0 chany_bottom_out[16]
rlabel metal2 5198 1520 5198 1520 0 chany_bottom_out[17]
rlabel metal1 14168 37094 14168 37094 0 chany_bottom_out[18]
rlabel metal1 8786 37094 8786 37094 0 chany_bottom_out[1]
rlabel metal2 38226 21233 38226 21233 0 chany_bottom_out[2]
rlabel metal2 38226 14297 38226 14297 0 chany_bottom_out[3]
rlabel metal1 38088 36890 38088 36890 0 chany_bottom_out[4]
rlabel metal2 3266 1520 3266 1520 0 chany_bottom_out[5]
rlabel metal2 38226 3077 38226 3077 0 chany_bottom_out[6]
rlabel metal2 38226 15793 38226 15793 0 chany_bottom_out[7]
rlabel metal3 1234 27268 1234 27268 0 chany_bottom_out[8]
rlabel metal2 2622 38209 2622 38209 0 chany_bottom_out[9]
rlabel metal2 36754 1588 36754 1588 0 chany_top_in[0]
rlabel metal3 1188 20468 1188 20468 0 chany_top_in[10]
rlabel metal1 2116 36754 2116 36754 0 chany_top_in[11]
rlabel metal1 38410 36822 38410 36822 0 chany_top_in[12]
rlabel metal2 8418 1588 8418 1588 0 chany_top_in[13]
rlabel metal3 1188 18428 1188 18428 0 chany_top_in[14]
rlabel metal2 23874 1588 23874 1588 0 chany_top_in[15]
rlabel metal2 38042 2064 38042 2064 0 chany_top_in[16]
rlabel metal1 14398 35054 14398 35054 0 chany_top_in[17]
rlabel metal2 30314 1588 30314 1588 0 chany_top_in[18]
rlabel metal2 3910 1588 3910 1588 0 chany_top_in[1]
rlabel metal3 1188 13668 1188 13668 0 chany_top_in[2]
rlabel metal2 38318 4369 38318 4369 0 chany_top_in[3]
rlabel metal2 37490 29461 37490 29461 0 chany_top_in[4]
rlabel metal1 37352 20910 37352 20910 0 chany_top_in[5]
rlabel metal2 32890 1554 32890 1554 0 chany_top_in[6]
rlabel metal3 1234 23868 1234 23868 0 chany_top_in[7]
rlabel metal1 37352 10030 37352 10030 0 chany_top_in[8]
rlabel metal3 1188 32028 1188 32028 0 chany_top_in[9]
rlabel via2 38226 22491 38226 22491 0 chany_top_out[0]
rlabel metal2 38226 34221 38226 34221 0 chany_top_out[10]
rlabel metal2 36110 1520 36110 1520 0 chany_top_out[11]
rlabel metal2 38226 36057 38226 36057 0 chany_top_out[12]
rlabel metal3 1234 33388 1234 33388 0 chany_top_out[13]
rlabel metal3 1188 2108 1188 2108 0 chany_top_out[14]
rlabel metal3 1234 12308 1234 12308 0 chany_top_out[15]
rlabel metal2 46 1826 46 1826 0 chany_top_out[16]
rlabel metal2 25806 1520 25806 1520 0 chany_top_out[17]
rlabel metal2 1794 37519 1794 37519 0 chany_top_out[18]
rlabel metal1 9844 37094 9844 37094 0 chany_top_out[1]
rlabel metal1 24656 37094 24656 37094 0 chany_top_out[2]
rlabel metal3 1234 29988 1234 29988 0 chany_top_out[3]
rlabel metal2 6486 1520 6486 1520 0 chany_top_out[4]
rlabel metal2 1978 1520 1978 1520 0 chany_top_out[5]
rlabel metal2 1794 8755 1794 8755 0 chany_top_out[6]
rlabel metal2 21942 38226 21942 38226 0 chany_top_out[7]
rlabel metal2 18078 1520 18078 1520 0 chany_top_out[8]
rlabel metal1 36156 37094 36156 37094 0 chany_top_out[9]
rlabel metal2 6210 29750 6210 29750 0 clknet_0_prog_clk
rlabel metal2 2622 17952 2622 17952 0 clknet_4_0_0_prog_clk
rlabel metal1 1840 33490 1840 33490 0 clknet_4_10_0_prog_clk
rlabel metal1 7728 31246 7728 31246 0 clknet_4_11_0_prog_clk
rlabel metal2 9154 29376 9154 29376 0 clknet_4_12_0_prog_clk
rlabel metal1 15180 32198 15180 32198 0 clknet_4_13_0_prog_clk
rlabel metal1 10626 30770 10626 30770 0 clknet_4_14_0_prog_clk
rlabel metal1 16698 35666 16698 35666 0 clknet_4_15_0_prog_clk
rlabel metal1 9246 22542 9246 22542 0 clknet_4_1_0_prog_clk
rlabel metal1 2852 24242 2852 24242 0 clknet_4_2_0_prog_clk
rlabel metal2 6762 25568 6762 25568 0 clknet_4_3_0_prog_clk
rlabel metal1 9936 23086 9936 23086 0 clknet_4_4_0_prog_clk
rlabel metal2 12926 17952 12926 17952 0 clknet_4_5_0_prog_clk
rlabel metal2 11822 24548 11822 24548 0 clknet_4_6_0_prog_clk
rlabel metal2 15502 22916 15502 22916 0 clknet_4_7_0_prog_clk
rlabel metal2 4922 28016 4922 28016 0 clknet_4_8_0_prog_clk
rlabel metal1 6256 30770 6256 30770 0 clknet_4_9_0_prog_clk
rlabel metal2 23782 12308 23782 12308 0 mem_bottom_track_1.DFFR_0_.D
rlabel metal2 20746 21250 20746 21250 0 mem_bottom_track_1.DFFR_0_.Q
rlabel metal2 15962 16592 15962 16592 0 mem_bottom_track_1.DFFR_1_.Q
rlabel metal1 11822 23188 11822 23188 0 mem_bottom_track_1.DFFR_2_.Q
rlabel metal2 12282 24616 12282 24616 0 mem_bottom_track_1.DFFR_3_.Q
rlabel metal2 11546 22304 11546 22304 0 mem_bottom_track_1.DFFR_4_.Q
rlabel metal1 11868 22134 11868 22134 0 mem_bottom_track_1.DFFR_5_.Q
rlabel metal1 9752 19414 9752 19414 0 mem_bottom_track_1.DFFR_6_.Q
rlabel metal1 11362 19482 11362 19482 0 mem_bottom_track_1.DFFR_7_.Q
rlabel metal2 21114 33660 21114 33660 0 mem_bottom_track_17.DFFR_0_.D
rlabel metal1 3496 31382 3496 31382 0 mem_bottom_track_17.DFFR_0_.Q
rlabel metal1 3995 28934 3995 28934 0 mem_bottom_track_17.DFFR_1_.Q
rlabel metal2 7038 27778 7038 27778 0 mem_bottom_track_17.DFFR_2_.Q
rlabel metal2 3542 27268 3542 27268 0 mem_bottom_track_17.DFFR_3_.Q
rlabel metal1 4462 27982 4462 27982 0 mem_bottom_track_17.DFFR_4_.Q
rlabel metal1 1564 24106 1564 24106 0 mem_bottom_track_17.DFFR_5_.Q
rlabel metal1 2024 23018 2024 23018 0 mem_bottom_track_17.DFFR_6_.Q
rlabel metal1 4324 28458 4324 28458 0 mem_bottom_track_17.DFFR_7_.Q
rlabel metal1 8096 28594 8096 28594 0 mem_bottom_track_25.DFFR_0_.Q
rlabel metal2 21896 35020 21896 35020 0 mem_bottom_track_25.DFFR_1_.Q
rlabel via2 9246 34901 9246 34901 0 mem_bottom_track_25.DFFR_2_.Q
rlabel metal1 8740 16218 8740 16218 0 mem_bottom_track_25.DFFR_3_.Q
rlabel metal2 14766 32776 14766 32776 0 mem_bottom_track_25.DFFR_4_.Q
rlabel metal1 17204 30158 17204 30158 0 mem_bottom_track_25.DFFR_5_.Q
rlabel metal2 18630 29886 18630 29886 0 mem_bottom_track_25.DFFR_6_.Q
rlabel metal1 16921 26554 16921 26554 0 mem_bottom_track_25.DFFR_7_.Q
rlabel metal1 14490 7378 14490 7378 0 mem_bottom_track_33.DFFR_0_.Q
rlabel metal1 17066 6290 17066 6290 0 mem_bottom_track_33.DFFR_1_.Q
rlabel metal1 10672 25330 10672 25330 0 mem_bottom_track_33.DFFR_2_.Q
rlabel metal2 10902 25602 10902 25602 0 mem_bottom_track_33.DFFR_3_.Q
rlabel metal2 13478 27676 13478 27676 0 mem_bottom_track_33.DFFR_4_.Q
rlabel metal1 10350 22746 10350 22746 0 mem_bottom_track_9.DFFR_0_.Q
rlabel metal2 11914 25466 11914 25466 0 mem_bottom_track_9.DFFR_1_.Q
rlabel metal2 20102 28849 20102 28849 0 mem_bottom_track_9.DFFR_2_.Q
rlabel metal1 27278 20468 27278 20468 0 mem_bottom_track_9.DFFR_3_.Q
rlabel metal1 21850 27064 21850 27064 0 mem_bottom_track_9.DFFR_4_.Q
rlabel metal1 8418 32810 8418 32810 0 mem_bottom_track_9.DFFR_5_.Q
rlabel metal2 9706 35394 9706 35394 0 mem_bottom_track_9.DFFR_6_.Q
rlabel metal1 6210 23494 6210 23494 0 mem_right_track_0.DFFR_0_.D
rlabel metal2 12466 18394 12466 18394 0 mem_right_track_0.DFFR_0_.Q
rlabel metal1 6762 20978 6762 20978 0 mem_right_track_0.DFFR_1_.Q
rlabel metal1 4094 18802 4094 18802 0 mem_right_track_0.DFFR_2_.Q
rlabel metal1 4922 20230 4922 20230 0 mem_right_track_0.DFFR_3_.Q
rlabel metal1 1886 17544 1886 17544 0 mem_right_track_0.DFFR_4_.Q
rlabel metal1 3450 17510 3450 17510 0 mem_right_track_0.DFFR_5_.Q
rlabel metal2 15778 23970 15778 23970 0 mem_right_track_10.DFFR_0_.D
rlabel metal1 22724 6766 22724 6766 0 mem_right_track_10.DFFR_0_.Q
rlabel metal1 12052 19754 12052 19754 0 mem_right_track_10.DFFR_1_.Q
rlabel metal1 10304 25806 10304 25806 0 mem_right_track_12.DFFR_0_.Q
rlabel metal2 11040 28900 11040 28900 0 mem_right_track_12.DFFR_1_.Q
rlabel metal1 11270 29070 11270 29070 0 mem_right_track_14.DFFR_0_.Q
rlabel metal2 4186 35802 4186 35802 0 mem_right_track_14.DFFR_1_.Q
rlabel metal3 17618 28900 17618 28900 0 mem_right_track_16.DFFR_0_.Q
rlabel metal2 8694 35020 8694 35020 0 mem_right_track_16.DFFR_1_.Q
rlabel metal1 19458 31926 19458 31926 0 mem_right_track_18.DFFR_0_.Q
rlabel metal1 16652 27982 16652 27982 0 mem_right_track_18.DFFR_1_.Q
rlabel metal1 14444 11730 14444 11730 0 mem_right_track_2.DFFR_0_.Q
rlabel metal1 25530 10778 25530 10778 0 mem_right_track_2.DFFR_1_.Q
rlabel metal1 7222 18666 7222 18666 0 mem_right_track_2.DFFR_2_.Q
rlabel metal1 5612 27370 5612 27370 0 mem_right_track_2.DFFR_3_.Q
rlabel metal1 8326 27574 8326 27574 0 mem_right_track_2.DFFR_4_.Q
rlabel metal1 10350 28186 10350 28186 0 mem_right_track_2.DFFR_5_.Q
rlabel metal1 23782 8976 23782 8976 0 mem_right_track_20.DFFR_0_.Q
rlabel metal1 21390 10098 21390 10098 0 mem_right_track_20.DFFR_1_.Q
rlabel metal1 15180 18190 15180 18190 0 mem_right_track_22.DFFR_0_.Q
rlabel metal1 16744 17714 16744 17714 0 mem_right_track_22.DFFR_1_.Q
rlabel metal1 18906 9996 18906 9996 0 mem_right_track_24.DFFR_0_.Q
rlabel metal1 16376 19142 16376 19142 0 mem_right_track_24.DFFR_1_.Q
rlabel metal1 17158 11730 17158 11730 0 mem_right_track_26.DFFR_0_.Q
rlabel metal1 8326 30566 8326 30566 0 mem_right_track_4.DFFR_0_.Q
rlabel metal1 2714 10064 2714 10064 0 mem_right_track_4.DFFR_1_.Q
rlabel metal2 1380 19244 1380 19244 0 mem_right_track_4.DFFR_2_.Q
rlabel metal1 8694 22576 8694 22576 0 mem_right_track_4.DFFR_3_.Q
rlabel metal1 12045 28934 12045 28934 0 mem_right_track_4.DFFR_4_.Q
rlabel metal2 9430 29410 9430 29410 0 mem_right_track_4.DFFR_5_.Q
rlabel metal1 6578 34442 6578 34442 0 mem_right_track_6.DFFR_0_.Q
rlabel metal2 5014 35224 5014 35224 0 mem_right_track_6.DFFR_1_.Q
rlabel via3 5405 22100 5405 22100 0 mem_right_track_6.DFFR_2_.Q
rlabel via2 5934 33915 5934 33915 0 mem_right_track_6.DFFR_3_.Q
rlabel metal1 14582 32300 14582 32300 0 mem_right_track_6.DFFR_4_.Q
rlabel metal1 16100 34986 16100 34986 0 mem_right_track_6.DFFR_5_.Q
rlabel metal1 17526 32334 17526 32334 0 mem_right_track_8.DFFR_0_.Q
rlabel metal1 6164 24174 6164 24174 0 mem_top_track_0.DFFR_0_.Q
rlabel metal2 16146 35615 16146 35615 0 mem_top_track_0.DFFR_1_.Q
rlabel metal1 21022 22610 21022 22610 0 mem_top_track_0.DFFR_2_.Q
rlabel metal1 15732 32810 15732 32810 0 mem_top_track_0.DFFR_3_.Q
rlabel metal1 17388 33422 17388 33422 0 mem_top_track_0.DFFR_4_.Q
rlabel metal1 18584 33286 18584 33286 0 mem_top_track_0.DFFR_5_.Q
rlabel metal2 17618 31620 17618 31620 0 mem_top_track_0.DFFR_6_.Q
rlabel metal2 17158 25993 17158 25993 0 mem_top_track_0.DFFR_7_.Q
rlabel via2 6026 22389 6026 22389 0 mem_top_track_16.DFFR_0_.D
rlabel metal1 9200 23630 9200 23630 0 mem_top_track_16.DFFR_0_.Q
rlabel metal1 2530 8976 2530 8976 0 mem_top_track_16.DFFR_1_.Q
rlabel via1 7859 30022 7859 30022 0 mem_top_track_16.DFFR_2_.Q
rlabel metal2 9338 29342 9338 29342 0 mem_top_track_16.DFFR_3_.Q
rlabel metal2 9890 22644 9890 22644 0 mem_top_track_16.DFFR_4_.Q
rlabel metal1 8602 25126 8602 25126 0 mem_top_track_16.DFFR_5_.Q
rlabel metal1 6164 19754 6164 19754 0 mem_top_track_16.DFFR_6_.Q
rlabel metal1 9374 27642 9374 27642 0 mem_top_track_16.DFFR_7_.Q
rlabel metal1 12098 27506 12098 27506 0 mem_top_track_24.DFFR_0_.Q
rlabel metal1 11822 31246 11822 31246 0 mem_top_track_24.DFFR_1_.Q
rlabel metal1 14306 31382 14306 31382 0 mem_top_track_24.DFFR_2_.Q
rlabel metal1 23230 35564 23230 35564 0 mem_top_track_24.DFFR_3_.Q
rlabel metal2 18630 34680 18630 34680 0 mem_top_track_24.DFFR_4_.Q
rlabel metal1 18768 35462 18768 35462 0 mem_top_track_24.DFFR_5_.Q
rlabel metal1 21206 33388 21206 33388 0 mem_top_track_32.DFFR_0_.Q
rlabel metal1 11086 32810 11086 32810 0 mem_top_track_32.DFFR_1_.Q
rlabel metal1 4876 30770 4876 30770 0 mem_top_track_32.DFFR_2_.Q
rlabel metal1 2530 13260 2530 13260 0 mem_top_track_32.DFFR_3_.Q
rlabel metal1 4646 23766 4646 23766 0 mem_top_track_32.DFFR_4_.Q
rlabel metal2 18630 25398 18630 25398 0 mem_top_track_8.DFFR_0_.Q
rlabel metal1 15686 24072 15686 24072 0 mem_top_track_8.DFFR_1_.Q
rlabel metal1 17480 20774 17480 20774 0 mem_top_track_8.DFFR_2_.Q
rlabel metal1 10626 23222 10626 23222 0 mem_top_track_8.DFFR_3_.Q
rlabel metal1 7544 22950 7544 22950 0 mem_top_track_8.DFFR_4_.Q
rlabel metal1 6847 22202 6847 22202 0 mem_top_track_8.DFFR_5_.Q
rlabel metal1 5704 22542 5704 22542 0 mem_top_track_8.DFFR_6_.Q
rlabel metal1 20976 14926 20976 14926 0 mux_bottom_track_1.INVTX1_0_.out
rlabel metal2 23414 12308 23414 12308 0 mux_bottom_track_1.INVTX1_1_.out
rlabel metal1 18906 9690 18906 9690 0 mux_bottom_track_1.INVTX1_2_.out
rlabel metal1 26956 14450 26956 14450 0 mux_bottom_track_1.INVTX1_3_.out
rlabel metal1 12834 36618 12834 36618 0 mux_bottom_track_1.INVTX1_4_.out
rlabel metal2 24702 21454 24702 21454 0 mux_bottom_track_1.INVTX1_5_.out
rlabel metal1 6762 10710 6762 10710 0 mux_bottom_track_1.INVTX1_6_.out
rlabel metal1 23736 32334 23736 32334 0 mux_bottom_track_1.INVTX1_7_.out
rlabel metal1 18630 4046 18630 4046 0 mux_bottom_track_1.INVTX1_8_.out
rlabel metal2 19366 12852 19366 12852 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 14766 13192 14766 13192 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 19642 5134 19642 5134 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 21942 3706 21942 3706 0 mux_bottom_track_1.out
rlabel metal1 8372 13430 8372 13430 0 mux_bottom_track_17.INVTX1_0_.out
rlabel metal2 20194 17527 20194 17527 0 mux_bottom_track_17.INVTX1_1_.out
rlabel metal1 18676 10098 18676 10098 0 mux_bottom_track_17.INVTX1_2_.out
rlabel metal1 19642 6630 19642 6630 0 mux_bottom_track_17.INVTX1_3_.out
rlabel metal2 27278 32946 27278 32946 0 mux_bottom_track_17.INVTX1_4_.out
rlabel metal1 6440 9078 6440 9078 0 mux_bottom_track_17.INVTX1_5_.out
rlabel metal1 25806 32198 25806 32198 0 mux_bottom_track_17.INVTX1_6_.out
rlabel metal2 2162 27404 2162 27404 0 mux_bottom_track_17.INVTX1_7_.out
rlabel metal1 2116 14042 2116 14042 0 mux_bottom_track_17.INVTX1_8_.out
rlabel metal1 2323 14926 2323 14926 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 1794 10540 1794 10540 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 2484 10574 2484 10574 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 2254 5610 2254 5610 0 mux_bottom_track_17.out
rlabel metal2 18262 29138 18262 29138 0 mux_bottom_track_25.INVTX1_0_.out
rlabel metal1 21344 27098 21344 27098 0 mux_bottom_track_25.INVTX1_1_.out
rlabel metal2 21022 23545 21022 23545 0 mux_bottom_track_25.INVTX1_2_.out
rlabel metal1 2990 15980 2990 15980 0 mux_bottom_track_25.INVTX1_3_.out
rlabel metal1 27416 11322 27416 11322 0 mux_bottom_track_25.INVTX1_4_.out
rlabel metal1 27830 36686 27830 36686 0 mux_bottom_track_25.INVTX1_5_.out
rlabel metal2 14030 36023 14030 36023 0 mux_bottom_track_25.INVTX1_6_.out
rlabel metal2 12742 36482 12742 36482 0 mux_bottom_track_25.INVTX1_7_.out
rlabel metal1 31510 28526 31510 28526 0 mux_bottom_track_25.INVTX1_8_.out
rlabel metal2 17250 24140 17250 24140 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 25576 35598 25576 35598 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 21022 26792 21022 26792 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 36478 8636 36478 8636 0 mux_bottom_track_25.out
rlabel metal2 29762 16388 29762 16388 0 mux_bottom_track_33.INVTX1_0_.out
rlabel metal2 27278 26894 27278 26894 0 mux_bottom_track_33.INVTX1_1_.out
rlabel via2 21942 27523 21942 27523 0 mux_bottom_track_33.INVTX1_2_.out
rlabel metal1 13616 6834 13616 6834 0 mux_bottom_track_33.INVTX1_3_.out
rlabel metal1 19872 7310 19872 7310 0 mux_bottom_track_33.INVTX1_4_.out
rlabel metal1 11868 6426 11868 6426 0 mux_bottom_track_33.INVTX1_5_.out
rlabel metal2 14398 6324 14398 6324 0 mux_bottom_track_33.INVTX1_6_.out
rlabel metal1 18124 6834 18124 6834 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem2_0_out
rlabel metal1 18676 27370 18676 27370 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 20102 7548 20102 7548 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 19228 7446 19228 7446 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 6762 6732 6762 6732 0 mux_bottom_track_33.out
rlabel metal1 15364 12274 15364 12274 0 mux_bottom_track_9.INVTX1_0_.out
rlabel metal1 28244 21114 28244 21114 0 mux_bottom_track_9.INVTX1_1_.out
rlabel metal1 19918 17714 19918 17714 0 mux_bottom_track_9.INVTX1_2_.out
rlabel metal2 27462 20604 27462 20604 0 mux_bottom_track_9.INVTX1_3_.out
rlabel metal2 20562 9554 20562 9554 0 mux_bottom_track_9.INVTX1_4_.out
rlabel metal1 21390 29104 21390 29104 0 mux_bottom_track_9.INVTX1_5_.out
rlabel metal1 26588 28594 26588 28594 0 mux_bottom_track_9.INVTX1_6_.out
rlabel metal1 30590 14042 30590 14042 0 mux_bottom_track_9.INVTX1_7_.out
rlabel via2 2438 31773 2438 31773 0 mux_bottom_track_9.INVTX1_8_.out
rlabel metal1 17986 17816 17986 17816 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 22954 12342 22954 12342 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 35098 36686 35098 36686 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 35558 36754 35558 36754 0 mux_bottom_track_9.out
rlabel metal2 24702 16184 24702 16184 0 mux_right_track_0.INVTX1_1_.out
rlabel metal2 7958 10268 7958 10268 0 mux_right_track_0.INVTX1_2_.out
rlabel metal2 21298 15334 21298 15334 0 mux_right_track_0.INVTX1_3_.out
rlabel metal2 20194 14484 20194 14484 0 mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 4002 13328 4002 13328 0 mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 4094 16116 4094 16116 0 mux_right_track_0.out
rlabel metal1 25300 6426 25300 6426 0 mux_right_track_10.INVTX1_1_.out
rlabel metal1 17618 8874 17618 8874 0 mux_right_track_10.INVTX1_2_.out
rlabel metal2 23506 8704 23506 8704 0 mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 13570 8296 13570 8296 0 mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 12466 8092 12466 8092 0 mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 8602 6766 8602 6766 0 mux_right_track_10.out
rlabel metal2 25622 24174 25622 24174 0 mux_right_track_12.INVTX1_1_.out
rlabel metal1 29854 20876 29854 20876 0 mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 31832 20434 31832 20434 0 mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 33350 18802 33350 18802 0 mux_right_track_12.out
rlabel metal1 21390 32946 21390 32946 0 mux_right_track_14.INVTX1_1_.out
rlabel metal1 22816 34986 22816 34986 0 mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 5888 36210 5888 36210 0 mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 2300 33082 2300 33082 0 mux_right_track_14.out
rlabel metal1 22816 27914 22816 27914 0 mux_right_track_16.INVTX1_1_.out
rlabel metal1 22954 35734 22954 35734 0 mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 14214 34952 14214 34952 0 mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 5934 35904 5934 35904 0 mux_right_track_16.out
rlabel metal1 27002 32334 27002 32334 0 mux_right_track_18.INVTX1_2_.out
rlabel metal2 28474 26146 28474 26146 0 mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 28152 32198 28152 32198 0 mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 28566 30192 28566 30192 0 mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 32982 29614 32982 29614 0 mux_right_track_18.out
rlabel metal2 24334 9860 24334 9860 0 mux_right_track_2.INVTX1_1_.out
rlabel metal1 2162 15572 2162 15572 0 mux_right_track_2.INVTX1_3_.out
rlabel metal2 26542 15266 26542 15266 0 mux_right_track_2.INVTX1_4_.out
rlabel metal2 21390 14535 21390 14535 0 mux_right_track_2.mux_2level_tapbuf_basis_input2_mem2_0_out
rlabel metal2 19274 11152 19274 11152 0 mux_right_track_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 20746 17680 20746 17680 0 mux_right_track_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 14858 36448 14858 36448 0 mux_right_track_2.out
rlabel metal1 29624 18394 29624 18394 0 mux_right_track_20.INVTX1_2_.out
rlabel metal2 19826 9248 19826 9248 0 mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 25438 11118 25438 11118 0 mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 25300 6290 25300 6290 0 mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 25714 5882 25714 5882 0 mux_right_track_20.out
rlabel metal2 22402 15062 22402 15062 0 mux_right_track_22.INVTX1_2_.out
rlabel metal2 20746 15504 20746 15504 0 mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 26358 16728 26358 16728 0 mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 27922 14654 27922 14654 0 mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 32522 12988 32522 12988 0 mux_right_track_22.out
rlabel metal1 17089 10030 17089 10030 0 mux_right_track_24.INVTX1_1_.out
rlabel metal2 17710 10982 17710 10982 0 mux_right_track_24.INVTX1_2_.out
rlabel metal1 21850 10234 21850 10234 0 mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 26496 11322 26496 11322 0 mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 29026 12274 29026 12274 0 mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 31326 19482 31326 19482 0 mux_right_track_24.out
rlabel metal1 17894 13226 17894 13226 0 mux_right_track_26.INVTX1_1_.out
rlabel metal1 27462 9554 27462 9554 0 mux_right_track_26.INVTX1_2_.out
rlabel metal1 20792 13226 20792 13226 0 mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 26358 10064 26358 10064 0 mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 25622 10540 25622 10540 0 mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 32246 3502 32246 3502 0 mux_right_track_26.out
rlabel metal1 2070 8534 2070 8534 0 mux_right_track_4.INVTX1_1_.out
rlabel metal1 3312 13838 3312 13838 0 mux_right_track_4.INVTX1_4_.out
rlabel metal1 8740 14586 8740 14586 0 mux_right_track_4.mux_2level_tapbuf_basis_input2_mem2_0_out
rlabel metal1 2392 15538 2392 15538 0 mux_right_track_4.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 12926 14620 12926 14620 0 mux_right_track_4.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 30590 22066 30590 22066 0 mux_right_track_4.out
rlabel metal1 8372 36686 8372 36686 0 mux_right_track_6.INVTX1_1_.out
rlabel metal2 19918 32266 19918 32266 0 mux_right_track_6.INVTX1_3_.out
rlabel metal2 8694 26220 8694 26220 0 mux_right_track_6.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 21850 36074 21850 36074 0 mux_right_track_6.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 26312 36346 26312 36346 0 mux_right_track_6.out
rlabel metal1 27416 8602 27416 8602 0 mux_right_track_8.INVTX1_1_.out
rlabel metal2 20930 29920 20930 29920 0 mux_right_track_8.INVTX1_2_.out
rlabel metal1 30452 16558 30452 16558 0 mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 27784 32266 27784 32266 0 mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 31878 26044 31878 26044 0 mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 31970 26758 31970 26758 0 mux_right_track_8.out
rlabel metal1 28290 26894 28290 26894 0 mux_top_track_0.INVTX1_0_.out
rlabel metal2 20930 34833 20930 34833 0 mux_top_track_0.INVTX1_1_.out
rlabel metal2 27922 33966 27922 33966 0 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 20332 18666 20332 18666 0 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 33258 24990 33258 24990 0 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 34454 23052 34454 23052 0 mux_top_track_0.out
rlabel metal1 28428 32946 28428 32946 0 mux_top_track_16.INVTX1_0_.out
rlabel metal2 3818 10880 3818 10880 0 mux_top_track_16.INVTX1_1_.out
rlabel metal1 15962 14824 15962 14824 0 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 15870 14688 15870 14688 0 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 13892 11254 13892 11254 0 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 15686 8092 15686 8092 0 mux_top_track_16.out
rlabel metal2 26358 35292 26358 35292 0 mux_top_track_24.INVTX1_0_.out
rlabel metal2 27278 34119 27278 34119 0 mux_top_track_24.INVTX1_1_.out
rlabel metal1 24610 34646 24610 34646 0 mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 20148 9554 20148 9554 0 mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 20194 23664 20194 23664 0 mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 23322 31892 23322 31892 0 mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 35282 34986 35282 34986 0 mux_top_track_24.out
rlabel metal1 6394 36244 6394 36244 0 mux_top_track_32.INVTX1_0_.out
rlabel metal1 28428 23834 28428 23834 0 mux_top_track_32.INVTX1_1_.out
rlabel metal2 17250 16898 17250 16898 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 23506 34476 23506 34476 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 9246 16796 9246 16796 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 1978 16830 1978 16830 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 3266 6970 3266 6970 0 mux_top_track_32.out
rlabel metal1 21850 7514 21850 7514 0 mux_top_track_8.INVTX1_0_.out
rlabel metal1 26680 7922 26680 7922 0 mux_top_track_8.INVTX1_1_.out
rlabel metal1 23138 7786 23138 7786 0 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 27278 15538 27278 15538 0 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 19320 11050 19320 11050 0 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 6762 3468 6762 3468 0 mux_top_track_8.out
rlabel metal2 1886 28730 1886 28730 0 net1
rlabel metal1 37536 8602 37536 8602 0 net10
rlabel metal1 36961 18258 36961 18258 0 net100
rlabel metal1 1748 31790 1748 31790 0 net101
rlabel metal1 2162 35054 2162 35054 0 net102
rlabel metal1 36754 32402 36754 32402 0 net103
rlabel metal1 22218 3366 22218 3366 0 net104
rlabel metal1 13478 14246 13478 14246 0 net105
rlabel metal2 29118 25262 29118 25262 0 net106
rlabel metal1 37168 8330 37168 8330 0 net107
rlabel metal1 27002 36890 27002 36890 0 net108
rlabel metal2 37306 25738 37306 25738 0 net109
rlabel metal3 4715 23596 4715 23596 0 net11
rlabel metal2 21206 36414 21206 36414 0 net110
rlabel metal1 1610 3060 1610 3060 0 net111
rlabel metal2 5290 2244 5290 2244 0 net112
rlabel metal1 21206 37196 21206 37196 0 net113
rlabel metal1 8510 26282 8510 26282 0 net114
rlabel metal1 37950 21522 37950 21522 0 net115
rlabel metal1 36961 14382 36961 14382 0 net116
rlabel metal1 36662 36788 36662 36788 0 net117
rlabel metal1 3634 2414 3634 2414 0 net118
rlabel metal1 37996 3502 37996 3502 0 net119
rlabel metal2 2162 18462 2162 18462 0 net12
rlabel metal2 36938 15606 36938 15606 0 net120
rlabel metal2 2070 5865 2070 5865 0 net121
rlabel metal2 8050 27744 8050 27744 0 net122
rlabel metal1 38042 22576 38042 22576 0 net123
rlabel metal2 36662 34374 36662 34374 0 net124
rlabel metal1 36041 2414 36041 2414 0 net125
rlabel metal1 37306 36074 37306 36074 0 net126
rlabel metal2 2438 34017 2438 34017 0 net127
rlabel metal1 2070 3502 2070 3502 0 net128
rlabel metal1 1610 12172 1610 12172 0 net129
rlabel metal1 29578 36720 29578 36720 0 net13
rlabel metal2 3082 4828 3082 4828 0 net130
rlabel metal1 21896 8330 21896 8330 0 net131
rlabel metal3 1863 36380 1863 36380 0 net132
rlabel metal2 10028 22780 10028 22780 0 net133
rlabel metal1 24242 20774 24242 20774 0 net134
rlabel via3 1955 6460 1955 6460 0 net135
rlabel metal2 6578 2618 6578 2618 0 net136
rlabel metal1 4370 2448 4370 2448 0 net137
rlabel metal1 1656 23494 1656 23494 0 net138
rlabel metal1 21804 36754 21804 36754 0 net139
rlabel metal1 2576 23494 2576 23494 0 net14
rlabel metal1 18032 2414 18032 2414 0 net140
rlabel metal2 36202 31212 36202 31212 0 net141
rlabel metal1 32660 26010 32660 26010 0 net142
rlabel metal2 2990 7922 2990 7922 0 net143
rlabel metal2 10718 11424 10718 11424 0 net144
rlabel metal1 15502 10098 15502 10098 0 net145
rlabel metal1 28290 34714 28290 34714 0 net146
rlabel metal1 3174 11662 3174 11662 0 net147
rlabel metal2 29854 23392 29854 23392 0 net148
rlabel metal2 18170 23902 18170 23902 0 net149
rlabel metal2 12834 36737 12834 36737 0 net15
rlabel metal2 20470 33694 20470 33694 0 net150
rlabel metal2 2346 10914 2346 10914 0 net151
rlabel metal2 25530 36652 25530 36652 0 net152
rlabel metal1 17434 31246 17434 31246 0 net153
rlabel metal1 21206 21658 21206 21658 0 net154
rlabel metal2 28566 24480 28566 24480 0 net155
rlabel metal2 12926 7548 12926 7548 0 net156
rlabel metal1 27830 31314 27830 31314 0 net157
rlabel metal2 28198 11424 28198 11424 0 net158
rlabel metal1 25668 17102 25668 17102 0 net159
rlabel metal1 37628 11322 37628 11322 0 net16
rlabel metal2 25806 11424 25806 11424 0 net160
rlabel metal2 25714 9724 25714 9724 0 net161
rlabel metal1 31234 19890 31234 19890 0 net162
rlabel metal2 4830 36448 4830 36448 0 net163
rlabel metal2 9246 35564 9246 35564 0 net164
rlabel metal1 17388 6834 17388 6834 0 net165
rlabel metal1 24564 7854 24564 7854 0 net17
rlabel metal2 13938 35836 13938 35836 0 net18
rlabel metal1 35374 36006 35374 36006 0 net19
rlabel metal1 12282 36720 12282 36720 0 net2
rlabel metal2 37490 32334 37490 32334 0 net20
rlabel metal2 6578 7990 6578 7990 0 net21
rlabel metal2 20746 4692 20746 4692 0 net22
rlabel metal1 37030 27846 37030 27846 0 net23
rlabel metal1 34937 12682 34937 12682 0 net24
rlabel metal1 18446 36856 18446 36856 0 net25
rlabel metal1 37766 2924 37766 2924 0 net26
rlabel metal2 33074 36686 33074 36686 0 net27
rlabel metal1 18492 7854 18492 7854 0 net28
rlabel metal1 10626 36754 10626 36754 0 net29
rlabel metal2 13018 4454 13018 4454 0 net3
rlabel metal1 11684 2550 11684 2550 0 net30
rlabel metal1 30038 3978 30038 3978 0 net31
rlabel metal1 22586 37230 22586 37230 0 net32
rlabel via2 15410 36805 15410 36805 0 net33
rlabel metal1 28842 32402 28842 32402 0 net34
rlabel metal1 38134 37298 38134 37298 0 net35
rlabel metal2 21942 12546 21942 12546 0 net36
rlabel metal1 13202 3060 13202 3060 0 net37
rlabel metal2 1886 16354 1886 16354 0 net38
rlabel metal2 1610 8194 1610 8194 0 net39
rlabel metal2 19458 3366 19458 3366 0 net4
rlabel metal1 28980 5678 28980 5678 0 net40
rlabel metal1 36156 3162 36156 3162 0 net41
rlabel metal2 3266 15130 3266 15130 0 net42
rlabel metal1 37260 7718 37260 7718 0 net43
rlabel metal4 20700 35156 20700 35156 0 net44
rlabel metal1 4416 24582 4416 24582 0 net45
rlabel metal1 19964 19346 19964 19346 0 net46
rlabel metal2 16882 5712 16882 5712 0 net47
rlabel metal1 6578 24276 6578 24276 0 net48
rlabel metal2 36846 35564 36846 35564 0 net49
rlabel metal1 1978 27098 1978 27098 0 net5
rlabel metal2 37766 7854 37766 7854 0 net50
rlabel metal1 14398 20876 14398 20876 0 net51
rlabel metal1 2346 36856 2346 36856 0 net52
rlabel metal2 38226 36414 38226 36414 0 net53
rlabel metal1 18814 9554 18814 9554 0 net54
rlabel metal1 18170 18088 18170 18088 0 net55
rlabel metal1 26726 8466 26726 8466 0 net56
rlabel metal2 37490 3230 37490 3230 0 net57
rlabel metal1 14674 35190 14674 35190 0 net58
rlabel metal1 26726 6290 26726 6290 0 net59
rlabel metal1 1518 6630 1518 6630 0 net6
rlabel metal1 4278 2516 4278 2516 0 net60
rlabel metal2 31970 13906 31970 13906 0 net61
rlabel metal1 37674 4794 37674 4794 0 net62
rlabel metal2 34638 28356 34638 28356 0 net63
rlabel metal1 37904 14994 37904 14994 0 net64
rlabel metal1 33902 2550 33902 2550 0 net65
rlabel metal1 1426 24582 1426 24582 0 net66
rlabel metal1 33212 10098 33212 10098 0 net67
rlabel metal1 2070 32266 2070 32266 0 net68
rlabel metal1 32798 6086 32798 6086 0 net69
rlabel metal2 38134 29580 38134 29580 0 net7
rlabel metal1 3680 11866 3680 11866 0 net70
rlabel metal1 6578 10030 6578 10030 0 net71
rlabel metal1 19550 2890 19550 2890 0 net72
rlabel metal2 5658 6766 5658 6766 0 net73
rlabel metal2 38134 26724 38134 26724 0 net74
rlabel metal2 22034 4998 22034 4998 0 net75
rlabel metal1 29026 33524 29026 33524 0 net76
rlabel metal1 26450 35632 26450 35632 0 net77
rlabel metal2 2990 36550 2990 36550 0 net78
rlabel metal1 13570 36822 13570 36822 0 net79
rlabel metal1 12144 2618 12144 2618 0 net8
rlabel metal1 27278 2618 27278 2618 0 net80
rlabel metal2 3726 9724 3726 9724 0 net81
rlabel metal1 5566 34646 5566 34646 0 net82
rlabel metal2 38134 20264 38134 20264 0 net83
rlabel metal1 18170 20910 18170 20910 0 net84
rlabel metal1 1610 16150 1610 16150 0 net85
rlabel metal1 25392 5542 25392 5542 0 net86
rlabel metal2 32338 13124 32338 13124 0 net87
rlabel metal2 38042 24548 38042 24548 0 net88
rlabel metal1 34362 2414 34362 2414 0 net89
rlabel metal1 24426 33524 24426 33524 0 net9
rlabel metal2 14950 2618 14950 2618 0 net90
rlabel metal1 32338 37196 32338 37196 0 net91
rlabel metal2 15962 8959 15962 8959 0 net92
rlabel metal2 34822 3196 34822 3196 0 net93
rlabel metal2 38042 16218 38042 16218 0 net94
rlabel metal2 20746 36567 20746 36567 0 net95
rlabel metal2 34730 23460 34730 23460 0 net96
rlabel metal2 21114 37264 21114 37264 0 net97
rlabel metal1 36110 32878 36110 32878 0 net98
rlabel metal2 6670 5610 6670 5610 0 net99
rlabel metal2 38318 6239 38318 6239 0 pReset
rlabel metal1 9430 27064 9430 27064 0 prog_clk
rlabel metal2 3634 11679 3634 11679 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal2 7130 1588 7130 1588 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal2 14214 1894 14214 1894 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
rlabel metal3 1050 3468 1050 3468 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
rlabel metal2 38318 26129 38318 26129 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 21942 1588 21942 1588 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 30406 37230 30406 37230 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 29486 37230 29486 37230 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 1564 36142 1564 36142 0 top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal1 6624 37230 6624 37230 0 top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal2 27094 1588 27094 1588 0 top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal2 3450 10149 3450 10149 0 top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal3 1234 34748 1234 34748 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 38318 19227 38318 19227 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
