// This is the unpowered netlist.
module cby_0__1_ (ccff_head,
    ccff_tail,
    left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_,
    left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_,
    left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_,
    left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_,
    left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_,
    left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_,
    left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_,
    left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_,
    pReset,
    prog_clk,
    right_grid_left_width_0_height_0_subtile_0__pin_I_11_,
    right_grid_left_width_0_height_0_subtile_0__pin_I_3_,
    right_grid_left_width_0_height_0_subtile_0__pin_I_7_,
    chany_bottom_in,
    chany_bottom_out,
    chany_top_in,
    chany_top_out);
 input ccff_head;
 output ccff_tail;
 output left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
 output left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
 output left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
 output left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
 output left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
 output left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
 output left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
 output left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
 input pReset;
 input prog_clk;
 output right_grid_left_width_0_height_0_subtile_0__pin_I_11_;
 output right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
 output right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
 input [0:18] chany_bottom_in;
 output [0:18] chany_bottom_out;
 input [0:18] chany_top_in;
 output [0:18] chany_top_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire \mem_left_ipin_0.DFFR_0_.Q ;
 wire \mem_left_ipin_0.DFFR_1_.Q ;
 wire \mem_left_ipin_0.DFFR_2_.Q ;
 wire \mem_left_ipin_0.DFFR_3_.Q ;
 wire \mem_left_ipin_0.DFFR_4_.Q ;
 wire \mem_left_ipin_0.DFFR_5_.Q ;
 wire \mem_left_ipin_1.DFFR_0_.Q ;
 wire \mem_left_ipin_1.DFFR_1_.Q ;
 wire \mem_left_ipin_1.DFFR_2_.Q ;
 wire \mem_left_ipin_1.DFFR_3_.Q ;
 wire \mem_left_ipin_1.DFFR_4_.Q ;
 wire \mem_left_ipin_1.DFFR_5_.Q ;
 wire \mem_left_ipin_2.DFFR_0_.Q ;
 wire \mem_left_ipin_2.DFFR_1_.Q ;
 wire \mem_left_ipin_2.DFFR_2_.Q ;
 wire \mem_left_ipin_2.DFFR_3_.Q ;
 wire \mem_left_ipin_2.DFFR_4_.Q ;
 wire \mem_left_ipin_2.DFFR_5_.Q ;
 wire \mem_right_ipin_0.DFFR_0_.Q ;
 wire \mem_right_ipin_0.DFFR_1_.Q ;
 wire \mem_right_ipin_0.DFFR_2_.Q ;
 wire \mem_right_ipin_0.DFFR_3_.Q ;
 wire \mem_right_ipin_0.DFFR_4_.Q ;
 wire \mem_right_ipin_0.DFFR_5_.Q ;
 wire \mem_right_ipin_1.DFFR_0_.Q ;
 wire \mem_right_ipin_1.DFFR_1_.Q ;
 wire \mem_right_ipin_1.DFFR_2_.Q ;
 wire \mem_right_ipin_1.DFFR_3_.Q ;
 wire \mem_right_ipin_1.DFFR_4_.Q ;
 wire \mem_right_ipin_1.DFFR_5_.Q ;
 wire \mem_right_ipin_2.DFFR_0_.Q ;
 wire \mem_right_ipin_2.DFFR_1_.Q ;
 wire \mem_right_ipin_2.DFFR_2_.Q ;
 wire \mem_right_ipin_2.DFFR_3_.Q ;
 wire \mem_right_ipin_2.DFFR_4_.Q ;
 wire \mem_right_ipin_2.DFFR_5_.Q ;
 wire \mem_right_ipin_3.DFFR_0_.Q ;
 wire \mem_right_ipin_3.DFFR_1_.Q ;
 wire \mem_right_ipin_3.DFFR_2_.Q ;
 wire \mem_right_ipin_3.DFFR_3_.Q ;
 wire \mem_right_ipin_3.DFFR_4_.Q ;
 wire \mem_right_ipin_3.DFFR_5_.Q ;
 wire \mem_right_ipin_4.DFFR_0_.Q ;
 wire \mem_right_ipin_4.DFFR_1_.Q ;
 wire \mem_right_ipin_4.DFFR_2_.Q ;
 wire \mem_right_ipin_4.DFFR_3_.Q ;
 wire \mem_right_ipin_4.DFFR_4_.Q ;
 wire \mem_right_ipin_4.DFFR_5_.Q ;
 wire \mem_right_ipin_5.DFFR_0_.Q ;
 wire \mem_right_ipin_5.DFFR_1_.Q ;
 wire \mem_right_ipin_5.DFFR_2_.Q ;
 wire \mem_right_ipin_5.DFFR_3_.Q ;
 wire \mem_right_ipin_5.DFFR_4_.Q ;
 wire \mem_right_ipin_5.DFFR_5_.Q ;
 wire \mem_right_ipin_6.DFFR_0_.Q ;
 wire \mem_right_ipin_6.DFFR_1_.Q ;
 wire \mem_right_ipin_6.DFFR_2_.Q ;
 wire \mem_right_ipin_6.DFFR_3_.Q ;
 wire \mem_right_ipin_6.DFFR_4_.Q ;
 wire \mem_right_ipin_6.DFFR_5_.Q ;
 wire \mem_right_ipin_7.DFFR_0_.Q ;
 wire \mem_right_ipin_7.DFFR_1_.Q ;
 wire \mem_right_ipin_7.DFFR_2_.Q ;
 wire \mem_right_ipin_7.DFFR_3_.Q ;
 wire \mem_right_ipin_7.DFFR_4_.Q ;
 wire \mux_left_ipin_0.INVTX1_0_.out ;
 wire \mux_left_ipin_0.INVTX1_1_.out ;
 wire \mux_left_ipin_0.INVTX1_2_.out ;
 wire \mux_left_ipin_0.INVTX1_3_.out ;
 wire \mux_left_ipin_0.INVTX1_4_.out ;
 wire \mux_left_ipin_0.INVTX1_5_.out ;
 wire \mux_left_ipin_0.INVTX1_6_.out ;
 wire \mux_left_ipin_0.INVTX1_7_.out ;
 wire \mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_left_ipin_1.INVTX1_2_.out ;
 wire \mux_left_ipin_1.INVTX1_3_.out ;
 wire \mux_left_ipin_1.INVTX1_4_.out ;
 wire \mux_left_ipin_1.INVTX1_5_.out ;
 wire \mux_left_ipin_1.INVTX1_6_.out ;
 wire \mux_left_ipin_1.INVTX1_7_.out ;
 wire \mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_left_ipin_2.INVTX1_2_.out ;
 wire \mux_left_ipin_2.INVTX1_3_.out ;
 wire \mux_left_ipin_2.INVTX1_4_.out ;
 wire \mux_left_ipin_2.INVTX1_5_.out ;
 wire \mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_right_ipin_0.INVTX1_2_.out ;
 wire \mux_right_ipin_0.INVTX1_3_.out ;
 wire \mux_right_ipin_0.INVTX1_4_.out ;
 wire \mux_right_ipin_0.INVTX1_5_.out ;
 wire \mux_right_ipin_0.INVTX1_6_.out ;
 wire \mux_right_ipin_0.INVTX1_7_.out ;
 wire \mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_right_ipin_1.INVTX1_2_.out ;
 wire \mux_right_ipin_1.INVTX1_3_.out ;
 wire \mux_right_ipin_1.INVTX1_4_.out ;
 wire \mux_right_ipin_1.INVTX1_5_.out ;
 wire \mux_right_ipin_1.INVTX1_6_.out ;
 wire \mux_right_ipin_1.INVTX1_7_.out ;
 wire \mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_right_ipin_2.INVTX1_2_.out ;
 wire \mux_right_ipin_2.INVTX1_3_.out ;
 wire \mux_right_ipin_2.INVTX1_6_.out ;
 wire \mux_right_ipin_2.INVTX1_7_.out ;
 wire \mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_right_ipin_5.INVTX1_4_.out ;
 wire \mux_right_ipin_5.INVTX1_5_.out ;
 wire \mux_right_ipin_5.INVTX1_6_.out ;
 wire \mux_right_ipin_5.INVTX1_7_.out ;
 wire \mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire \mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out ;
 wire \mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out ;
 wire \mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out ;
 wire \mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;

 sky130_fd_sc_hd__inv_2 _213_ (.A(\mem_left_ipin_2.DFFR_3_.Q ),
    .Y(_199_));
 sky130_fd_sc_hd__inv_2 _214_ (.A(\mem_left_ipin_2.DFFR_0_.Q ),
    .Y(_201_));
 sky130_fd_sc_hd__inv_2 _215_ (.A(\mem_left_ipin_2.DFFR_2_.Q ),
    .Y(_198_));
 sky130_fd_sc_hd__inv_2 _216_ (.A(\mem_left_ipin_2.DFFR_1_.Q ),
    .Y(_197_));
 sky130_fd_sc_hd__inv_2 _217_ (.A(\mem_left_ipin_2.DFFR_5_.Q ),
    .Y(_194_));
 sky130_fd_sc_hd__inv_2 _218_ (.A(\mem_left_ipin_2.DFFR_4_.Q ),
    .Y(_193_));
 sky130_fd_sc_hd__inv_2 _219_ (.A(\mem_left_ipin_2.DFFR_0_.Q ),
    .Y(_200_));
 sky130_fd_sc_hd__inv_2 _220_ (.A(\mem_left_ipin_2.DFFR_2_.Q ),
    .Y(_196_));
 sky130_fd_sc_hd__inv_2 _221_ (.A(\mem_left_ipin_2.DFFR_1_.Q ),
    .Y(_195_));
 sky130_fd_sc_hd__inv_2 _222_ (.A(\mem_right_ipin_7.DFFR_3_.Q ),
    .Y(_189_));
 sky130_fd_sc_hd__inv_2 _223_ (.A(\mem_right_ipin_7.DFFR_0_.Q ),
    .Y(_192_));
 sky130_fd_sc_hd__inv_2 _224_ (.A(\mem_right_ipin_7.DFFR_2_.Q ),
    .Y(_188_));
 sky130_fd_sc_hd__inv_2 _225_ (.A(\mem_right_ipin_7.DFFR_1_.Q ),
    .Y(_187_));
 sky130_fd_sc_hd__inv_2 _226_ (.A(net41),
    .Y(_182_));
 sky130_fd_sc_hd__inv_2 _227_ (.A(\mem_right_ipin_7.DFFR_0_.Q ),
    .Y(_190_));
 sky130_fd_sc_hd__inv_2 _228_ (.A(\mem_right_ipin_7.DFFR_2_.Q ),
    .Y(_184_));
 sky130_fd_sc_hd__inv_2 _229_ (.A(\mem_right_ipin_7.DFFR_1_.Q ),
    .Y(_183_));
 sky130_fd_sc_hd__inv_2 _230_ (.A(\mem_right_ipin_7.DFFR_4_.Q ),
    .Y(_181_));
 sky130_fd_sc_hd__inv_2 _231_ (.A(\mem_right_ipin_7.DFFR_0_.Q ),
    .Y(_191_));
 sky130_fd_sc_hd__inv_2 _232_ (.A(\mem_right_ipin_7.DFFR_2_.Q ),
    .Y(_186_));
 sky130_fd_sc_hd__inv_2 _233_ (.A(\mem_right_ipin_7.DFFR_1_.Q ),
    .Y(_185_));
 sky130_fd_sc_hd__inv_2 _234_ (.A(\mem_right_ipin_6.DFFR_3_.Q ),
    .Y(_177_));
 sky130_fd_sc_hd__inv_2 _235_ (.A(\mem_right_ipin_6.DFFR_0_.Q ),
    .Y(_180_));
 sky130_fd_sc_hd__inv_2 _236_ (.A(\mem_right_ipin_6.DFFR_2_.Q ),
    .Y(_176_));
 sky130_fd_sc_hd__inv_2 _237_ (.A(\mem_right_ipin_6.DFFR_1_.Q ),
    .Y(_175_));
 sky130_fd_sc_hd__inv_2 _238_ (.A(\mem_right_ipin_6.DFFR_5_.Q ),
    .Y(_170_));
 sky130_fd_sc_hd__inv_2 _239_ (.A(\mem_right_ipin_6.DFFR_0_.Q ),
    .Y(_178_));
 sky130_fd_sc_hd__inv_2 _240_ (.A(\mem_right_ipin_6.DFFR_2_.Q ),
    .Y(_172_));
 sky130_fd_sc_hd__inv_2 _241_ (.A(\mem_right_ipin_6.DFFR_1_.Q ),
    .Y(_171_));
 sky130_fd_sc_hd__inv_2 _242_ (.A(\mem_right_ipin_6.DFFR_4_.Q ),
    .Y(_169_));
 sky130_fd_sc_hd__inv_2 _243_ (.A(\mem_right_ipin_6.DFFR_0_.Q ),
    .Y(_179_));
 sky130_fd_sc_hd__inv_2 _244_ (.A(\mem_right_ipin_6.DFFR_2_.Q ),
    .Y(_174_));
 sky130_fd_sc_hd__inv_2 _245_ (.A(\mem_right_ipin_6.DFFR_1_.Q ),
    .Y(_173_));
 sky130_fd_sc_hd__inv_2 _246_ (.A(\mem_right_ipin_5.DFFR_3_.Q ),
    .Y(_165_));
 sky130_fd_sc_hd__inv_2 _247_ (.A(\mem_right_ipin_5.DFFR_0_.Q ),
    .Y(_168_));
 sky130_fd_sc_hd__inv_2 _248_ (.A(\mem_right_ipin_5.DFFR_2_.Q ),
    .Y(_164_));
 sky130_fd_sc_hd__inv_2 _249_ (.A(\mem_right_ipin_5.DFFR_1_.Q ),
    .Y(_163_));
 sky130_fd_sc_hd__inv_2 _250_ (.A(\mem_right_ipin_5.DFFR_5_.Q ),
    .Y(_158_));
 sky130_fd_sc_hd__inv_2 _251_ (.A(\mem_right_ipin_5.DFFR_0_.Q ),
    .Y(_166_));
 sky130_fd_sc_hd__inv_2 _252_ (.A(\mem_right_ipin_5.DFFR_2_.Q ),
    .Y(_160_));
 sky130_fd_sc_hd__inv_2 _253_ (.A(\mem_right_ipin_5.DFFR_1_.Q ),
    .Y(_159_));
 sky130_fd_sc_hd__inv_2 _254_ (.A(\mem_right_ipin_5.DFFR_4_.Q ),
    .Y(_157_));
 sky130_fd_sc_hd__inv_2 _255_ (.A(\mem_right_ipin_5.DFFR_0_.Q ),
    .Y(_167_));
 sky130_fd_sc_hd__inv_2 _256_ (.A(\mem_right_ipin_5.DFFR_2_.Q ),
    .Y(_162_));
 sky130_fd_sc_hd__inv_2 _257_ (.A(\mem_right_ipin_5.DFFR_1_.Q ),
    .Y(_161_));
 sky130_fd_sc_hd__inv_2 _258_ (.A(\mem_right_ipin_4.DFFR_3_.Q ),
    .Y(_153_));
 sky130_fd_sc_hd__inv_2 _259_ (.A(\mem_right_ipin_4.DFFR_0_.Q ),
    .Y(_156_));
 sky130_fd_sc_hd__inv_2 _260_ (.A(\mem_right_ipin_4.DFFR_2_.Q ),
    .Y(_152_));
 sky130_fd_sc_hd__inv_2 _261_ (.A(\mem_right_ipin_4.DFFR_1_.Q ),
    .Y(_151_));
 sky130_fd_sc_hd__inv_2 _262_ (.A(\mem_right_ipin_4.DFFR_5_.Q ),
    .Y(_146_));
 sky130_fd_sc_hd__inv_2 _263_ (.A(\mem_right_ipin_4.DFFR_0_.Q ),
    .Y(_154_));
 sky130_fd_sc_hd__inv_2 _264_ (.A(\mem_right_ipin_4.DFFR_2_.Q ),
    .Y(_148_));
 sky130_fd_sc_hd__inv_2 _265_ (.A(\mem_right_ipin_4.DFFR_1_.Q ),
    .Y(_147_));
 sky130_fd_sc_hd__inv_2 _266_ (.A(\mem_right_ipin_4.DFFR_4_.Q ),
    .Y(_145_));
 sky130_fd_sc_hd__inv_2 _267_ (.A(\mem_right_ipin_4.DFFR_0_.Q ),
    .Y(_155_));
 sky130_fd_sc_hd__inv_2 _268_ (.A(\mem_right_ipin_4.DFFR_2_.Q ),
    .Y(_150_));
 sky130_fd_sc_hd__inv_2 _269_ (.A(\mem_right_ipin_4.DFFR_1_.Q ),
    .Y(_149_));
 sky130_fd_sc_hd__inv_2 _270_ (.A(\mem_right_ipin_3.DFFR_3_.Q ),
    .Y(_141_));
 sky130_fd_sc_hd__inv_2 _271_ (.A(\mem_right_ipin_3.DFFR_0_.Q ),
    .Y(_144_));
 sky130_fd_sc_hd__inv_2 _272_ (.A(\mem_right_ipin_3.DFFR_2_.Q ),
    .Y(_140_));
 sky130_fd_sc_hd__inv_2 _273_ (.A(\mem_right_ipin_3.DFFR_1_.Q ),
    .Y(_139_));
 sky130_fd_sc_hd__inv_2 _274_ (.A(\mem_right_ipin_3.DFFR_5_.Q ),
    .Y(_134_));
 sky130_fd_sc_hd__inv_2 _275_ (.A(\mem_right_ipin_3.DFFR_0_.Q ),
    .Y(_142_));
 sky130_fd_sc_hd__inv_2 _276_ (.A(\mem_right_ipin_3.DFFR_2_.Q ),
    .Y(_136_));
 sky130_fd_sc_hd__inv_2 _277_ (.A(\mem_right_ipin_3.DFFR_1_.Q ),
    .Y(_135_));
 sky130_fd_sc_hd__inv_2 _278_ (.A(\mem_right_ipin_3.DFFR_4_.Q ),
    .Y(_133_));
 sky130_fd_sc_hd__inv_2 _279_ (.A(\mem_right_ipin_3.DFFR_0_.Q ),
    .Y(_143_));
 sky130_fd_sc_hd__inv_2 _280_ (.A(\mem_right_ipin_3.DFFR_2_.Q ),
    .Y(_138_));
 sky130_fd_sc_hd__inv_2 _281_ (.A(\mem_right_ipin_3.DFFR_1_.Q ),
    .Y(_137_));
 sky130_fd_sc_hd__inv_2 _282_ (.A(\mem_right_ipin_2.DFFR_3_.Q ),
    .Y(_129_));
 sky130_fd_sc_hd__inv_2 _283_ (.A(\mem_right_ipin_2.DFFR_0_.Q ),
    .Y(_132_));
 sky130_fd_sc_hd__inv_2 _284_ (.A(\mem_right_ipin_2.DFFR_2_.Q ),
    .Y(_128_));
 sky130_fd_sc_hd__inv_2 _285_ (.A(\mem_right_ipin_2.DFFR_1_.Q ),
    .Y(_127_));
 sky130_fd_sc_hd__inv_2 _286_ (.A(\mem_right_ipin_2.DFFR_5_.Q ),
    .Y(_122_));
 sky130_fd_sc_hd__inv_2 _287_ (.A(\mem_right_ipin_2.DFFR_0_.Q ),
    .Y(_130_));
 sky130_fd_sc_hd__inv_2 _288_ (.A(\mem_right_ipin_2.DFFR_2_.Q ),
    .Y(_124_));
 sky130_fd_sc_hd__inv_2 _289_ (.A(\mem_right_ipin_2.DFFR_1_.Q ),
    .Y(_123_));
 sky130_fd_sc_hd__inv_2 _290_ (.A(\mem_right_ipin_2.DFFR_4_.Q ),
    .Y(_121_));
 sky130_fd_sc_hd__inv_2 _291_ (.A(\mem_right_ipin_2.DFFR_0_.Q ),
    .Y(_131_));
 sky130_fd_sc_hd__inv_2 _292_ (.A(\mem_right_ipin_2.DFFR_2_.Q ),
    .Y(_126_));
 sky130_fd_sc_hd__inv_2 _293_ (.A(\mem_right_ipin_2.DFFR_1_.Q ),
    .Y(_125_));
 sky130_fd_sc_hd__inv_2 _294_ (.A(\mem_right_ipin_1.DFFR_3_.Q ),
    .Y(_117_));
 sky130_fd_sc_hd__inv_2 _295_ (.A(\mem_right_ipin_1.DFFR_0_.Q ),
    .Y(_120_));
 sky130_fd_sc_hd__inv_2 _296_ (.A(\mem_right_ipin_1.DFFR_2_.Q ),
    .Y(_116_));
 sky130_fd_sc_hd__inv_2 _297_ (.A(\mem_right_ipin_1.DFFR_1_.Q ),
    .Y(_115_));
 sky130_fd_sc_hd__inv_2 _298_ (.A(\mem_right_ipin_1.DFFR_5_.Q ),
    .Y(_110_));
 sky130_fd_sc_hd__inv_2 _299_ (.A(\mem_right_ipin_1.DFFR_0_.Q ),
    .Y(_118_));
 sky130_fd_sc_hd__inv_2 _300_ (.A(\mem_right_ipin_1.DFFR_2_.Q ),
    .Y(_112_));
 sky130_fd_sc_hd__inv_2 _301_ (.A(\mem_right_ipin_1.DFFR_1_.Q ),
    .Y(_111_));
 sky130_fd_sc_hd__inv_2 _302_ (.A(\mem_right_ipin_1.DFFR_4_.Q ),
    .Y(_109_));
 sky130_fd_sc_hd__inv_2 _303_ (.A(\mem_right_ipin_1.DFFR_0_.Q ),
    .Y(_119_));
 sky130_fd_sc_hd__inv_2 _304_ (.A(\mem_right_ipin_1.DFFR_2_.Q ),
    .Y(_114_));
 sky130_fd_sc_hd__inv_2 _305_ (.A(\mem_right_ipin_1.DFFR_1_.Q ),
    .Y(_113_));
 sky130_fd_sc_hd__inv_2 _306_ (.A(\mem_right_ipin_0.DFFR_3_.Q ),
    .Y(_105_));
 sky130_fd_sc_hd__inv_2 _307_ (.A(\mem_right_ipin_0.DFFR_0_.Q ),
    .Y(_108_));
 sky130_fd_sc_hd__inv_2 _308_ (.A(\mem_right_ipin_0.DFFR_2_.Q ),
    .Y(_104_));
 sky130_fd_sc_hd__inv_2 _309_ (.A(\mem_right_ipin_0.DFFR_1_.Q ),
    .Y(_103_));
 sky130_fd_sc_hd__inv_2 _310_ (.A(\mem_right_ipin_0.DFFR_5_.Q ),
    .Y(_098_));
 sky130_fd_sc_hd__inv_2 _311_ (.A(\mem_right_ipin_0.DFFR_0_.Q ),
    .Y(_106_));
 sky130_fd_sc_hd__inv_2 _312_ (.A(\mem_right_ipin_0.DFFR_2_.Q ),
    .Y(_100_));
 sky130_fd_sc_hd__inv_2 _313_ (.A(\mem_right_ipin_0.DFFR_1_.Q ),
    .Y(_099_));
 sky130_fd_sc_hd__inv_2 _314_ (.A(\mem_right_ipin_0.DFFR_4_.Q ),
    .Y(_097_));
 sky130_fd_sc_hd__inv_2 _315_ (.A(\mem_right_ipin_0.DFFR_0_.Q ),
    .Y(_107_));
 sky130_fd_sc_hd__inv_2 _316_ (.A(\mem_right_ipin_0.DFFR_2_.Q ),
    .Y(_102_));
 sky130_fd_sc_hd__inv_2 _317_ (.A(\mem_right_ipin_0.DFFR_1_.Q ),
    .Y(_101_));
 sky130_fd_sc_hd__inv_2 _318_ (.A(\mem_left_ipin_1.DFFR_3_.Q ),
    .Y(_093_));
 sky130_fd_sc_hd__inv_2 _319_ (.A(\mem_left_ipin_1.DFFR_0_.Q ),
    .Y(_096_));
 sky130_fd_sc_hd__inv_2 _320_ (.A(\mem_left_ipin_1.DFFR_1_.Q ),
    .Y(_090_));
 sky130_fd_sc_hd__inv_2 _321_ (.A(\mem_left_ipin_1.DFFR_2_.Q ),
    .Y(_089_));
 sky130_fd_sc_hd__inv_2 _322_ (.A(\mem_left_ipin_1.DFFR_5_.Q ),
    .Y(_088_));
 sky130_fd_sc_hd__inv_2 _323_ (.A(\mem_left_ipin_1.DFFR_0_.Q ),
    .Y(_094_));
 sky130_fd_sc_hd__inv_2 _324_ (.A(\mem_left_ipin_1.DFFR_1_.Q ),
    .Y(_087_));
 sky130_fd_sc_hd__inv_2 _325_ (.A(\mem_left_ipin_1.DFFR_2_.Q ),
    .Y(_086_));
 sky130_fd_sc_hd__inv_2 _326_ (.A(\mem_left_ipin_1.DFFR_4_.Q ),
    .Y(_085_));
 sky130_fd_sc_hd__inv_2 _327_ (.A(\mem_left_ipin_1.DFFR_0_.Q ),
    .Y(_095_));
 sky130_fd_sc_hd__inv_2 _328_ (.A(\mem_left_ipin_1.DFFR_1_.Q ),
    .Y(_092_));
 sky130_fd_sc_hd__inv_2 _329_ (.A(\mem_left_ipin_1.DFFR_2_.Q ),
    .Y(_091_));
 sky130_fd_sc_hd__inv_2 _330_ (.A(\mem_left_ipin_0.DFFR_3_.Q ),
    .Y(_084_));
 sky130_fd_sc_hd__inv_2 _331_ (.A(\mem_left_ipin_0.DFFR_0_.Q ),
    .Y(_081_));
 sky130_fd_sc_hd__inv_2 _332_ (.A(\mem_left_ipin_0.DFFR_4_.Q ),
    .Y(_080_));
 sky130_fd_sc_hd__inv_2 _333_ (.A(\mem_left_ipin_0.DFFR_0_.Q ),
    .Y(_082_));
 sky130_fd_sc_hd__inv_2 _334_ (.A(\mem_left_ipin_0.DFFR_5_.Q ),
    .Y(_079_));
 sky130_fd_sc_hd__inv_2 _335_ (.A(\mem_left_ipin_0.DFFR_0_.Q ),
    .Y(_083_));
 sky130_fd_sc_hd__inv_2 _336_ (.A(\mem_left_ipin_0.DFFR_1_.Q ),
    .Y(_078_));
 sky130_fd_sc_hd__inv_2 _337_ (.A(\mem_left_ipin_0.DFFR_2_.Q ),
    .Y(_077_));
 sky130_fd_sc_hd__inv_2 _338_ (.A(\mem_left_ipin_0.DFFR_1_.Q ),
    .Y(_076_));
 sky130_fd_sc_hd__inv_2 _339_ (.A(\mem_left_ipin_0.DFFR_2_.Q ),
    .Y(_075_));
 sky130_fd_sc_hd__inv_2 _340_ (.A(\mem_left_ipin_0.DFFR_1_.Q ),
    .Y(_074_));
 sky130_fd_sc_hd__inv_2 _341_ (.A(\mem_left_ipin_0.DFFR_2_.Q ),
    .Y(_073_));
 sky130_fd_sc_hd__inv_2 _342_ (.A(net24),
    .Y(\mux_left_ipin_0.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _343_ (.A(net11),
    .Y(\mux_left_ipin_0.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _344_ (.A(\mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net89));
 sky130_fd_sc_hd__inv_2 _345_ (.A(net30),
    .Y(\mux_left_ipin_0.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _346_ (.A(net2),
    .Y(\mux_left_ipin_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _347_ (.A(net21),
    .Y(\mux_left_ipin_0.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _348_ (.A(net17),
    .Y(\mux_left_ipin_0.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _349_ (.A(net36),
    .Y(\mux_left_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _350_ (.A(net5),
    .Y(\mux_left_ipin_0.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _351_ (.A(\mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net90));
 sky130_fd_sc_hd__inv_2 _352_ (.A(net6),
    .Y(\mux_left_ipin_1.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _353_ (.A(net37),
    .Y(\mux_left_ipin_1.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _354_ (.A(net18),
    .Y(\mux_left_ipin_1.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _355_ (.A(net31),
    .Y(\mux_left_ipin_1.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _356_ (.A(net12),
    .Y(\mux_left_ipin_1.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _357_ (.A(net25),
    .Y(\mux_left_ipin_1.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _358_ (.A(\mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net80));
 sky130_fd_sc_hd__inv_2 _359_ (.A(net8),
    .Y(\mux_right_ipin_0.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _360_ (.A(net39),
    .Y(\mux_right_ipin_0.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _361_ (.A(net20),
    .Y(\mux_right_ipin_0.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _362_ (.A(net33),
    .Y(\mux_right_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _363_ (.A(net14),
    .Y(\mux_right_ipin_0.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _364_ (.A(net27),
    .Y(\mux_right_ipin_0.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _365_ (.A(\mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net81));
 sky130_fd_sc_hd__inv_2 _366_ (.A(net9),
    .Y(\mux_right_ipin_1.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _367_ (.A(net22),
    .Y(\mux_right_ipin_1.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _368_ (.A(net3),
    .Y(\mux_right_ipin_1.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _369_ (.A(net34),
    .Y(\mux_right_ipin_1.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _370_ (.A(net15),
    .Y(\mux_right_ipin_1.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _371_ (.A(net28),
    .Y(\mux_right_ipin_1.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _372_ (.A(\mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net82));
 sky130_fd_sc_hd__inv_2 _373_ (.A(net10),
    .Y(\mux_right_ipin_2.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _374_ (.A(net35),
    .Y(\mux_right_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _375_ (.A(net16),
    .Y(\mux_right_ipin_2.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _376_ (.A(net29),
    .Y(\mux_right_ipin_2.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _377_ (.A(\mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net83));
 sky130_fd_sc_hd__inv_2 _378_ (.A(\mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net84));
 sky130_fd_sc_hd__inv_2 _379_ (.A(\mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net85));
 sky130_fd_sc_hd__clkinv_2 _380_ (.A(net7),
    .Y(\mux_right_ipin_5.INVTX1_6_.out ));
 sky130_fd_sc_hd__inv_2 _381_ (.A(net38),
    .Y(\mux_right_ipin_5.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_2 _382_ (.A(net19),
    .Y(\mux_right_ipin_5.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _383_ (.A(net26),
    .Y(\mux_right_ipin_5.INVTX1_7_.out ));
 sky130_fd_sc_hd__inv_2 _384_ (.A(\mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net86));
 sky130_fd_sc_hd__inv_2 _385_ (.A(\mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out ),
    .Y(net87));
 sky130_fd_sc_hd__inv_2 _386_ (.A(\mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .Y(net88));
 sky130_fd_sc_hd__inv_2 _387_ (.A(net4),
    .Y(\mux_left_ipin_2.INVTX1_4_.out ));
 sky130_fd_sc_hd__inv_2 _388_ (.A(net32),
    .Y(\mux_left_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__inv_2 _389_ (.A(net13),
    .Y(\mux_left_ipin_2.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _390_ (.A(net23),
    .Y(\mux_left_ipin_2.INVTX1_5_.out ));
 sky130_fd_sc_hd__clkbuf_4 _391_ (.A(net40),
    .X(_066_));
 sky130_fd_sc_hd__buf_4 _392_ (.A(_066_),
    .X(_067_));
 sky130_fd_sc_hd__inv_2 _393_ (.A(_067_),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _394_ (.A(_067_),
    .Y(_001_));
 sky130_fd_sc_hd__inv_2 _395_ (.A(_067_),
    .Y(_002_));
 sky130_fd_sc_hd__inv_2 _396_ (.A(_067_),
    .Y(_003_));
 sky130_fd_sc_hd__inv_2 _397_ (.A(_067_),
    .Y(_004_));
 sky130_fd_sc_hd__inv_2 _398_ (.A(_067_),
    .Y(_005_));
 sky130_fd_sc_hd__inv_2 _399_ (.A(_067_),
    .Y(_006_));
 sky130_fd_sc_hd__inv_2 _400_ (.A(_067_),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _401_ (.A(_067_),
    .Y(_008_));
 sky130_fd_sc_hd__inv_2 _402_ (.A(_067_),
    .Y(_009_));
 sky130_fd_sc_hd__buf_4 _403_ (.A(_066_),
    .X(_068_));
 sky130_fd_sc_hd__inv_2 _404_ (.A(_068_),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _405_ (.A(_068_),
    .Y(_011_));
 sky130_fd_sc_hd__inv_2 _406_ (.A(_068_),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _407_ (.A(_068_),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _408_ (.A(_068_),
    .Y(_014_));
 sky130_fd_sc_hd__inv_2 _409_ (.A(_068_),
    .Y(_015_));
 sky130_fd_sc_hd__inv_2 _410_ (.A(_068_),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _411_ (.A(_068_),
    .Y(_017_));
 sky130_fd_sc_hd__inv_2 _412_ (.A(_068_),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _413_ (.A(_068_),
    .Y(_019_));
 sky130_fd_sc_hd__buf_4 _414_ (.A(_066_),
    .X(_069_));
 sky130_fd_sc_hd__inv_2 _415_ (.A(_069_),
    .Y(_020_));
 sky130_fd_sc_hd__inv_2 _416_ (.A(_069_),
    .Y(_021_));
 sky130_fd_sc_hd__inv_2 _417_ (.A(_069_),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _418_ (.A(_069_),
    .Y(_023_));
 sky130_fd_sc_hd__inv_2 _419_ (.A(_069_),
    .Y(_024_));
 sky130_fd_sc_hd__inv_2 _420_ (.A(_069_),
    .Y(_025_));
 sky130_fd_sc_hd__inv_2 _421_ (.A(_069_),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _422_ (.A(_069_),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _423_ (.A(_069_),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _424_ (.A(_069_),
    .Y(_029_));
 sky130_fd_sc_hd__clkbuf_8 _425_ (.A(_066_),
    .X(_070_));
 sky130_fd_sc_hd__inv_2 _426_ (.A(_070_),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _427_ (.A(_070_),
    .Y(_031_));
 sky130_fd_sc_hd__inv_2 _428_ (.A(_070_),
    .Y(_032_));
 sky130_fd_sc_hd__inv_2 _429_ (.A(_070_),
    .Y(_033_));
 sky130_fd_sc_hd__inv_2 _430_ (.A(_070_),
    .Y(_034_));
 sky130_fd_sc_hd__inv_2 _431_ (.A(_070_),
    .Y(_035_));
 sky130_fd_sc_hd__inv_2 _432_ (.A(_070_),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _433_ (.A(_070_),
    .Y(_037_));
 sky130_fd_sc_hd__inv_2 _434_ (.A(_070_),
    .Y(_038_));
 sky130_fd_sc_hd__inv_2 _435_ (.A(_070_),
    .Y(_039_));
 sky130_fd_sc_hd__buf_4 _436_ (.A(net40),
    .X(_071_));
 sky130_fd_sc_hd__inv_2 _437_ (.A(_071_),
    .Y(_040_));
 sky130_fd_sc_hd__inv_2 _438_ (.A(_071_),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _439_ (.A(_071_),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _440_ (.A(_071_),
    .Y(_043_));
 sky130_fd_sc_hd__inv_2 _441_ (.A(_071_),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _442_ (.A(_071_),
    .Y(_045_));
 sky130_fd_sc_hd__inv_2 _443_ (.A(_071_),
    .Y(_046_));
 sky130_fd_sc_hd__inv_2 _444_ (.A(_071_),
    .Y(_047_));
 sky130_fd_sc_hd__inv_2 _445_ (.A(_071_),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _446_ (.A(_071_),
    .Y(_049_));
 sky130_fd_sc_hd__buf_4 _447_ (.A(net40),
    .X(_072_));
 sky130_fd_sc_hd__inv_2 _448_ (.A(_072_),
    .Y(_050_));
 sky130_fd_sc_hd__inv_2 _449_ (.A(_072_),
    .Y(_051_));
 sky130_fd_sc_hd__inv_2 _450_ (.A(_072_),
    .Y(_052_));
 sky130_fd_sc_hd__inv_2 _451_ (.A(_072_),
    .Y(_053_));
 sky130_fd_sc_hd__inv_2 _452_ (.A(_072_),
    .Y(_054_));
 sky130_fd_sc_hd__inv_2 _453_ (.A(_072_),
    .Y(_055_));
 sky130_fd_sc_hd__inv_2 _454_ (.A(_072_),
    .Y(_056_));
 sky130_fd_sc_hd__inv_2 _455_ (.A(_072_),
    .Y(_057_));
 sky130_fd_sc_hd__inv_2 _456_ (.A(_072_),
    .Y(_058_));
 sky130_fd_sc_hd__inv_2 _457_ (.A(_072_),
    .Y(_059_));
 sky130_fd_sc_hd__inv_2 _458_ (.A(_066_),
    .Y(_060_));
 sky130_fd_sc_hd__inv_2 _459_ (.A(_066_),
    .Y(_061_));
 sky130_fd_sc_hd__inv_2 _460_ (.A(_066_),
    .Y(_062_));
 sky130_fd_sc_hd__inv_2 _461_ (.A(_066_),
    .Y(_063_));
 sky130_fd_sc_hd__inv_2 _462_ (.A(_066_),
    .Y(_064_));
 sky130_fd_sc_hd__inv_2 _463_ (.A(_066_),
    .Y(_065_));
 sky130_fd_sc_hd__dfrtp_1 _464_ (.CLK(prog_clk),
    .D(\mem_left_ipin_0.DFFR_4_.Q ),
    .RESET_B(_000_),
    .Q(\mem_left_ipin_0.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _465_ (.CLK(prog_clk),
    .D(\mem_left_ipin_0.DFFR_3_.Q ),
    .RESET_B(_001_),
    .Q(\mem_left_ipin_0.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _466_ (.CLK(prog_clk),
    .D(\mem_left_ipin_0.DFFR_2_.Q ),
    .RESET_B(_002_),
    .Q(\mem_left_ipin_0.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _467_ (.CLK(prog_clk),
    .D(\mem_left_ipin_0.DFFR_1_.Q ),
    .RESET_B(_003_),
    .Q(\mem_left_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _468_ (.CLK(prog_clk),
    .D(\mem_left_ipin_0.DFFR_0_.Q ),
    .RESET_B(_004_),
    .Q(\mem_left_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _469_ (.CLK(prog_clk),
    .D(net1),
    .RESET_B(_005_),
    .Q(\mem_left_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _470_ (.CLK(prog_clk),
    .D(\mem_left_ipin_1.DFFR_4_.Q ),
    .RESET_B(_006_),
    .Q(\mem_left_ipin_1.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _471_ (.CLK(prog_clk),
    .D(\mem_left_ipin_1.DFFR_3_.Q ),
    .RESET_B(_007_),
    .Q(\mem_left_ipin_1.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _472_ (.CLK(prog_clk),
    .D(\mem_left_ipin_1.DFFR_2_.Q ),
    .RESET_B(_008_),
    .Q(\mem_left_ipin_1.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _473_ (.CLK(prog_clk),
    .D(\mem_left_ipin_1.DFFR_1_.Q ),
    .RESET_B(_009_),
    .Q(\mem_left_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _474_ (.CLK(prog_clk),
    .D(\mem_left_ipin_1.DFFR_0_.Q ),
    .RESET_B(_010_),
    .Q(\mem_left_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _475_ (.CLK(prog_clk),
    .D(\mem_left_ipin_0.DFFR_5_.Q ),
    .RESET_B(_011_),
    .Q(\mem_left_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _476_ (.CLK(prog_clk),
    .D(\mem_right_ipin_0.DFFR_4_.Q ),
    .RESET_B(_012_),
    .Q(\mem_right_ipin_0.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _477_ (.CLK(prog_clk),
    .D(\mem_right_ipin_0.DFFR_3_.Q ),
    .RESET_B(_013_),
    .Q(\mem_right_ipin_0.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _478_ (.CLK(prog_clk),
    .D(\mem_right_ipin_0.DFFR_2_.Q ),
    .RESET_B(_014_),
    .Q(\mem_right_ipin_0.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _479_ (.CLK(prog_clk),
    .D(\mem_right_ipin_0.DFFR_1_.Q ),
    .RESET_B(_015_),
    .Q(\mem_right_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _480_ (.CLK(prog_clk),
    .D(\mem_right_ipin_0.DFFR_0_.Q ),
    .RESET_B(_016_),
    .Q(\mem_right_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _481_ (.CLK(prog_clk),
    .D(\mem_left_ipin_2.DFFR_5_.Q ),
    .RESET_B(_017_),
    .Q(\mem_right_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _482_ (.CLK(prog_clk),
    .D(\mem_right_ipin_1.DFFR_4_.Q ),
    .RESET_B(_018_),
    .Q(\mem_right_ipin_1.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _483_ (.CLK(prog_clk),
    .D(\mem_right_ipin_1.DFFR_3_.Q ),
    .RESET_B(_019_),
    .Q(\mem_right_ipin_1.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _484_ (.CLK(prog_clk),
    .D(\mem_right_ipin_1.DFFR_2_.Q ),
    .RESET_B(_020_),
    .Q(\mem_right_ipin_1.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _485_ (.CLK(prog_clk),
    .D(\mem_right_ipin_1.DFFR_1_.Q ),
    .RESET_B(_021_),
    .Q(\mem_right_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _486_ (.CLK(prog_clk),
    .D(\mem_right_ipin_1.DFFR_0_.Q ),
    .RESET_B(_022_),
    .Q(\mem_right_ipin_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _487_ (.CLK(prog_clk),
    .D(\mem_right_ipin_0.DFFR_5_.Q ),
    .RESET_B(_023_),
    .Q(\mem_right_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _488_ (.CLK(prog_clk),
    .D(\mem_right_ipin_2.DFFR_4_.Q ),
    .RESET_B(_024_),
    .Q(\mem_right_ipin_2.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _489_ (.CLK(prog_clk),
    .D(\mem_right_ipin_2.DFFR_3_.Q ),
    .RESET_B(_025_),
    .Q(\mem_right_ipin_2.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _490_ (.CLK(prog_clk),
    .D(\mem_right_ipin_2.DFFR_2_.Q ),
    .RESET_B(_026_),
    .Q(\mem_right_ipin_2.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _491_ (.CLK(prog_clk),
    .D(\mem_right_ipin_2.DFFR_1_.Q ),
    .RESET_B(_027_),
    .Q(\mem_right_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _492_ (.CLK(prog_clk),
    .D(\mem_right_ipin_2.DFFR_0_.Q ),
    .RESET_B(_028_),
    .Q(\mem_right_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _493_ (.CLK(prog_clk),
    .D(\mem_right_ipin_1.DFFR_5_.Q ),
    .RESET_B(_029_),
    .Q(\mem_right_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _494_ (.CLK(prog_clk),
    .D(\mem_right_ipin_3.DFFR_4_.Q ),
    .RESET_B(_030_),
    .Q(\mem_right_ipin_3.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _495_ (.CLK(prog_clk),
    .D(\mem_right_ipin_3.DFFR_3_.Q ),
    .RESET_B(_031_),
    .Q(\mem_right_ipin_3.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _496_ (.CLK(prog_clk),
    .D(\mem_right_ipin_3.DFFR_2_.Q ),
    .RESET_B(_032_),
    .Q(\mem_right_ipin_3.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _497_ (.CLK(prog_clk),
    .D(\mem_right_ipin_3.DFFR_1_.Q ),
    .RESET_B(_033_),
    .Q(\mem_right_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _498_ (.CLK(prog_clk),
    .D(\mem_right_ipin_3.DFFR_0_.Q ),
    .RESET_B(_034_),
    .Q(\mem_right_ipin_3.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _499_ (.CLK(prog_clk),
    .D(\mem_right_ipin_2.DFFR_5_.Q ),
    .RESET_B(_035_),
    .Q(\mem_right_ipin_3.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _500_ (.CLK(prog_clk),
    .D(\mem_right_ipin_4.DFFR_4_.Q ),
    .RESET_B(_036_),
    .Q(\mem_right_ipin_4.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _501_ (.CLK(prog_clk),
    .D(\mem_right_ipin_4.DFFR_3_.Q ),
    .RESET_B(_037_),
    .Q(\mem_right_ipin_4.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _502_ (.CLK(prog_clk),
    .D(\mem_right_ipin_4.DFFR_2_.Q ),
    .RESET_B(_038_),
    .Q(\mem_right_ipin_4.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _503_ (.CLK(prog_clk),
    .D(\mem_right_ipin_4.DFFR_1_.Q ),
    .RESET_B(_039_),
    .Q(\mem_right_ipin_4.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _504_ (.CLK(prog_clk),
    .D(\mem_right_ipin_4.DFFR_0_.Q ),
    .RESET_B(_040_),
    .Q(\mem_right_ipin_4.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _505_ (.CLK(prog_clk),
    .D(\mem_right_ipin_3.DFFR_5_.Q ),
    .RESET_B(_041_),
    .Q(\mem_right_ipin_4.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _506_ (.CLK(prog_clk),
    .D(\mem_right_ipin_5.DFFR_4_.Q ),
    .RESET_B(_042_),
    .Q(\mem_right_ipin_5.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _507_ (.CLK(prog_clk),
    .D(\mem_right_ipin_5.DFFR_3_.Q ),
    .RESET_B(_043_),
    .Q(\mem_right_ipin_5.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _508_ (.CLK(prog_clk),
    .D(\mem_right_ipin_5.DFFR_2_.Q ),
    .RESET_B(_044_),
    .Q(\mem_right_ipin_5.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _509_ (.CLK(prog_clk),
    .D(\mem_right_ipin_5.DFFR_1_.Q ),
    .RESET_B(_045_),
    .Q(\mem_right_ipin_5.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _510_ (.CLK(prog_clk),
    .D(\mem_right_ipin_5.DFFR_0_.Q ),
    .RESET_B(_046_),
    .Q(\mem_right_ipin_5.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _511_ (.CLK(prog_clk),
    .D(\mem_right_ipin_4.DFFR_5_.Q ),
    .RESET_B(_047_),
    .Q(\mem_right_ipin_5.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _512_ (.CLK(prog_clk),
    .D(\mem_right_ipin_6.DFFR_4_.Q ),
    .RESET_B(_048_),
    .Q(\mem_right_ipin_6.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _513_ (.CLK(prog_clk),
    .D(\mem_right_ipin_6.DFFR_3_.Q ),
    .RESET_B(_049_),
    .Q(\mem_right_ipin_6.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _514_ (.CLK(prog_clk),
    .D(\mem_right_ipin_6.DFFR_2_.Q ),
    .RESET_B(_050_),
    .Q(\mem_right_ipin_6.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _515_ (.CLK(prog_clk),
    .D(\mem_right_ipin_6.DFFR_1_.Q ),
    .RESET_B(_051_),
    .Q(\mem_right_ipin_6.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _516_ (.CLK(prog_clk),
    .D(\mem_right_ipin_6.DFFR_0_.Q ),
    .RESET_B(_052_),
    .Q(\mem_right_ipin_6.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _517_ (.CLK(prog_clk),
    .D(\mem_right_ipin_5.DFFR_5_.Q ),
    .RESET_B(_053_),
    .Q(\mem_right_ipin_6.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _518_ (.CLK(prog_clk),
    .D(\mem_right_ipin_7.DFFR_4_.Q ),
    .RESET_B(_054_),
    .Q(net41));
 sky130_fd_sc_hd__dfrtp_1 _519_ (.CLK(prog_clk),
    .D(\mem_right_ipin_7.DFFR_3_.Q ),
    .RESET_B(_055_),
    .Q(\mem_right_ipin_7.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _520_ (.CLK(prog_clk),
    .D(\mem_right_ipin_7.DFFR_2_.Q ),
    .RESET_B(_056_),
    .Q(\mem_right_ipin_7.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _521_ (.CLK(prog_clk),
    .D(\mem_right_ipin_7.DFFR_1_.Q ),
    .RESET_B(_057_),
    .Q(\mem_right_ipin_7.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _522_ (.CLK(prog_clk),
    .D(\mem_right_ipin_7.DFFR_0_.Q ),
    .RESET_B(_058_),
    .Q(\mem_right_ipin_7.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _523_ (.CLK(prog_clk),
    .D(\mem_right_ipin_6.DFFR_5_.Q ),
    .RESET_B(_059_),
    .Q(\mem_right_ipin_7.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _524_ (.CLK(prog_clk),
    .D(\mem_left_ipin_2.DFFR_4_.Q ),
    .RESET_B(_060_),
    .Q(\mem_left_ipin_2.DFFR_5_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _525_ (.CLK(prog_clk),
    .D(\mem_left_ipin_2.DFFR_3_.Q ),
    .RESET_B(_061_),
    .Q(\mem_left_ipin_2.DFFR_4_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _526_ (.CLK(prog_clk),
    .D(\mem_left_ipin_2.DFFR_2_.Q ),
    .RESET_B(_062_),
    .Q(\mem_left_ipin_2.DFFR_3_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _527_ (.CLK(prog_clk),
    .D(\mem_left_ipin_2.DFFR_1_.Q ),
    .RESET_B(_063_),
    .Q(\mem_left_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _528_ (.CLK(prog_clk),
    .D(\mem_left_ipin_2.DFFR_0_.Q ),
    .RESET_B(_064_),
    .Q(\mem_left_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _529_ (.CLK(prog_clk),
    .D(\mem_left_ipin_1.DFFR_5_.Q ),
    .RESET_B(_065_),
    .Q(\mem_left_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__conb_1 _592__92 (.HI(net92));
 sky130_fd_sc_hd__conb_1 _606__93 (.HI(net93));
 sky130_fd_sc_hd__conb_1 _618__94 (.HI(net94));
 sky130_fd_sc_hd__conb_1 _630__95 (.HI(net95));
 sky130_fd_sc_hd__conb_1 _642__96 (.HI(net96));
 sky130_fd_sc_hd__conb_1 _654__97 (.HI(net97));
 sky130_fd_sc_hd__conb_1 _666__98 (.HI(net98));
 sky130_fd_sc_hd__conb_1 _678__99 (.HI(net99));
 sky130_fd_sc_hd__conb_1 _690__100 (.HI(net100));
 sky130_fd_sc_hd__conb_1 _700__101 (.HI(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__402__A (.DIODE(_067_));
 sky130_fd_sc_hd__clkbuf_1 _541_ (.A(net4),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 _542_ (.A(net3),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 _543_ (.A(net20),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 _544_ (.A(net19),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 _545_ (.A(net18),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 _546_ (.A(net17),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _547_ (.A(net16),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _548_ (.A(net15),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 _549_ (.A(net14),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 _550_ (.A(net13),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 _551_ (.A(net12),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 _552_ (.A(net2),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 _553_ (.A(net30),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 _554_ (.A(net29),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 _555_ (.A(net28),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 _556_ (.A(net27),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 _557_ (.A(net26),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 _558_ (.A(net25),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 _559_ (.A(net24),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 _560_ (.A(net23),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 _561_ (.A(net22),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 _562_ (.A(net39),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 _563_ (.A(net38),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 _564_ (.A(net37),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 _565_ (.A(net36),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 _566_ (.A(net35),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 _567_ (.A(net34),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 _568_ (.A(net33),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 _569_ (.A(net32),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 _570_ (.A(net31),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 _571_ (.A(net21),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 _572_ (.A(net11),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 _573_ (.A(net10),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 _574_ (.A(net9),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 _575_ (.A(net8),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 _576_ (.A(net7),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 _577_ (.A(net6),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 _578_ (.A(net5),
    .X(net64));
 sky130_fd_sc_hd__ebufn_1 _579_ (.A(\mux_left_ipin_0.INVTX1_2_.out ),
    .TE_B(_073_),
    .Z(\mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_1 _580_ (.A(\mux_left_ipin_0.INVTX1_1_.out ),
    .TE_B(_074_),
    .Z(\mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_1 _581_ (.A(\mux_left_ipin_0.INVTX1_5_.out ),
    .TE_B(_075_),
    .Z(\mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_1 _582_ (.A(\mux_left_ipin_0.INVTX1_4_.out ),
    .TE_B(_076_),
    .Z(\mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _583_ (.A(net91),
    .TE_B(_077_),
    .Z(\mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _584_ (.A(\mux_left_ipin_0.INVTX1_7_.out ),
    .TE_B(_078_),
    .Z(\mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_4 _585_ (.A(\mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_079_),
    .Z(\mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_4 _586_ (.A(\mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_080_),
    .Z(\mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_1 _587_ (.A(\mux_left_ipin_0.INVTX1_0_.out ),
    .TE_B(_081_),
    .Z(\mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_1 _588_ (.A(\mux_left_ipin_0.INVTX1_3_.out ),
    .TE_B(_082_),
    .Z(\mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _589_ (.A(\mux_left_ipin_0.INVTX1_6_.out ),
    .TE_B(_083_),
    .Z(\mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_4 _590_ (.A(\mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_084_),
    .Z(\mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _591_ (.A(\mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_085_),
    .Z(\mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _592_ (.A(net92),
    .TE_B(_086_),
    .Z(\mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _593_ (.A(\mux_left_ipin_1.INVTX1_7_.out ),
    .TE_B(_087_),
    .Z(\mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _594_ (.A(\mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_088_),
    .Z(\mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _595_ (.A(\mux_left_ipin_1.INVTX1_2_.out ),
    .TE_B(_089_),
    .Z(\mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _596_ (.A(\mux_left_ipin_0.INVTX1_1_.out ),
    .TE_B(_090_),
    .Z(\mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _597_ (.A(\mux_left_ipin_1.INVTX1_5_.out ),
    .TE_B(_091_),
    .Z(\mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _598_ (.A(\mux_left_ipin_1.INVTX1_4_.out ),
    .TE_B(_092_),
    .Z(\mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _599_ (.A(\mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_093_),
    .Z(\mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _600_ (.A(\mux_left_ipin_1.INVTX1_6_.out ),
    .TE_B(_094_),
    .Z(\mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _601_ (.A(\mux_left_ipin_1.INVTX1_3_.out ),
    .TE_B(_095_),
    .Z(\mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _602_ (.A(\mux_left_ipin_0.INVTX1_0_.out ),
    .TE_B(_096_),
    .Z(\mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _603_ (.A(\mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_097_),
    .Z(\mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _604_ (.A(\mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_098_),
    .Z(\mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _605_ (.A(\mux_right_ipin_0.INVTX1_7_.out ),
    .TE_B(_099_),
    .Z(\mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _606_ (.A(net93),
    .TE_B(_100_),
    .Z(\mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _607_ (.A(\mux_right_ipin_0.INVTX1_4_.out ),
    .TE_B(_101_),
    .Z(\mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _608_ (.A(\mux_right_ipin_0.INVTX1_5_.out ),
    .TE_B(_102_),
    .Z(\mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _609_ (.A(\mux_left_ipin_2.INVTX1_3_.out ),
    .TE_B(_103_),
    .Z(\mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _610_ (.A(\mux_right_ipin_0.INVTX1_2_.out ),
    .TE_B(_104_),
    .Z(\mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _611_ (.A(\mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_105_),
    .Z(\mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _612_ (.A(\mux_right_ipin_0.INVTX1_6_.out ),
    .TE_B(_106_),
    .Z(\mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _613_ (.A(\mux_right_ipin_0.INVTX1_3_.out ),
    .TE_B(_107_),
    .Z(\mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _614_ (.A(\mux_left_ipin_2.INVTX1_2_.out ),
    .TE_B(_108_),
    .Z(\mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _615_ (.A(\mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_109_),
    .Z(\mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _616_ (.A(\mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_110_),
    .Z(\mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _617_ (.A(\mux_right_ipin_1.INVTX1_7_.out ),
    .TE_B(_111_),
    .Z(\mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _618_ (.A(net94),
    .TE_B(_112_),
    .Z(\mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _619_ (.A(\mux_right_ipin_1.INVTX1_4_.out ),
    .TE_B(_113_),
    .Z(\mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _620_ (.A(\mux_right_ipin_1.INVTX1_5_.out ),
    .TE_B(_114_),
    .Z(\mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _621_ (.A(\mux_right_ipin_0.INVTX1_3_.out ),
    .TE_B(_115_),
    .Z(\mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _622_ (.A(\mux_right_ipin_1.INVTX1_2_.out ),
    .TE_B(_116_),
    .Z(\mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _623_ (.A(\mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_117_),
    .Z(\mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _624_ (.A(\mux_right_ipin_1.INVTX1_6_.out ),
    .TE_B(_118_),
    .Z(\mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _625_ (.A(\mux_right_ipin_1.INVTX1_3_.out ),
    .TE_B(_119_),
    .Z(\mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _626_ (.A(\mux_right_ipin_0.INVTX1_2_.out ),
    .TE_B(_120_),
    .Z(\mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _627_ (.A(\mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_121_),
    .Z(\mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _628_ (.A(\mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_122_),
    .Z(\mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _629_ (.A(\mux_right_ipin_2.INVTX1_7_.out ),
    .TE_B(_123_),
    .Z(\mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _630_ (.A(net95),
    .TE_B(_124_),
    .Z(\mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _631_ (.A(\mux_left_ipin_2.INVTX1_4_.out ),
    .TE_B(_125_),
    .Z(\mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _632_ (.A(\mux_left_ipin_2.INVTX1_5_.out ),
    .TE_B(_126_),
    .Z(\mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _633_ (.A(\mux_right_ipin_1.INVTX1_3_.out ),
    .TE_B(_127_),
    .Z(\mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _634_ (.A(\mux_right_ipin_2.INVTX1_2_.out ),
    .TE_B(_128_),
    .Z(\mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _635_ (.A(\mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_129_),
    .Z(\mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _636_ (.A(\mux_right_ipin_2.INVTX1_6_.out ),
    .TE_B(_130_),
    .Z(\mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _637_ (.A(\mux_right_ipin_2.INVTX1_3_.out ),
    .TE_B(_131_),
    .Z(\mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _638_ (.A(\mux_right_ipin_1.INVTX1_2_.out ),
    .TE_B(_132_),
    .Z(\mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _639_ (.A(\mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_133_),
    .Z(\mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _640_ (.A(\mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_134_),
    .Z(\mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _641_ (.A(\mux_left_ipin_0.INVTX1_7_.out ),
    .TE_B(_135_),
    .Z(\mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _642_ (.A(net96),
    .TE_B(_136_),
    .Z(\mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _643_ (.A(\mux_left_ipin_0.INVTX1_4_.out ),
    .TE_B(_137_),
    .Z(\mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _644_ (.A(\mux_left_ipin_0.INVTX1_5_.out ),
    .TE_B(_138_),
    .Z(\mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _645_ (.A(\mux_right_ipin_2.INVTX1_3_.out ),
    .TE_B(_139_),
    .Z(\mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _646_ (.A(\mux_left_ipin_0.INVTX1_2_.out ),
    .TE_B(_140_),
    .Z(\mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _647_ (.A(\mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_141_),
    .Z(\mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _648_ (.A(\mux_left_ipin_0.INVTX1_6_.out ),
    .TE_B(_142_),
    .Z(\mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _649_ (.A(\mux_left_ipin_0.INVTX1_3_.out ),
    .TE_B(_143_),
    .Z(\mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _650_ (.A(\mux_right_ipin_2.INVTX1_2_.out ),
    .TE_B(_144_),
    .Z(\mux_right_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _651_ (.A(\mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_145_),
    .Z(\mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _652_ (.A(\mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_146_),
    .Z(\mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_1 _653_ (.A(\mux_left_ipin_1.INVTX1_7_.out ),
    .TE_B(_147_),
    .Z(\mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_1 _654_ (.A(net97),
    .TE_B(_148_),
    .Z(\mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _655_ (.A(\mux_left_ipin_1.INVTX1_4_.out ),
    .TE_B(_149_),
    .Z(\mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _656_ (.A(\mux_left_ipin_1.INVTX1_5_.out ),
    .TE_B(_150_),
    .Z(\mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _657_ (.A(\mux_left_ipin_0.INVTX1_1_.out ),
    .TE_B(_151_),
    .Z(\mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _658_ (.A(\mux_left_ipin_0.INVTX1_2_.out ),
    .TE_B(_152_),
    .Z(\mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _659_ (.A(\mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_153_),
    .Z(\mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_1 _660_ (.A(\mux_left_ipin_1.INVTX1_6_.out ),
    .TE_B(_154_),
    .Z(\mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _661_ (.A(\mux_left_ipin_0.INVTX1_3_.out ),
    .TE_B(_155_),
    .Z(\mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _662_ (.A(\mux_left_ipin_0.INVTX1_0_.out ),
    .TE_B(_156_),
    .Z(\mux_right_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _663_ (.A(\mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_157_),
    .Z(\mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _664_ (.A(\mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_158_),
    .Z(\mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _665_ (.A(\mux_right_ipin_5.INVTX1_7_.out ),
    .TE_B(_159_),
    .Z(\mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _666_ (.A(net98),
    .TE_B(_160_),
    .Z(\mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _667_ (.A(\mux_right_ipin_5.INVTX1_4_.out ),
    .TE_B(_161_),
    .Z(\mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _668_ (.A(\mux_right_ipin_5.INVTX1_5_.out ),
    .TE_B(_162_),
    .Z(\mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _669_ (.A(\mux_left_ipin_1.INVTX1_3_.out ),
    .TE_B(_163_),
    .Z(\mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _670_ (.A(\mux_left_ipin_1.INVTX1_4_.out ),
    .TE_B(_164_),
    .Z(\mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _671_ (.A(\mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_165_),
    .Z(\mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _672_ (.A(\mux_right_ipin_5.INVTX1_6_.out ),
    .TE_B(_166_),
    .Z(\mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _673_ (.A(\mux_left_ipin_1.INVTX1_5_.out ),
    .TE_B(_167_),
    .Z(\mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _674_ (.A(\mux_left_ipin_1.INVTX1_2_.out ),
    .TE_B(_168_),
    .Z(\mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _675_ (.A(\mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_169_),
    .Z(\mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_4 _676_ (.A(\mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_170_),
    .Z(\mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _677_ (.A(\mux_right_ipin_0.INVTX1_7_.out ),
    .TE_B(_171_),
    .Z(\mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _678_ (.A(net99),
    .TE_B(_172_),
    .Z(\mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _679_ (.A(\mux_right_ipin_0.INVTX1_4_.out ),
    .TE_B(_173_),
    .Z(\mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _680_ (.A(\mux_right_ipin_0.INVTX1_5_.out ),
    .TE_B(_174_),
    .Z(\mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _681_ (.A(\mux_left_ipin_2.INVTX1_3_.out ),
    .TE_B(_175_),
    .Z(\mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _682_ (.A(\mux_right_ipin_5.INVTX1_4_.out ),
    .TE_B(_176_),
    .Z(\mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _683_ (.A(\mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_177_),
    .Z(\mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _684_ (.A(\mux_right_ipin_0.INVTX1_6_.out ),
    .TE_B(_178_),
    .Z(\mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _685_ (.A(\mux_right_ipin_5.INVTX1_5_.out ),
    .TE_B(_179_),
    .Z(\mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _686_ (.A(\mux_left_ipin_2.INVTX1_2_.out ),
    .TE_B(_180_),
    .Z(\mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _687_ (.A(\mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_181_),
    .Z(\mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_4 _688_ (.A(\mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out ),
    .TE_B(_182_),
    .Z(\mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _689_ (.A(\mux_right_ipin_1.INVTX1_7_.out ),
    .TE_B(_183_),
    .Z(\mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _690_ (.A(net100),
    .TE_B(_184_),
    .Z(\mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _691_ (.A(\mux_right_ipin_1.INVTX1_4_.out ),
    .TE_B(_185_),
    .Z(\mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _692_ (.A(\mux_right_ipin_1.INVTX1_5_.out ),
    .TE_B(_186_),
    .Z(\mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _693_ (.A(\mux_right_ipin_0.INVTX1_3_.out ),
    .TE_B(_187_),
    .Z(\mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _694_ (.A(\mux_right_ipin_0.INVTX1_4_.out ),
    .TE_B(_188_),
    .Z(\mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_4 _695_ (.A(\mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_189_),
    .Z(\mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__ebufn_2 _696_ (.A(\mux_right_ipin_1.INVTX1_6_.out ),
    .TE_B(_190_),
    .Z(\mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _697_ (.A(\mux_right_ipin_0.INVTX1_5_.out ),
    .TE_B(_191_),
    .Z(\mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _698_ (.A(\mux_right_ipin_0.INVTX1_2_.out ),
    .TE_B(_192_),
    .Z(\mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _699_ (.A(\mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ),
    .TE_B(_193_),
    .Z(\mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _700_ (.A(net101),
    .TE_B(_194_),
    .Z(\mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _701_ (.A(\mux_left_ipin_2.INVTX1_4_.out ),
    .TE_B(_195_),
    .Z(\mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _702_ (.A(\mux_left_ipin_2.INVTX1_5_.out ),
    .TE_B(_196_),
    .Z(\mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _703_ (.A(\mux_left_ipin_1.INVTX1_3_.out ),
    .TE_B(_197_),
    .Z(\mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _704_ (.A(\mux_left_ipin_2.INVTX1_2_.out ),
    .TE_B(_198_),
    .Z(\mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__ebufn_2 _705_ (.A(\mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ),
    .TE_B(_199_),
    .Z(\mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__ebufn_2 _706_ (.A(\mux_left_ipin_2.INVTX1_3_.out ),
    .TE_B(_200_),
    .Z(\mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__ebufn_2 _707_ (.A(\mux_left_ipin_1.INVTX1_2_.out ),
    .TE_B(_201_),
    .Z(\mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(ccff_head),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(chany_bottom_in[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(chany_bottom_in[10]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(chany_bottom_in[11]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(chany_bottom_in[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(chany_bottom_in[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(chany_bottom_in[14]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(chany_bottom_in[15]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(chany_bottom_in[16]),
    .X(net9));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(chany_bottom_in[17]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(chany_bottom_in[18]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(chany_bottom_in[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(chany_bottom_in[2]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input14 (.A(chany_bottom_in[3]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(chany_bottom_in[4]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(chany_bottom_in[5]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(chany_bottom_in[6]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(chany_bottom_in[7]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(chany_bottom_in[8]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(chany_bottom_in[9]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(chany_top_in[0]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(chany_top_in[10]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(chany_top_in[11]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(chany_top_in[12]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(chany_top_in[13]),
    .X(net25));
 sky130_fd_sc_hd__dlymetal6s2s_1 input26 (.A(chany_top_in[14]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(chany_top_in[15]),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(chany_top_in[16]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(chany_top_in[17]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(chany_top_in[18]),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(chany_top_in[1]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(chany_top_in[2]),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 input33 (.A(chany_top_in[3]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(chany_top_in[4]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(chany_top_in[5]),
    .X(net35));
 sky130_fd_sc_hd__dlymetal6s2s_1 input36 (.A(chany_top_in[6]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(chany_top_in[7]),
    .X(net37));
 sky130_fd_sc_hd__dlymetal6s2s_1 input38 (.A(chany_top_in[8]),
    .X(net38));
 sky130_fd_sc_hd__dlymetal6s2s_1 input39 (.A(chany_top_in[9]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(pReset),
    .X(net40));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(ccff_tail));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(chany_bottom_out[0]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(chany_bottom_out[10]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(chany_bottom_out[11]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(chany_bottom_out[12]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(chany_bottom_out[13]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(chany_bottom_out[14]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(chany_bottom_out[15]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(chany_bottom_out[16]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(chany_bottom_out[17]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(chany_bottom_out[18]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(chany_bottom_out[1]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(chany_bottom_out[2]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(chany_bottom_out[3]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(chany_bottom_out[4]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(chany_bottom_out[5]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(chany_bottom_out[6]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(chany_bottom_out[7]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(chany_bottom_out[8]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(chany_bottom_out[9]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(chany_top_out[0]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(chany_top_out[10]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(chany_top_out[11]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(chany_top_out[12]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(chany_top_out[13]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(chany_top_out[14]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(chany_top_out[15]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(chany_top_out[16]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(chany_top_out[17]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(chany_top_out[18]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(chany_top_out[1]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(chany_top_out[2]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(chany_top_out[3]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(chany_top_out[4]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(chany_top_out[5]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(chany_top_out[6]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(chany_top_out[7]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(chany_top_out[8]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(chany_top_out[9]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(right_grid_left_width_0_height_0_subtile_0__pin_I_11_));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(right_grid_left_width_0_height_0_subtile_0__pin_I_3_));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(right_grid_left_width_0_height_0_subtile_0__pin_I_7_));
 sky130_fd_sc_hd__conb_1 _583__91 (.HI(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__401__A (.DIODE(_067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__400__A (.DIODE(_067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__399__A (.DIODE(_067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__398__A (.DIODE(_067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__397__A (.DIODE(_067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__396__A (.DIODE(_067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__395__A (.DIODE(_067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__394__A (.DIODE(_067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__393__A (.DIODE(_067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__413__A (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__412__A (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__411__A (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__410__A (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__409__A (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__408__A (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__407__A (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__406__A (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__405__A (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__404__A (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__424__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__423__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__422__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__421__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__420__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__419__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__418__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__417__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__416__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__415__A (.DIODE(_069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__435__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__434__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__433__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__432__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__431__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__430__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__429__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__428__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__427__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__426__A (.DIODE(_070_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(ccff_head));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(chany_bottom_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(chany_bottom_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(chany_bottom_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(chany_bottom_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(chany_bottom_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(chany_bottom_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(chany_bottom_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(chany_bottom_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(chany_bottom_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(chany_bottom_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(chany_bottom_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(chany_bottom_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(chany_bottom_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(chany_bottom_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(chany_bottom_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(chany_bottom_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(chany_bottom_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(chany_bottom_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(chany_bottom_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(chany_top_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(chany_top_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(chany_top_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(chany_top_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(chany_top_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(chany_top_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(chany_top_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(chany_top_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(chany_top_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(chany_top_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(chany_top_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(chany_top_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(chany_top_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(chany_top_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(chany_top_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(chany_top_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(chany_top_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(chany_top_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(chany_top_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__468__D (.DIODE(\mem_left_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__335__A (.DIODE(\mem_left_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__333__A (.DIODE(\mem_left_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__331__A (.DIODE(\mem_left_ipin_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__467__D (.DIODE(\mem_left_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__340__A (.DIODE(\mem_left_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__338__A (.DIODE(\mem_left_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__336__A (.DIODE(\mem_left_ipin_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__475__D (.DIODE(\mem_left_ipin_0.DFFR_5_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__334__A (.DIODE(\mem_left_ipin_0.DFFR_5_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__474__D (.DIODE(\mem_left_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__327__A (.DIODE(\mem_left_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__323__A (.DIODE(\mem_left_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__319__A (.DIODE(\mem_left_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__478__D (.DIODE(\mem_right_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__316__A (.DIODE(\mem_right_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__312__A (.DIODE(\mem_right_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__308__A (.DIODE(\mem_right_ipin_0.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__486__D (.DIODE(\mem_right_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__303__A (.DIODE(\mem_right_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__299__A (.DIODE(\mem_right_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__295__A (.DIODE(\mem_right_ipin_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__484__D (.DIODE(\mem_right_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__304__A (.DIODE(\mem_right_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__300__A (.DIODE(\mem_right_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__296__A (.DIODE(\mem_right_ipin_1.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__482__D (.DIODE(\mem_right_ipin_1.DFFR_4_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__302__A (.DIODE(\mem_right_ipin_1.DFFR_4_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__493__D (.DIODE(\mem_right_ipin_1.DFFR_5_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__298__A (.DIODE(\mem_right_ipin_1.DFFR_5_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__492__D (.DIODE(\mem_right_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__291__A (.DIODE(\mem_right_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__287__A (.DIODE(\mem_right_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__283__A (.DIODE(\mem_right_ipin_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__491__D (.DIODE(\mem_right_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__293__A (.DIODE(\mem_right_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__289__A (.DIODE(\mem_right_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__285__A (.DIODE(\mem_right_ipin_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__490__D (.DIODE(\mem_right_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__292__A (.DIODE(\mem_right_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__288__A (.DIODE(\mem_right_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__284__A (.DIODE(\mem_right_ipin_2.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__498__D (.DIODE(\mem_right_ipin_3.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__279__A (.DIODE(\mem_right_ipin_3.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__275__A (.DIODE(\mem_right_ipin_3.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__271__A (.DIODE(\mem_right_ipin_3.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__496__D (.DIODE(\mem_right_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__280__A (.DIODE(\mem_right_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__276__A (.DIODE(\mem_right_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__272__A (.DIODE(\mem_right_ipin_3.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__504__D (.DIODE(\mem_right_ipin_4.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__267__A (.DIODE(\mem_right_ipin_4.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__263__A (.DIODE(\mem_right_ipin_4.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__259__A (.DIODE(\mem_right_ipin_4.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__502__D (.DIODE(\mem_right_ipin_4.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__268__A (.DIODE(\mem_right_ipin_4.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__264__A (.DIODE(\mem_right_ipin_4.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__260__A (.DIODE(\mem_right_ipin_4.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__510__D (.DIODE(\mem_right_ipin_5.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__255__A (.DIODE(\mem_right_ipin_5.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__251__A (.DIODE(\mem_right_ipin_5.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__247__A (.DIODE(\mem_right_ipin_5.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__508__D (.DIODE(\mem_right_ipin_5.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__256__A (.DIODE(\mem_right_ipin_5.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__252__A (.DIODE(\mem_right_ipin_5.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__248__A (.DIODE(\mem_right_ipin_5.DFFR_2_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__516__D (.DIODE(\mem_right_ipin_6.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__243__A (.DIODE(\mem_right_ipin_6.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__239__A (.DIODE(\mem_right_ipin_6.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__235__A (.DIODE(\mem_right_ipin_6.DFFR_0_.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__344__A (.DIODE(\mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__635__A (.DIODE(\mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__663__A (.DIODE(\mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__664__A (.DIODE(\mux_right_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__384__A (.DIODE(\mux_right_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__385__A (.DIODE(\mux_right_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(pReset));
 sky130_fd_sc_hd__diode_2 ANTENNA__529__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__528__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__527__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__526__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__525__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__524__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__523__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__522__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__521__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__520__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__519__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__518__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__517__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__516__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__515__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__514__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__513__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__512__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__511__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__510__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__509__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__508__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__507__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__506__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__505__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__504__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__503__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__502__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__501__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__500__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__499__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__498__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__497__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__496__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__495__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__494__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__493__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__492__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__491__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__490__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__489__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__488__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__487__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__486__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__485__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__484__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__483__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__482__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__481__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__480__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__479__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__478__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__477__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__476__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__475__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__474__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__473__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__472__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__471__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__470__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__469__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__468__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__467__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__466__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__465__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__464__CLK (.DIODE(prog_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__469__D (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__552__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__346__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__542__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__368__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__578__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__350__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__577__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__352__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__575__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__359__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__574__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__366__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__572__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__343__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__551__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__356__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__550__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__389__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__548__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__370__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__547__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__375__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__546__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__348__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__545__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__354__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__544__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__382__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__543__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__361__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__571__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__347__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__561__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__367__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__560__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__390__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__559__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__342__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__558__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__357__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__556__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__364__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__555__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__371__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__570__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__355__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__569__A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__388__A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__567__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__369__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__566__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__374__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__565__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__349__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__447__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__436__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__391__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_output41_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__226__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_output43_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_output52_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_output54_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_output55_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_output56_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_output57_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_output62_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net79));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_405 ();
endmodule

