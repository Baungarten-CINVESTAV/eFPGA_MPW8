magic
tech sky130A
magscale 1 2
timestamp 1672422468
<< viali >>
rect 36829 37417 36863 37451
rect 23305 37349 23339 37383
rect 3985 37281 4019 37315
rect 6837 37281 6871 37315
rect 9321 37281 9355 37315
rect 10057 37281 10091 37315
rect 13737 37281 13771 37315
rect 14289 37281 14323 37315
rect 20821 37281 20855 37315
rect 21465 37281 21499 37315
rect 22017 37281 22051 37315
rect 24777 37281 24811 37315
rect 1685 37213 1719 37247
rect 2697 37213 2731 37247
rect 4905 37213 4939 37247
rect 6009 37213 6043 37247
rect 6653 37213 6687 37247
rect 8125 37213 8159 37247
rect 9873 37213 9907 37247
rect 13461 37213 13495 37247
rect 15209 37213 15243 37247
rect 17141 37213 17175 37247
rect 18429 37213 18463 37247
rect 20361 37213 20395 37247
rect 22293 37213 22327 37247
rect 23489 37213 23523 37247
rect 25329 37213 25363 37247
rect 26617 37213 26651 37247
rect 27169 37213 27203 37247
rect 28457 37213 28491 37247
rect 30389 37213 30423 37247
rect 32321 37213 32355 37247
rect 33609 37213 33643 37247
rect 35541 37213 35575 37247
rect 36645 37213 36679 37247
rect 37473 37213 37507 37247
rect 1777 37077 1811 37111
rect 2881 37077 2915 37111
rect 4721 37077 4755 37111
rect 5457 37077 5491 37111
rect 7941 37077 7975 37111
rect 15025 37077 15059 37111
rect 16957 37077 16991 37111
rect 18245 37077 18279 37111
rect 20177 37077 20211 37111
rect 25421 37077 25455 37111
rect 27353 37077 27387 37111
rect 28641 37077 28675 37111
rect 30573 37077 30607 37111
rect 32505 37077 32539 37111
rect 33793 37077 33827 37111
rect 34989 37077 35023 37111
rect 35725 37077 35759 37111
rect 37657 37077 37691 37111
rect 2421 36873 2455 36907
rect 6561 36873 6595 36907
rect 10517 36873 10551 36907
rect 23213 36873 23247 36907
rect 27353 36873 27387 36907
rect 34989 36873 35023 36907
rect 36461 36873 36495 36907
rect 38209 36873 38243 36907
rect 1685 36805 1719 36839
rect 3065 36805 3099 36839
rect 2605 36737 2639 36771
rect 6745 36737 6779 36771
rect 10701 36737 10735 36771
rect 11713 36737 11747 36771
rect 27169 36737 27203 36771
rect 34897 36737 34931 36771
rect 38025 36737 38059 36771
rect 11989 36669 12023 36703
rect 1869 36601 1903 36635
rect 35541 36533 35575 36567
rect 11621 36329 11655 36363
rect 38209 36329 38243 36363
rect 37565 36261 37599 36295
rect 1869 36125 1903 36159
rect 37381 36125 37415 36159
rect 38025 36125 38059 36159
rect 1685 35989 1719 36023
rect 29561 35785 29595 35819
rect 29377 35649 29411 35683
rect 38025 35581 38059 35615
rect 38301 35581 38335 35615
rect 38301 35241 38335 35275
rect 2421 34697 2455 34731
rect 1869 34561 1903 34595
rect 2513 34561 2547 34595
rect 3065 34493 3099 34527
rect 1685 34357 1719 34391
rect 37473 33473 37507 33507
rect 38025 33473 38059 33507
rect 38209 33337 38243 33371
rect 27353 32521 27387 32555
rect 1869 32385 1903 32419
rect 27169 32385 27203 32419
rect 38025 32317 38059 32351
rect 38301 32317 38335 32351
rect 1685 32181 1719 32215
rect 27905 32181 27939 32215
rect 38301 31977 38335 32011
rect 2513 30889 2547 30923
rect 27353 30889 27387 30923
rect 2329 30685 2363 30719
rect 2973 30685 3007 30719
rect 27169 30685 27203 30719
rect 27813 30685 27847 30719
rect 1685 30617 1719 30651
rect 1869 30617 1903 30651
rect 1685 30345 1719 30379
rect 30205 30209 30239 30243
rect 30849 30209 30883 30243
rect 37565 30209 37599 30243
rect 38209 30209 38243 30243
rect 30389 30073 30423 30107
rect 38117 30005 38151 30039
rect 23121 29529 23155 29563
rect 23029 29461 23063 29495
rect 23673 29461 23707 29495
rect 1685 29121 1719 29155
rect 1869 28985 1903 29019
rect 19993 28713 20027 28747
rect 1593 28645 1627 28679
rect 15577 28509 15611 28543
rect 20085 28509 20119 28543
rect 15669 28373 15703 28407
rect 20637 28373 20671 28407
rect 19257 28169 19291 28203
rect 25605 28169 25639 28203
rect 26341 28169 26375 28203
rect 18429 28101 18463 28135
rect 18521 28033 18555 28067
rect 19349 28033 19383 28067
rect 22201 28033 22235 28067
rect 26157 28033 26191 28067
rect 28549 28033 28583 28067
rect 37565 28033 37599 28067
rect 38209 28033 38243 28067
rect 28457 27897 28491 27931
rect 38025 27897 38059 27931
rect 22109 27829 22143 27863
rect 14841 27421 14875 27455
rect 32413 27421 32447 27455
rect 14933 27285 14967 27319
rect 18705 27285 18739 27319
rect 32321 27285 32355 27319
rect 1869 26945 1903 26979
rect 38025 26877 38059 26911
rect 38301 26877 38335 26911
rect 1685 26741 1719 26775
rect 38301 26537 38335 26571
rect 7205 25449 7239 25483
rect 9137 25449 9171 25483
rect 1593 25245 1627 25279
rect 1869 25245 1903 25279
rect 7389 25245 7423 25279
rect 9321 25245 9355 25279
rect 7849 25109 7883 25143
rect 9781 25109 9815 25143
rect 1593 24905 1627 24939
rect 38025 24701 38059 24735
rect 38301 24701 38335 24735
rect 38301 24361 38335 24395
rect 1593 23613 1627 23647
rect 1869 23613 1903 23647
rect 23857 23273 23891 23307
rect 1593 23205 1627 23239
rect 23397 23069 23431 23103
rect 23305 22933 23339 22967
rect 38025 22593 38059 22627
rect 38209 22457 38243 22491
rect 23581 22049 23615 22083
rect 23029 21981 23063 22015
rect 22937 21845 22971 21879
rect 6929 21641 6963 21675
rect 25697 21641 25731 21675
rect 32781 21641 32815 21675
rect 1869 21505 1903 21539
rect 7113 21505 7147 21539
rect 25605 21505 25639 21539
rect 32597 21505 32631 21539
rect 33241 21505 33275 21539
rect 38025 21505 38059 21539
rect 1685 21301 1719 21335
rect 7665 21301 7699 21335
rect 24961 21301 24995 21335
rect 38209 21301 38243 21335
rect 1777 21097 1811 21131
rect 1961 20893 1995 20927
rect 24777 20893 24811 20927
rect 22109 20757 22143 20791
rect 24685 20757 24719 20791
rect 22293 20417 22327 20451
rect 22937 20417 22971 20451
rect 24133 20417 24167 20451
rect 24777 20417 24811 20451
rect 25421 20417 25455 20451
rect 24593 20349 24627 20383
rect 23121 20281 23155 20315
rect 22385 20213 22419 20247
rect 23673 20213 23707 20247
rect 25329 20213 25363 20247
rect 26065 20009 26099 20043
rect 24869 19941 24903 19975
rect 23581 19873 23615 19907
rect 25421 19873 25455 19907
rect 21649 19805 21683 19839
rect 22293 19805 22327 19839
rect 23765 19805 23799 19839
rect 26157 19805 26191 19839
rect 1685 19737 1719 19771
rect 25329 19737 25363 19771
rect 1777 19669 1811 19703
rect 22201 19669 22235 19703
rect 23121 19669 23155 19703
rect 26709 19669 26743 19703
rect 1685 19465 1719 19499
rect 22661 19465 22695 19499
rect 24041 19397 24075 19431
rect 24133 19397 24167 19431
rect 24685 19397 24719 19431
rect 9321 19329 9355 19363
rect 9413 19329 9447 19363
rect 20821 19329 20855 19363
rect 21281 19329 21315 19363
rect 22201 19329 22235 19363
rect 25881 19329 25915 19363
rect 25973 19329 26007 19363
rect 26525 19329 26559 19363
rect 26617 19329 26651 19363
rect 38025 19329 38059 19363
rect 22017 19261 22051 19295
rect 23857 19261 23891 19295
rect 25145 19261 25179 19295
rect 25329 19261 25363 19295
rect 21373 19125 21407 19159
rect 27261 19125 27295 19159
rect 27721 19125 27755 19159
rect 38209 19125 38243 19159
rect 19717 18921 19751 18955
rect 22109 18921 22143 18955
rect 28273 18853 28307 18887
rect 21649 18785 21683 18819
rect 22661 18785 22695 18819
rect 23765 18785 23799 18819
rect 25145 18785 25179 18819
rect 27721 18785 27755 18819
rect 10149 18717 10183 18751
rect 10793 18717 10827 18751
rect 20821 18717 20855 18751
rect 21465 18717 21499 18751
rect 25329 18717 25363 18751
rect 25881 18717 25915 18751
rect 25973 18717 26007 18751
rect 26617 18717 26651 18751
rect 27261 18717 27295 18751
rect 10241 18649 10275 18683
rect 22753 18649 22787 18683
rect 23305 18649 23339 18683
rect 17601 18581 17635 18615
rect 20269 18581 20303 18615
rect 20913 18581 20947 18615
rect 24685 18581 24719 18615
rect 26525 18581 26559 18615
rect 27169 18581 27203 18615
rect 28917 18581 28951 18615
rect 17509 18309 17543 18343
rect 17601 18309 17635 18343
rect 19441 18309 19475 18343
rect 21373 18309 21407 18343
rect 22569 18309 22603 18343
rect 23397 18309 23431 18343
rect 27813 18309 27847 18343
rect 28365 18309 28399 18343
rect 1869 18241 1903 18275
rect 18705 18241 18739 18275
rect 20453 18241 20487 18275
rect 21281 18241 21315 18275
rect 24501 18241 24535 18275
rect 25237 18241 25271 18275
rect 26433 18241 26467 18275
rect 18153 18173 18187 18207
rect 19901 18173 19935 18207
rect 22661 18173 22695 18207
rect 23305 18173 23339 18207
rect 23949 18173 23983 18207
rect 26617 18173 26651 18207
rect 27169 18173 27203 18207
rect 18797 18105 18831 18139
rect 22109 18105 22143 18139
rect 25421 18105 25455 18139
rect 1685 18037 1719 18071
rect 20545 18037 20579 18071
rect 24501 18037 24535 18071
rect 25973 18037 26007 18071
rect 29009 18037 29043 18071
rect 29469 18037 29503 18071
rect 17141 17833 17175 17867
rect 22477 17833 22511 17867
rect 23397 17833 23431 17867
rect 29745 17833 29779 17867
rect 17785 17697 17819 17731
rect 24041 17697 24075 17731
rect 28733 17697 28767 17731
rect 17049 17629 17083 17663
rect 20269 17629 20303 17663
rect 22385 17629 22419 17663
rect 23857 17629 23891 17663
rect 26065 17629 26099 17663
rect 26893 17629 26927 17663
rect 27537 17629 27571 17663
rect 28181 17629 28215 17663
rect 28825 17629 28859 17663
rect 18797 17561 18831 17595
rect 20821 17561 20855 17595
rect 20913 17561 20947 17595
rect 21465 17561 21499 17595
rect 24961 17561 24995 17595
rect 25053 17561 25087 17595
rect 25605 17561 25639 17595
rect 26801 17561 26835 17595
rect 18245 17493 18279 17527
rect 19533 17493 19567 17527
rect 20177 17493 20211 17527
rect 26157 17493 26191 17527
rect 27445 17493 27479 17527
rect 28089 17493 28123 17527
rect 23305 17289 23339 17323
rect 25789 17289 25823 17323
rect 19533 17221 19567 17255
rect 22109 17221 22143 17255
rect 22201 17221 22235 17255
rect 22753 17221 22787 17255
rect 24869 17221 24903 17255
rect 29653 17221 29687 17255
rect 16313 17153 16347 17187
rect 16865 17153 16899 17187
rect 19993 17153 20027 17187
rect 20637 17153 20671 17187
rect 21281 17153 21315 17187
rect 23213 17153 23247 17187
rect 26249 17153 26283 17187
rect 26433 17153 26467 17187
rect 27169 17153 27203 17187
rect 27997 17153 28031 17187
rect 28641 17153 28675 17187
rect 18981 17085 19015 17119
rect 24685 17085 24719 17119
rect 24961 17085 24995 17119
rect 38025 17085 38059 17119
rect 38301 17085 38335 17119
rect 17785 17017 17819 17051
rect 20085 17017 20119 17051
rect 29101 17017 29135 17051
rect 16957 16949 16991 16983
rect 18337 16949 18371 16983
rect 20729 16949 20763 16983
rect 21373 16949 21407 16983
rect 27261 16949 27295 16983
rect 27905 16949 27939 16983
rect 28549 16949 28583 16983
rect 17049 16745 17083 16779
rect 17693 16745 17727 16779
rect 21557 16745 21591 16779
rect 22201 16745 22235 16779
rect 38301 16745 38335 16779
rect 18153 16677 18187 16711
rect 22845 16677 22879 16711
rect 29101 16677 29135 16711
rect 19441 16609 19475 16643
rect 23581 16609 23615 16643
rect 24685 16609 24719 16643
rect 24961 16609 24995 16643
rect 26801 16609 26835 16643
rect 27353 16609 27387 16643
rect 27813 16609 27847 16643
rect 28549 16609 28583 16643
rect 29745 16609 29779 16643
rect 18705 16541 18739 16575
rect 20913 16541 20947 16575
rect 23397 16541 23431 16575
rect 27997 16541 28031 16575
rect 28641 16541 28675 16575
rect 19993 16473 20027 16507
rect 20085 16473 20119 16507
rect 21005 16473 21039 16507
rect 22293 16473 22327 16507
rect 24777 16473 24811 16507
rect 25789 16473 25823 16507
rect 26709 16473 26743 16507
rect 18797 16405 18831 16439
rect 24041 16405 24075 16439
rect 30297 16405 30331 16439
rect 15117 16133 15151 16167
rect 17049 16133 17083 16167
rect 17601 16133 17635 16167
rect 18337 16133 18371 16167
rect 20361 16133 20395 16167
rect 22661 16133 22695 16167
rect 23213 16133 23247 16167
rect 23857 16133 23891 16167
rect 25421 16133 25455 16167
rect 27353 16133 27387 16167
rect 1869 16065 1903 16099
rect 15025 16065 15059 16099
rect 19533 16065 19567 16099
rect 20269 16065 20303 16099
rect 21097 16065 21131 16099
rect 28549 16065 28583 16099
rect 29193 16065 29227 16099
rect 29837 16065 29871 16099
rect 30481 16065 30515 16099
rect 38025 16065 38059 16099
rect 16957 15997 16991 16031
rect 18245 15997 18279 16031
rect 19441 15997 19475 16031
rect 22569 15997 22603 16031
rect 23765 15997 23799 16031
rect 24041 15997 24075 16031
rect 24869 15997 24903 16031
rect 25513 15997 25547 16031
rect 26065 15997 26099 16031
rect 27261 15997 27295 16031
rect 27537 15997 27571 16031
rect 29101 15997 29135 16031
rect 18797 15929 18831 15963
rect 29745 15929 29779 15963
rect 1685 15861 1719 15895
rect 2421 15861 2455 15895
rect 16221 15861 16255 15895
rect 20913 15861 20947 15895
rect 28457 15861 28491 15895
rect 30389 15861 30423 15895
rect 38209 15861 38243 15895
rect 22293 15657 22327 15691
rect 28733 15657 28767 15691
rect 31309 15657 31343 15691
rect 33609 15657 33643 15691
rect 38025 15657 38059 15691
rect 23121 15589 23155 15623
rect 24685 15589 24719 15623
rect 17233 15521 17267 15555
rect 17509 15521 17543 15555
rect 18705 15521 18739 15555
rect 19533 15521 19567 15555
rect 26341 15521 26375 15555
rect 26525 15521 26559 15555
rect 30481 15521 30515 15555
rect 20637 15453 20671 15487
rect 21465 15453 21499 15487
rect 22201 15453 22235 15487
rect 23305 15453 23339 15487
rect 23489 15453 23523 15487
rect 28181 15453 28215 15487
rect 28825 15453 28859 15487
rect 29929 15453 29963 15487
rect 30389 15453 30423 15487
rect 31401 15453 31435 15487
rect 33517 15453 33551 15487
rect 37841 15453 37875 15487
rect 16037 15385 16071 15419
rect 16221 15385 16255 15419
rect 17417 15385 17451 15419
rect 18061 15385 18095 15419
rect 18613 15385 18647 15419
rect 19625 15385 19659 15419
rect 20177 15385 20211 15419
rect 25237 15385 25271 15419
rect 25329 15385 25363 15419
rect 25881 15385 25915 15419
rect 27537 15385 27571 15419
rect 27629 15385 27663 15419
rect 15577 15317 15611 15351
rect 20729 15317 20763 15351
rect 21281 15317 21315 15351
rect 23949 15317 23983 15351
rect 26985 15317 27019 15351
rect 29837 15317 29871 15351
rect 18705 15113 18739 15147
rect 30757 15113 30791 15147
rect 17233 15045 17267 15079
rect 19441 15045 19475 15079
rect 20361 15045 20395 15079
rect 23397 15045 23431 15079
rect 23489 15045 23523 15079
rect 24593 15045 24627 15079
rect 25237 15045 25271 15079
rect 27445 15045 27479 15079
rect 27537 15045 27571 15079
rect 14749 14977 14783 15011
rect 16129 14977 16163 15011
rect 18797 14977 18831 15011
rect 22201 14977 22235 15011
rect 25697 14977 25731 15011
rect 26525 14977 26559 15011
rect 28089 14977 28123 15011
rect 28549 14977 28583 15011
rect 28733 14977 28767 15011
rect 31401 14977 31435 15011
rect 15577 14909 15611 14943
rect 17141 14909 17175 14943
rect 19349 14909 19383 14943
rect 21097 14909 21131 14943
rect 24685 14909 24719 14943
rect 25881 14909 25915 14943
rect 30113 14909 30147 14943
rect 30297 14909 30331 14943
rect 14657 14841 14691 14875
rect 17693 14841 17727 14875
rect 22937 14841 22971 14875
rect 24133 14841 24167 14875
rect 26341 14841 26375 14875
rect 31493 14841 31527 14875
rect 16221 14773 16255 14807
rect 22293 14773 22327 14807
rect 29009 14773 29043 14807
rect 29653 14773 29687 14807
rect 9229 14569 9263 14603
rect 15117 14569 15151 14603
rect 22201 14569 22235 14603
rect 30481 14569 30515 14603
rect 31769 14569 31803 14603
rect 32321 14569 32355 14603
rect 13737 14501 13771 14535
rect 16221 14501 16255 14535
rect 23121 14501 23155 14535
rect 27905 14501 27939 14535
rect 14565 14433 14599 14467
rect 23581 14433 23615 14467
rect 25237 14433 25271 14467
rect 26433 14433 26467 14467
rect 31125 14433 31159 14467
rect 1593 14365 1627 14399
rect 1869 14365 1903 14399
rect 9321 14365 9355 14399
rect 16865 14365 16899 14399
rect 17509 14365 17543 14399
rect 19441 14365 19475 14399
rect 20269 14365 20303 14399
rect 22109 14365 22143 14399
rect 23765 14365 23799 14399
rect 24593 14365 24627 14399
rect 25789 14365 25823 14399
rect 28365 14365 28399 14399
rect 28551 14365 28585 14399
rect 29193 14365 29227 14399
rect 29929 14365 29963 14399
rect 30389 14365 30423 14399
rect 31033 14365 31067 14399
rect 31861 14365 31895 14399
rect 15669 14297 15703 14331
rect 15761 14297 15795 14331
rect 16957 14297 16991 14331
rect 18245 14297 18279 14331
rect 18337 14297 18371 14331
rect 18889 14297 18923 14331
rect 20177 14297 20211 14331
rect 21005 14297 21039 14331
rect 21097 14297 21131 14331
rect 21649 14297 21683 14331
rect 25145 14297 25179 14331
rect 26525 14297 26559 14331
rect 27445 14297 27479 14331
rect 29837 14297 29871 14331
rect 32873 14297 32907 14331
rect 17601 14229 17635 14263
rect 19533 14229 19567 14263
rect 29101 14229 29135 14263
rect 1593 14025 1627 14059
rect 14013 14025 14047 14059
rect 14565 14025 14599 14059
rect 16221 14025 16255 14059
rect 26341 14025 26375 14059
rect 27169 14025 27203 14059
rect 32413 14025 32447 14059
rect 38117 14025 38151 14059
rect 13461 13957 13495 13991
rect 17601 13957 17635 13991
rect 18337 13957 18371 13991
rect 18889 13957 18923 13991
rect 20269 13957 20303 13991
rect 20913 13957 20947 13991
rect 23857 13957 23891 13991
rect 23949 13957 23983 13991
rect 25053 13957 25087 13991
rect 28365 13957 28399 13991
rect 28457 13957 28491 13991
rect 31217 13957 31251 13991
rect 16129 13889 16163 13923
rect 17049 13889 17083 13923
rect 17509 13889 17543 13923
rect 19441 13889 19475 13923
rect 22017 13889 22051 13923
rect 22845 13889 22879 13923
rect 27813 13889 27847 13923
rect 29653 13889 29687 13923
rect 30113 13889 30147 13923
rect 32505 13889 32539 13923
rect 37565 13889 37599 13923
rect 38301 13889 38335 13923
rect 15117 13821 15151 13855
rect 16957 13821 16991 13855
rect 18245 13821 18279 13855
rect 19533 13821 19567 13855
rect 20821 13821 20855 13855
rect 22109 13821 22143 13855
rect 23673 13821 23707 13855
rect 24501 13821 24535 13855
rect 25145 13821 25179 13855
rect 25697 13821 25731 13855
rect 25881 13821 25915 13855
rect 27629 13821 27663 13855
rect 30205 13821 30239 13855
rect 31125 13821 31159 13855
rect 32965 13821 32999 13855
rect 21373 13753 21407 13787
rect 28917 13753 28951 13787
rect 31677 13753 31711 13787
rect 15577 13685 15611 13719
rect 22753 13685 22787 13719
rect 29561 13685 29595 13719
rect 13737 13481 13771 13515
rect 14749 13481 14783 13515
rect 31033 13481 31067 13515
rect 31677 13481 31711 13515
rect 15945 13413 15979 13447
rect 20085 13413 20119 13447
rect 12633 13345 12667 13379
rect 17969 13345 18003 13379
rect 19533 13345 19567 13379
rect 20821 13345 20855 13379
rect 21189 13345 21223 13379
rect 22293 13345 22327 13379
rect 23305 13345 23339 13379
rect 24869 13345 24903 13379
rect 32965 13345 32999 13379
rect 15209 13277 15243 13311
rect 15853 13277 15887 13311
rect 16497 13277 16531 13311
rect 16589 13277 16623 13311
rect 24041 13277 24075 13311
rect 30481 13277 30515 13311
rect 31125 13277 31159 13311
rect 31769 13277 31803 13311
rect 32229 13277 32263 13311
rect 32873 13277 32907 13311
rect 13185 13209 13219 13243
rect 17325 13209 17359 13243
rect 18061 13209 18095 13243
rect 18613 13209 18647 13243
rect 19625 13209 19659 13243
rect 20913 13209 20947 13243
rect 23213 13209 23247 13243
rect 25697 13209 25731 13243
rect 25789 13209 25823 13243
rect 26617 13209 26651 13243
rect 26709 13209 26743 13243
rect 27629 13209 27663 13243
rect 28181 13209 28215 13243
rect 28273 13209 28307 13243
rect 29193 13209 29227 13243
rect 29837 13209 29871 13243
rect 29929 13209 29963 13243
rect 32321 13209 32355 13243
rect 15301 13141 15335 13175
rect 17233 13141 17267 13175
rect 23949 13141 23983 13175
rect 13369 12937 13403 12971
rect 14473 12937 14507 12971
rect 24869 12937 24903 12971
rect 30113 12937 30147 12971
rect 32413 12937 32447 12971
rect 12817 12869 12851 12903
rect 15669 12869 15703 12903
rect 15761 12869 15795 12903
rect 16313 12869 16347 12903
rect 17969 12869 18003 12903
rect 19165 12869 19199 12903
rect 20821 12869 20855 12903
rect 20913 12869 20947 12903
rect 21465 12869 21499 12903
rect 22201 12869 22235 12903
rect 23673 12869 23707 12903
rect 23765 12869 23799 12903
rect 25973 12869 26007 12903
rect 26065 12869 26099 12903
rect 27721 12869 27755 12903
rect 27813 12869 27847 12903
rect 32965 12869 32999 12903
rect 1869 12801 1903 12835
rect 14933 12801 14967 12835
rect 17141 12801 17175 12835
rect 24961 12801 24995 12835
rect 28365 12801 28399 12835
rect 29009 12801 29043 12835
rect 29653 12799 29687 12833
rect 30941 12801 30975 12835
rect 31585 12801 31619 12835
rect 32505 12801 32539 12835
rect 17877 12733 17911 12767
rect 19073 12733 19107 12767
rect 20085 12733 20119 12767
rect 22109 12733 22143 12767
rect 23029 12733 23063 12767
rect 23949 12733 23983 12767
rect 25789 12733 25823 12767
rect 29561 12733 29595 12767
rect 30849 12733 30883 12767
rect 13921 12665 13955 12699
rect 18429 12665 18463 12699
rect 1685 12597 1719 12631
rect 15025 12597 15059 12631
rect 17233 12597 17267 12631
rect 28917 12597 28951 12631
rect 31493 12597 31527 12631
rect 37933 12597 37967 12631
rect 29837 12393 29871 12427
rect 31769 12393 31803 12427
rect 14565 12325 14599 12359
rect 27169 12325 27203 12359
rect 31125 12325 31159 12359
rect 32965 12325 32999 12359
rect 12633 12257 12667 12291
rect 17049 12257 17083 12291
rect 18153 12257 18187 12291
rect 20453 12257 20487 12291
rect 21189 12257 21223 12291
rect 22017 12257 22051 12291
rect 23121 12257 23155 12291
rect 23765 12257 23799 12291
rect 25237 12257 25271 12291
rect 26157 12257 26191 12291
rect 27721 12257 27755 12291
rect 29101 12257 29135 12291
rect 32413 12257 32447 12291
rect 12081 12189 12115 12223
rect 14473 12189 14507 12223
rect 15117 12189 15151 12223
rect 15945 12189 15979 12223
rect 16405 12189 16439 12223
rect 18797 12189 18831 12223
rect 19809 12189 19843 12223
rect 29929 12189 29963 12223
rect 30389 12189 30423 12223
rect 31217 12189 31251 12223
rect 31677 12189 31711 12223
rect 32505 12189 32539 12223
rect 13737 12121 13771 12155
rect 16957 12121 16991 12155
rect 18245 12121 18279 12155
rect 20361 12121 20395 12155
rect 21281 12121 21315 12155
rect 23673 12121 23707 12155
rect 24593 12121 24627 12155
rect 25145 12121 25179 12155
rect 26433 12121 26467 12155
rect 26525 12121 26559 12155
rect 27629 12121 27663 12155
rect 28457 12121 28491 12155
rect 29009 12121 29043 12155
rect 30481 12121 30515 12155
rect 13185 12053 13219 12087
rect 15209 12053 15243 12087
rect 15853 12053 15887 12087
rect 37473 12053 37507 12087
rect 37933 12053 37967 12087
rect 6561 11849 6595 11883
rect 19901 11849 19935 11883
rect 22661 11849 22695 11883
rect 29101 11849 29135 11883
rect 31677 11849 31711 11883
rect 12909 11781 12943 11815
rect 15025 11781 15059 11815
rect 16129 11781 16163 11815
rect 17693 11781 17727 11815
rect 17785 11781 17819 11815
rect 18613 11781 18647 11815
rect 19165 11781 19199 11815
rect 21005 11781 21039 11815
rect 21097 11781 21131 11815
rect 23673 11781 23707 11815
rect 23765 11781 23799 11815
rect 24869 11781 24903 11815
rect 24961 11781 24995 11815
rect 26341 11781 26375 11815
rect 27169 11781 27203 11815
rect 27721 11781 27755 11815
rect 31033 11781 31067 11815
rect 5917 11713 5951 11747
rect 12357 11713 12391 11747
rect 13369 11713 13403 11747
rect 14289 11713 14323 11747
rect 15117 11713 15151 11747
rect 19809 11713 19843 11747
rect 22201 11713 22235 11747
rect 28365 11713 28399 11747
rect 29193 11713 29227 11747
rect 29837 11713 29871 11747
rect 30481 11713 30515 11747
rect 31125 11713 31159 11747
rect 31769 11713 31803 11747
rect 37565 11713 37599 11747
rect 38209 11713 38243 11747
rect 13461 11645 13495 11679
rect 16221 11645 16255 11679
rect 18521 11645 18555 11679
rect 20453 11645 20487 11679
rect 22017 11645 22051 11679
rect 26433 11645 26467 11679
rect 27813 11645 27847 11679
rect 30389 11645 30423 11679
rect 32965 11645 32999 11679
rect 15669 11577 15703 11611
rect 17233 11577 17267 11611
rect 23213 11577 23247 11611
rect 24409 11577 24443 11611
rect 25881 11577 25915 11611
rect 28457 11577 28491 11611
rect 38025 11577 38059 11611
rect 5733 11509 5767 11543
rect 14381 11509 14415 11543
rect 29745 11509 29779 11543
rect 32413 11509 32447 11543
rect 33425 11509 33459 11543
rect 36921 11509 36955 11543
rect 12449 11305 12483 11339
rect 23949 11305 23983 11339
rect 27077 11305 27111 11339
rect 30481 11305 30515 11339
rect 31677 11305 31711 11339
rect 32229 11305 32263 11339
rect 15577 11237 15611 11271
rect 27721 11237 27755 11271
rect 29837 11237 29871 11271
rect 14381 11169 14415 11203
rect 16405 11169 16439 11203
rect 17049 11169 17083 11203
rect 17693 11169 17727 11203
rect 18245 11169 18279 11203
rect 18613 11169 18647 11203
rect 20269 11169 20303 11203
rect 22109 11169 22143 11203
rect 25237 11169 25271 11203
rect 26157 11169 26191 11203
rect 11805 11101 11839 11135
rect 12357 11101 12391 11135
rect 13553 11101 13587 11135
rect 14289 11101 14323 11135
rect 21465 11101 21499 11135
rect 24041 11101 24075 11135
rect 28549 11101 28583 11135
rect 28641 11101 28675 11135
rect 29101 11101 29135 11135
rect 29929 11101 29963 11135
rect 30573 11101 30607 11135
rect 13645 11033 13679 11067
rect 15025 11033 15059 11067
rect 15117 11033 15151 11067
rect 16497 11033 16531 11067
rect 18337 11033 18371 11067
rect 19993 11033 20027 11067
rect 20085 11033 20119 11067
rect 22017 11033 22051 11067
rect 22661 11033 22695 11067
rect 23213 11033 23247 11067
rect 23305 11033 23339 11067
rect 24593 11033 24627 11067
rect 25145 11033 25179 11067
rect 25881 11033 25915 11067
rect 25973 11033 26007 11067
rect 27169 11033 27203 11067
rect 27905 11033 27939 11067
rect 31033 11033 31067 11067
rect 32781 11033 32815 11067
rect 35633 11033 35667 11067
rect 36093 11033 36127 11067
rect 36737 11033 36771 11067
rect 37289 11033 37323 11067
rect 38209 11033 38243 11067
rect 13093 10965 13127 10999
rect 35081 10965 35115 10999
rect 23765 10761 23799 10795
rect 29285 10761 29319 10795
rect 33333 10761 33367 10795
rect 15117 10693 15151 10727
rect 17325 10693 17359 10727
rect 18521 10693 18555 10727
rect 19073 10693 19107 10727
rect 19717 10693 19751 10727
rect 20913 10693 20947 10727
rect 21465 10693 21499 10727
rect 24777 10693 24811 10727
rect 24869 10693 24903 10727
rect 25421 10693 25455 10727
rect 25973 10693 26007 10727
rect 29929 10693 29963 10727
rect 1869 10625 1903 10659
rect 14473 10625 14507 10659
rect 16129 10625 16163 10659
rect 20269 10625 20303 10659
rect 22017 10625 22051 10659
rect 30021 10625 30055 10659
rect 33425 10625 33459 10659
rect 38025 10625 38059 10659
rect 15025 10557 15059 10591
rect 17233 10557 17267 10591
rect 18429 10557 18463 10591
rect 19625 10557 19659 10591
rect 20821 10557 20855 10591
rect 24225 10557 24259 10591
rect 26065 10557 26099 10591
rect 27537 10557 27571 10591
rect 27813 10557 27847 10591
rect 38301 10557 38335 10591
rect 14381 10489 14415 10523
rect 15577 10489 15611 10523
rect 17785 10489 17819 10523
rect 31585 10489 31619 10523
rect 34805 10489 34839 10523
rect 35449 10489 35483 10523
rect 36829 10489 36863 10523
rect 1685 10421 1719 10455
rect 13277 10421 13311 10455
rect 13829 10421 13863 10455
rect 16221 10421 16255 10455
rect 22280 10421 22314 10455
rect 30481 10421 30515 10455
rect 31033 10421 31067 10455
rect 32413 10421 32447 10455
rect 33885 10421 33919 10455
rect 36277 10421 36311 10455
rect 14657 10217 14691 10251
rect 18797 10217 18831 10251
rect 24685 10217 24719 10251
rect 29745 10217 29779 10251
rect 32045 10217 32079 10251
rect 36645 10217 36679 10251
rect 37657 10217 37691 10251
rect 38301 10217 38335 10251
rect 16681 10149 16715 10183
rect 22293 10149 22327 10183
rect 22937 10149 22971 10183
rect 28457 10149 28491 10183
rect 31401 10149 31435 10183
rect 15853 10081 15887 10115
rect 17233 10081 17267 10115
rect 17877 10081 17911 10115
rect 20821 10081 20855 10115
rect 23489 10081 23523 10115
rect 25697 10081 25731 10115
rect 13553 10013 13587 10047
rect 14749 10013 14783 10047
rect 16589 10013 16623 10047
rect 18889 10013 18923 10047
rect 19901 10013 19935 10047
rect 20545 10013 20579 10047
rect 24593 10013 24627 10047
rect 25421 10013 25455 10047
rect 27813 10013 27847 10047
rect 27905 10013 27939 10047
rect 28549 10013 28583 10047
rect 32137 10013 32171 10047
rect 32689 10013 32723 10047
rect 33241 10013 33275 10047
rect 33793 10013 33827 10047
rect 34253 10013 34287 10047
rect 15209 9945 15243 9979
rect 15761 9945 15795 9979
rect 17785 9945 17819 9979
rect 23404 9945 23438 9979
rect 29101 9945 29135 9979
rect 30297 9945 30331 9979
rect 30849 9945 30883 9979
rect 36001 9945 36035 9979
rect 37105 9945 37139 9979
rect 13001 9877 13035 9911
rect 13645 9877 13679 9911
rect 19993 9877 20027 9911
rect 27169 9877 27203 9911
rect 34989 9877 35023 9911
rect 35449 9877 35483 9911
rect 13829 9673 13863 9707
rect 4721 9605 4755 9639
rect 13277 9605 13311 9639
rect 14381 9605 14415 9639
rect 15761 9605 15795 9639
rect 17049 9605 17083 9639
rect 19073 9605 19107 9639
rect 19993 9605 20027 9639
rect 24041 9605 24075 9639
rect 36277 9605 36311 9639
rect 36829 9605 36863 9639
rect 4813 9537 4847 9571
rect 5365 9537 5399 9571
rect 14289 9537 14323 9571
rect 14933 9537 14967 9571
rect 16313 9537 16347 9571
rect 24501 9537 24535 9571
rect 15669 9469 15703 9503
rect 16957 9469 16991 9503
rect 17601 9469 17635 9503
rect 18889 9469 18923 9503
rect 19165 9469 19199 9503
rect 19717 9469 19751 9503
rect 22017 9469 22051 9503
rect 24777 9469 24811 9503
rect 26525 9469 26559 9503
rect 27169 9469 27203 9503
rect 28917 9469 28951 9503
rect 29193 9469 29227 9503
rect 29745 9469 29779 9503
rect 31401 9469 31435 9503
rect 33517 9469 33551 9503
rect 34069 9469 34103 9503
rect 35173 9469 35207 9503
rect 37473 9469 37507 9503
rect 34621 9401 34655 9435
rect 15025 9333 15059 9367
rect 21465 9333 21499 9367
rect 22280 9333 22314 9367
rect 30205 9333 30239 9367
rect 30757 9333 30791 9367
rect 32321 9333 32355 9367
rect 32873 9333 32907 9367
rect 35725 9333 35759 9367
rect 38209 9333 38243 9367
rect 15025 9129 15059 9163
rect 23489 9129 23523 9163
rect 24685 9129 24719 9163
rect 25329 9129 25363 9163
rect 26138 9129 26172 9163
rect 35541 9129 35575 9163
rect 1869 9061 1903 9095
rect 16957 9061 16991 9095
rect 15669 8993 15703 9027
rect 16313 8993 16347 9027
rect 19809 8993 19843 9027
rect 21189 8993 21223 9027
rect 22937 8993 22971 9027
rect 13737 8925 13771 8959
rect 14289 8925 14323 8959
rect 14933 8925 14967 8959
rect 16865 8925 16899 8959
rect 17693 8925 17727 8959
rect 20913 8925 20947 8959
rect 23397 8925 23431 8959
rect 24777 8925 24811 8959
rect 25421 8925 25455 8959
rect 25881 8925 25915 8959
rect 27905 8925 27939 8959
rect 31769 8925 31803 8959
rect 1685 8857 1719 8891
rect 15754 8857 15788 8891
rect 18153 8857 18187 8891
rect 18705 8857 18739 8891
rect 18797 8857 18831 8891
rect 19533 8857 19567 8891
rect 19625 8857 19659 8891
rect 29745 8857 29779 8891
rect 31493 8857 31527 8891
rect 36001 8857 36035 8891
rect 38209 8857 38243 8891
rect 14381 8789 14415 8823
rect 17601 8789 17635 8823
rect 28365 8789 28399 8823
rect 28917 8789 28951 8823
rect 32321 8789 32355 8823
rect 32873 8789 32907 8823
rect 33333 8789 33367 8823
rect 33885 8789 33919 8823
rect 34897 8789 34931 8823
rect 36553 8789 36587 8823
rect 37197 8789 37231 8823
rect 37657 8789 37691 8823
rect 1685 8585 1719 8619
rect 10885 8585 10919 8619
rect 19717 8585 19751 8619
rect 38117 8585 38151 8619
rect 14105 8517 14139 8551
rect 14657 8517 14691 8551
rect 15853 8517 15887 8551
rect 17049 8517 17083 8551
rect 18245 8517 18279 8551
rect 31125 8517 31159 8551
rect 10793 8449 10827 8483
rect 18797 8449 18831 8483
rect 22109 8449 22143 8483
rect 31401 8449 31435 8483
rect 35725 8449 35759 8483
rect 36185 8449 36219 8483
rect 37657 8449 37691 8483
rect 38301 8449 38335 8483
rect 13645 8381 13679 8415
rect 14749 8381 14783 8415
rect 15945 8381 15979 8415
rect 16957 8381 16991 8415
rect 18153 8381 18187 8415
rect 21189 8381 21223 8415
rect 21465 8381 21499 8415
rect 22385 8381 22419 8415
rect 23857 8381 23891 8415
rect 24501 8381 24535 8415
rect 25973 8381 26007 8415
rect 26249 8381 26283 8415
rect 27169 8381 27203 8415
rect 27445 8381 27479 8415
rect 29193 8381 29227 8415
rect 29653 8381 29687 8415
rect 32321 8381 32355 8415
rect 15393 8313 15427 8347
rect 17509 8313 17543 8347
rect 34529 8313 34563 8347
rect 35173 8313 35207 8347
rect 32965 8245 32999 8279
rect 33517 8245 33551 8279
rect 34069 8245 34103 8279
rect 36829 8245 36863 8279
rect 16221 8041 16255 8075
rect 17509 8041 17543 8075
rect 18153 8041 18187 8075
rect 18797 8041 18831 8075
rect 19809 8041 19843 8075
rect 27426 8041 27460 8075
rect 32597 8041 32631 8075
rect 33149 8041 33183 8075
rect 33701 8041 33735 8075
rect 34253 8041 34287 8075
rect 34897 8041 34931 8075
rect 35541 8041 35575 8075
rect 36553 8041 36587 8075
rect 37657 8041 37691 8075
rect 38209 8041 38243 8075
rect 15669 7973 15703 8007
rect 16865 7973 16899 8007
rect 28917 7973 28951 8007
rect 29745 7973 29779 8007
rect 30297 7973 30331 8007
rect 14657 7905 14691 7939
rect 31953 7905 31987 7939
rect 16129 7837 16163 7871
rect 16957 7837 16991 7871
rect 17601 7837 17635 7871
rect 18245 7837 18279 7871
rect 18705 7837 18739 7871
rect 19717 7837 19751 7871
rect 20361 7837 20395 7871
rect 21005 7837 21039 7871
rect 23029 7837 23063 7871
rect 24593 7837 24627 7871
rect 27169 7837 27203 7871
rect 30849 7837 30883 7871
rect 31401 7837 31435 7871
rect 14933 7769 14967 7803
rect 15025 7769 15059 7803
rect 22753 7769 22787 7803
rect 24869 7769 24903 7803
rect 20453 7701 20487 7735
rect 23489 7701 23523 7735
rect 26341 7701 26375 7735
rect 36001 7701 36035 7735
rect 37197 7701 37231 7735
rect 13737 7497 13771 7531
rect 15025 7497 15059 7531
rect 18613 7497 18647 7531
rect 19165 7497 19199 7531
rect 24501 7497 24535 7531
rect 28917 7497 28951 7531
rect 32413 7497 32447 7531
rect 33517 7497 33551 7531
rect 34069 7497 34103 7531
rect 34621 7497 34655 7531
rect 35173 7497 35207 7531
rect 35725 7497 35759 7531
rect 37473 7497 37507 7531
rect 15577 7429 15611 7463
rect 16129 7429 16163 7463
rect 17417 7429 17451 7463
rect 17509 7429 17543 7463
rect 21189 7429 21223 7463
rect 25973 7429 26007 7463
rect 30573 7429 30607 7463
rect 36737 7429 36771 7463
rect 1869 7361 1903 7395
rect 2513 7361 2547 7395
rect 13645 7361 13679 7395
rect 19073 7361 19107 7395
rect 21465 7361 21499 7395
rect 22017 7361 22051 7395
rect 26249 7361 26283 7395
rect 36829 7361 36863 7395
rect 16221 7293 16255 7327
rect 22293 7293 22327 7327
rect 23765 7293 23799 7327
rect 27169 7293 27203 7327
rect 27445 7293 27479 7327
rect 2329 7225 2363 7259
rect 16957 7225 16991 7259
rect 29469 7225 29503 7259
rect 31125 7225 31159 7259
rect 1685 7157 1719 7191
rect 19717 7157 19751 7191
rect 30021 7157 30055 7191
rect 31677 7157 31711 7191
rect 32873 7157 32907 7191
rect 38025 7157 38059 7191
rect 27261 6953 27295 6987
rect 28751 6953 28785 6987
rect 30002 6953 30036 6987
rect 31493 6953 31527 6987
rect 15301 6817 15335 6851
rect 15945 6817 15979 6851
rect 16589 6817 16623 6851
rect 18429 6817 18463 6851
rect 19533 6817 19567 6851
rect 20361 6817 20395 6851
rect 22845 6817 22879 6851
rect 24777 6817 24811 6851
rect 36553 6817 36587 6851
rect 6377 6749 6411 6783
rect 7021 6749 7055 6783
rect 16037 6749 16071 6783
rect 16681 6749 16715 6783
rect 17325 6749 17359 6783
rect 18521 6749 18555 6783
rect 19625 6749 19659 6783
rect 22385 6749 22419 6783
rect 23397 6749 23431 6783
rect 26525 6749 26559 6783
rect 29009 6749 29043 6783
rect 29745 6749 29779 6783
rect 33425 6749 33459 6783
rect 33517 6749 33551 6783
rect 34069 6749 34103 6783
rect 34161 6749 34195 6783
rect 36645 6749 36679 6783
rect 38209 6749 38243 6783
rect 14657 6681 14691 6715
rect 15209 6681 15243 6715
rect 17233 6681 17267 6715
rect 17785 6681 17819 6715
rect 22109 6681 22143 6715
rect 26249 6681 26283 6715
rect 32597 6681 32631 6715
rect 37657 6681 37691 6715
rect 6561 6613 6595 6647
rect 24041 6613 24075 6647
rect 32045 6613 32079 6647
rect 34897 6613 34931 6647
rect 35449 6613 35483 6647
rect 37105 6613 37139 6647
rect 17233 6409 17267 6443
rect 18521 6409 18555 6443
rect 24225 6409 24259 6443
rect 32689 6409 32723 6443
rect 33333 6409 33367 6443
rect 34621 6409 34655 6443
rect 35265 6409 35299 6443
rect 36645 6409 36679 6443
rect 22753 6341 22787 6375
rect 24961 6341 24995 6375
rect 28825 6341 28859 6375
rect 31309 6341 31343 6375
rect 33977 6341 34011 6375
rect 36001 6341 36035 6375
rect 17325 6273 17359 6307
rect 22477 6273 22511 6307
rect 30849 6273 30883 6307
rect 32781 6273 32815 6307
rect 33425 6273 33459 6307
rect 34069 6273 34103 6307
rect 34713 6273 34747 6307
rect 35357 6273 35391 6307
rect 36093 6273 36127 6307
rect 36737 6273 36771 6307
rect 38025 6273 38059 6307
rect 38301 6273 38335 6307
rect 15669 6205 15703 6239
rect 19717 6205 19751 6239
rect 19993 6205 20027 6239
rect 24685 6205 24719 6239
rect 30573 6205 30607 6239
rect 16313 6137 16347 6171
rect 21465 6137 21499 6171
rect 27169 6137 27203 6171
rect 27721 6137 27755 6171
rect 28273 6137 28307 6171
rect 13277 6069 13311 6103
rect 13921 6069 13955 6103
rect 14657 6069 14691 6103
rect 15209 6069 15243 6103
rect 17877 6069 17911 6103
rect 19073 6069 19107 6103
rect 26433 6069 26467 6103
rect 14565 5865 14599 5899
rect 16681 5865 16715 5899
rect 18889 5865 18923 5899
rect 21005 5865 21039 5899
rect 23765 5865 23799 5899
rect 32873 5865 32907 5899
rect 36277 5865 36311 5899
rect 17325 5797 17359 5831
rect 23213 5797 23247 5831
rect 29745 5797 29779 5831
rect 34989 5797 35023 5831
rect 15393 5729 15427 5763
rect 16037 5729 16071 5763
rect 26801 5729 26835 5763
rect 27445 5729 27479 5763
rect 28917 5729 28951 5763
rect 31217 5729 31251 5763
rect 31493 5729 31527 5763
rect 31953 5729 31987 5763
rect 37105 5729 37139 5763
rect 2881 5661 2915 5695
rect 13185 5661 13219 5695
rect 13737 5661 13771 5695
rect 14473 5661 14507 5695
rect 16773 5661 16807 5695
rect 17417 5661 17451 5695
rect 20269 5661 20303 5695
rect 21465 5661 21499 5695
rect 26341 5661 26375 5695
rect 29193 5661 29227 5695
rect 32965 5661 32999 5695
rect 33609 5661 33643 5695
rect 34161 5661 34195 5695
rect 34253 5661 34287 5695
rect 35081 5661 35115 5695
rect 35725 5661 35759 5695
rect 36369 5661 36403 5695
rect 37197 5661 37231 5695
rect 37841 5661 37875 5695
rect 15945 5593 15979 5627
rect 21741 5593 21775 5627
rect 26065 5593 26099 5627
rect 33517 5593 33551 5627
rect 35633 5593 35667 5627
rect 2789 5525 2823 5559
rect 18337 5525 18371 5559
rect 19717 5525 19751 5559
rect 24593 5525 24627 5559
rect 37749 5525 37783 5559
rect 10517 5321 10551 5355
rect 15025 5321 15059 5355
rect 22109 5321 22143 5355
rect 30573 5321 30607 5355
rect 13093 5253 13127 5287
rect 13737 5253 13771 5287
rect 23121 5253 23155 5287
rect 24409 5253 24443 5287
rect 26157 5253 26191 5287
rect 29837 5253 29871 5287
rect 33793 5253 33827 5287
rect 38025 5253 38059 5287
rect 38209 5253 38243 5287
rect 1869 5185 1903 5219
rect 2329 5185 2363 5219
rect 9965 5185 9999 5219
rect 11897 5185 11931 5219
rect 12357 5185 12391 5219
rect 13001 5185 13035 5219
rect 13829 5185 13863 5219
rect 14289 5185 14323 5219
rect 14933 5185 14967 5219
rect 15853 5185 15887 5219
rect 15945 5185 15979 5219
rect 17049 5185 17083 5219
rect 21465 5185 21499 5219
rect 24133 5185 24167 5219
rect 30113 5185 30147 5219
rect 31585 5185 31619 5219
rect 34621 5185 34655 5219
rect 34713 5185 34747 5219
rect 35357 5185 35391 5219
rect 36001 5185 36035 5219
rect 36645 5185 36679 5219
rect 18705 5117 18739 5151
rect 21189 5117 21223 5151
rect 28089 5117 28123 5151
rect 31677 5117 31711 5151
rect 34069 5117 34103 5151
rect 12449 5049 12483 5083
rect 35265 5049 35299 5083
rect 1685 4981 1719 5015
rect 9781 4981 9815 5015
rect 11805 4981 11839 5015
rect 14381 4981 14415 5015
rect 16865 4981 16899 5015
rect 17601 4981 17635 5015
rect 18153 4981 18187 5015
rect 19257 4981 19291 5015
rect 19717 4981 19751 5015
rect 22661 4981 22695 5015
rect 27169 4981 27203 5015
rect 32321 4981 32355 5015
rect 35909 4981 35943 5015
rect 36553 4981 36587 5015
rect 37565 4981 37599 5015
rect 12357 4777 12391 4811
rect 13645 4777 13679 4811
rect 14657 4777 14691 4811
rect 15301 4777 15335 4811
rect 22937 4777 22971 4811
rect 26801 4777 26835 4811
rect 31493 4777 31527 4811
rect 32216 4777 32250 4811
rect 13001 4709 13035 4743
rect 22385 4709 22419 4743
rect 23949 4709 23983 4743
rect 33701 4709 33735 4743
rect 37565 4709 37599 4743
rect 20637 4641 20671 4675
rect 24593 4641 24627 4675
rect 26065 4641 26099 4675
rect 28273 4641 28307 4675
rect 28549 4641 28583 4675
rect 29745 4641 29779 4675
rect 11805 4573 11839 4607
rect 12265 4573 12299 4607
rect 12909 4573 12943 4607
rect 13553 4573 13587 4607
rect 14565 4573 14599 4607
rect 15393 4573 15427 4607
rect 15853 4573 15887 4607
rect 16489 4567 16523 4601
rect 17141 4573 17175 4607
rect 19625 4573 19659 4607
rect 20177 4573 20211 4607
rect 23857 4573 23891 4607
rect 26341 4573 26375 4607
rect 31953 4573 31987 4607
rect 34345 4573 34379 4607
rect 35081 4573 35115 4607
rect 35725 4573 35759 4607
rect 36369 4573 36403 4607
rect 37013 4573 37047 4607
rect 37657 4573 37691 4607
rect 38117 4573 38151 4607
rect 11713 4505 11747 4539
rect 17233 4505 17267 4539
rect 20913 4505 20947 4539
rect 30021 4505 30055 4539
rect 36921 4505 36955 4539
rect 38209 4505 38243 4539
rect 15945 4437 15979 4471
rect 16589 4437 16623 4471
rect 18337 4437 18371 4471
rect 18797 4437 18831 4471
rect 29009 4437 29043 4471
rect 34161 4437 34195 4471
rect 34989 4437 35023 4471
rect 35633 4437 35667 4471
rect 36277 4437 36311 4471
rect 12909 4165 12943 4199
rect 14289 4165 14323 4199
rect 11161 4097 11195 4131
rect 11897 4097 11931 4131
rect 12449 4097 12483 4131
rect 13461 4097 13495 4131
rect 15301 4097 15335 4131
rect 16129 4097 16163 4131
rect 16221 4097 16255 4131
rect 17049 4097 17083 4131
rect 17141 4097 17175 4131
rect 17609 4097 17643 4131
rect 19717 4097 19751 4131
rect 22017 4097 22051 4131
rect 24225 4097 24259 4131
rect 26433 4097 26467 4131
rect 26525 4097 26559 4131
rect 31493 4097 31527 4131
rect 34713 4097 34747 4131
rect 35357 4097 35391 4131
rect 36001 4097 36035 4131
rect 36645 4097 36679 4131
rect 37657 4097 37691 4131
rect 38117 4097 38151 4131
rect 14197 4029 14231 4063
rect 14565 4029 14599 4063
rect 15393 4029 15427 4063
rect 17693 4029 17727 4063
rect 19993 4029 20027 4063
rect 22293 4029 22327 4063
rect 24501 4029 24535 4063
rect 27537 4029 27571 4063
rect 27813 4029 27847 4063
rect 29745 4029 29779 4063
rect 31217 4029 31251 4063
rect 32321 4029 32355 4063
rect 32597 4029 32631 4063
rect 37565 4029 37599 4063
rect 13553 3961 13587 3995
rect 19257 3961 19291 3995
rect 21465 3961 21499 3995
rect 23765 3961 23799 3995
rect 36553 3961 36587 3995
rect 18613 3893 18647 3927
rect 25973 3893 26007 3927
rect 29285 3893 29319 3927
rect 34069 3893 34103 3927
rect 34621 3893 34655 3927
rect 35265 3893 35299 3927
rect 35909 3893 35943 3927
rect 38209 3893 38243 3927
rect 2329 3689 2363 3723
rect 10609 3689 10643 3723
rect 11621 3689 11655 3723
rect 12265 3689 12299 3723
rect 13645 3689 13679 3723
rect 23213 3689 23247 3723
rect 29193 3689 29227 3723
rect 31953 3689 31987 3723
rect 34253 3689 34287 3723
rect 27537 3621 27571 3655
rect 29745 3621 29779 3655
rect 20545 3553 20579 3587
rect 25053 3553 25087 3587
rect 31493 3553 31527 3587
rect 33701 3553 33735 3587
rect 1869 3485 1903 3519
rect 12173 3485 12207 3519
rect 13553 3485 13587 3519
rect 14289 3485 14323 3519
rect 14565 3485 14599 3519
rect 17141 3485 17175 3519
rect 17601 3485 17635 3519
rect 17877 3485 17911 3519
rect 18521 3485 18555 3519
rect 23121 3485 23155 3519
rect 24041 3485 24075 3519
rect 29009 3485 29043 3519
rect 34345 3485 34379 3519
rect 35081 3485 35115 3519
rect 35725 3485 35759 3519
rect 36369 3485 36403 3519
rect 36829 3485 36863 3519
rect 38025 3485 38059 3519
rect 11161 3417 11195 3451
rect 15209 3417 15243 3451
rect 15945 3417 15979 3451
rect 16497 3417 16531 3451
rect 16589 3417 16623 3451
rect 19625 3417 19659 3451
rect 20821 3417 20855 3451
rect 22569 3417 22603 3451
rect 25329 3417 25363 3451
rect 27077 3417 27111 3451
rect 31217 3417 31251 3451
rect 33425 3417 33459 3451
rect 1685 3349 1719 3383
rect 13093 3349 13127 3383
rect 18613 3349 18647 3383
rect 19533 3349 19567 3383
rect 23857 3349 23891 3383
rect 28089 3349 28123 3383
rect 34989 3349 35023 3383
rect 35633 3349 35667 3383
rect 36277 3349 36311 3383
rect 37013 3349 37047 3383
rect 37565 3349 37599 3383
rect 38209 3349 38243 3383
rect 5089 3145 5123 3179
rect 11161 3145 11195 3179
rect 12541 3145 12575 3179
rect 15301 3145 15335 3179
rect 16957 3145 16991 3179
rect 21465 3145 21499 3179
rect 38209 3145 38243 3179
rect 10609 3077 10643 3111
rect 13369 3077 13403 3111
rect 17785 3077 17819 3111
rect 19993 3077 20027 3111
rect 24869 3077 24903 3111
rect 27905 3077 27939 3111
rect 29653 3077 29687 3111
rect 32597 3077 32631 3111
rect 37473 3077 37507 3111
rect 1869 3009 1903 3043
rect 2605 3009 2639 3043
rect 5273 3009 5307 3043
rect 11805 3009 11839 3043
rect 12449 3009 12483 3043
rect 13093 3009 13127 3043
rect 14013 3009 14047 3043
rect 15209 3009 15243 3043
rect 16221 3009 16255 3043
rect 17049 3009 17083 3043
rect 17509 3009 17543 3043
rect 19717 3009 19751 3043
rect 22017 3009 22051 3043
rect 24593 3009 24627 3043
rect 26617 3009 26651 3043
rect 27261 3009 27295 3043
rect 27445 3009 27479 3043
rect 29929 3009 29963 3043
rect 30665 3009 30699 3043
rect 31769 3009 31803 3043
rect 34713 3009 34747 3043
rect 35357 3009 35391 3043
rect 36001 3009 36035 3043
rect 36461 3009 36495 3043
rect 37657 3009 37691 3043
rect 14197 2941 14231 2975
rect 15945 2941 15979 2975
rect 22293 2941 22327 2975
rect 32321 2941 32355 2975
rect 19257 2873 19291 2907
rect 23765 2873 23799 2907
rect 31585 2873 31619 2907
rect 35817 2873 35851 2907
rect 1685 2805 1719 2839
rect 2421 2805 2455 2839
rect 3065 2805 3099 2839
rect 9689 2805 9723 2839
rect 11897 2805 11931 2839
rect 30481 2805 30515 2839
rect 34069 2805 34103 2839
rect 34621 2805 34655 2839
rect 35265 2805 35299 2839
rect 36645 2805 36679 2839
rect 10057 2601 10091 2635
rect 11161 2601 11195 2635
rect 12909 2601 12943 2635
rect 19717 2601 19751 2635
rect 22017 2601 22051 2635
rect 24593 2601 24627 2635
rect 29193 2601 29227 2635
rect 31493 2601 31527 2635
rect 9413 2533 9447 2567
rect 13461 2533 13495 2567
rect 18705 2533 18739 2567
rect 32321 2533 32355 2567
rect 2145 2465 2179 2499
rect 4077 2465 4111 2499
rect 17601 2465 17635 2499
rect 21465 2465 21499 2499
rect 23765 2465 23799 2499
rect 26065 2465 26099 2499
rect 29745 2465 29779 2499
rect 30021 2465 30055 2499
rect 33793 2465 33827 2499
rect 34069 2465 34103 2499
rect 37473 2465 37507 2499
rect 37749 2465 37783 2499
rect 2421 2397 2455 2431
rect 3433 2397 3467 2431
rect 4905 2397 4939 2431
rect 6561 2397 6595 2431
rect 9873 2397 9907 2431
rect 11989 2397 12023 2431
rect 14289 2397 14323 2431
rect 15485 2397 15519 2431
rect 16313 2397 16347 2431
rect 17417 2397 17451 2431
rect 18889 2397 18923 2431
rect 26341 2397 26375 2431
rect 27445 2397 27479 2431
rect 35173 2397 35207 2431
rect 35633 2397 35667 2431
rect 36645 2397 36679 2431
rect 9229 2329 9263 2363
rect 10609 2329 10643 2363
rect 13645 2329 13679 2363
rect 14565 2329 14599 2363
rect 21189 2329 21223 2363
rect 23489 2329 23523 2363
rect 27721 2329 27755 2363
rect 3249 2261 3283 2295
rect 4721 2261 4755 2295
rect 6745 2261 6779 2295
rect 8493 2261 8527 2295
rect 11805 2261 11839 2295
rect 15301 2261 15335 2295
rect 16129 2261 16163 2295
rect 16957 2261 16991 2295
rect 34989 2261 35023 2295
rect 35817 2261 35851 2295
rect 36829 2261 36863 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 36814 37448 36820 37460
rect 36775 37420 36820 37448
rect 36814 37408 36820 37420
rect 36872 37408 36878 37460
rect 17310 37340 17316 37392
rect 17368 37380 17374 37392
rect 23293 37383 23351 37389
rect 23293 37380 23305 37383
rect 17368 37352 23305 37380
rect 17368 37340 17374 37352
rect 23293 37349 23305 37352
rect 23339 37349 23351 37383
rect 23293 37343 23351 37349
rect 3973 37315 4031 37321
rect 3973 37312 3985 37315
rect 1688 37284 3985 37312
rect 1394 37204 1400 37256
rect 1452 37244 1458 37256
rect 1688 37253 1716 37284
rect 3973 37281 3985 37284
rect 4019 37281 4031 37315
rect 3973 37275 4031 37281
rect 6546 37272 6552 37324
rect 6604 37312 6610 37324
rect 6825 37315 6883 37321
rect 6825 37312 6837 37315
rect 6604 37284 6837 37312
rect 6604 37272 6610 37284
rect 6825 37281 6837 37284
rect 6871 37281 6883 37315
rect 6825 37275 6883 37281
rect 9309 37315 9367 37321
rect 9309 37281 9321 37315
rect 9355 37312 9367 37315
rect 10045 37315 10103 37321
rect 9355 37284 9720 37312
rect 9355 37281 9367 37284
rect 9309 37275 9367 37281
rect 9692 37256 9720 37284
rect 10045 37281 10057 37315
rect 10091 37312 10103 37315
rect 11514 37312 11520 37324
rect 10091 37284 11520 37312
rect 10091 37281 10103 37284
rect 10045 37275 10103 37281
rect 11514 37272 11520 37284
rect 11572 37272 11578 37324
rect 12894 37272 12900 37324
rect 12952 37312 12958 37324
rect 13725 37315 13783 37321
rect 13725 37312 13737 37315
rect 12952 37284 13737 37312
rect 12952 37272 12958 37284
rect 13725 37281 13737 37284
rect 13771 37312 13783 37315
rect 14277 37315 14335 37321
rect 14277 37312 14289 37315
rect 13771 37284 14289 37312
rect 13771 37281 13783 37284
rect 13725 37275 13783 37281
rect 14277 37281 14289 37284
rect 14323 37281 14335 37315
rect 14277 37275 14335 37281
rect 20809 37315 20867 37321
rect 20809 37281 20821 37315
rect 20855 37281 20867 37315
rect 20809 37275 20867 37281
rect 21453 37315 21511 37321
rect 21453 37281 21465 37315
rect 21499 37312 21511 37315
rect 21910 37312 21916 37324
rect 21499 37284 21916 37312
rect 21499 37281 21511 37284
rect 21453 37275 21511 37281
rect 1673 37247 1731 37253
rect 1673 37244 1685 37247
rect 1452 37216 1685 37244
rect 1452 37204 1458 37216
rect 1673 37213 1685 37216
rect 1719 37213 1731 37247
rect 1673 37207 1731 37213
rect 2498 37204 2504 37256
rect 2556 37244 2562 37256
rect 2685 37247 2743 37253
rect 2685 37244 2697 37247
rect 2556 37216 2697 37244
rect 2556 37204 2562 37216
rect 2685 37213 2697 37216
rect 2731 37213 2743 37247
rect 2685 37207 2743 37213
rect 4893 37247 4951 37253
rect 4893 37213 4905 37247
rect 4939 37244 4951 37247
rect 5997 37247 6055 37253
rect 4939 37216 5488 37244
rect 4939 37213 4951 37216
rect 4893 37207 4951 37213
rect 5460 37120 5488 37216
rect 5997 37213 6009 37247
rect 6043 37244 6055 37247
rect 6454 37244 6460 37256
rect 6043 37216 6460 37244
rect 6043 37213 6055 37216
rect 5997 37207 6055 37213
rect 6454 37204 6460 37216
rect 6512 37244 6518 37256
rect 6641 37247 6699 37253
rect 6641 37244 6653 37247
rect 6512 37216 6653 37244
rect 6512 37204 6518 37216
rect 6641 37213 6653 37216
rect 6687 37213 6699 37247
rect 8110 37244 8116 37256
rect 8071 37216 8116 37244
rect 6641 37207 6699 37213
rect 8110 37204 8116 37216
rect 8168 37204 8174 37256
rect 9674 37204 9680 37256
rect 9732 37244 9738 37256
rect 9861 37247 9919 37253
rect 9861 37244 9873 37247
rect 9732 37216 9873 37244
rect 9732 37204 9738 37216
rect 9861 37213 9873 37216
rect 9907 37213 9919 37247
rect 9861 37207 9919 37213
rect 13449 37247 13507 37253
rect 13449 37213 13461 37247
rect 13495 37213 13507 37247
rect 15194 37244 15200 37256
rect 15155 37216 15200 37244
rect 13449 37207 13507 37213
rect 10686 37136 10692 37188
rect 10744 37176 10750 37188
rect 13464 37176 13492 37207
rect 15194 37204 15200 37216
rect 15252 37204 15258 37256
rect 17126 37244 17132 37256
rect 17087 37216 17132 37244
rect 17126 37204 17132 37216
rect 17184 37204 17190 37256
rect 18414 37244 18420 37256
rect 18375 37216 18420 37244
rect 18414 37204 18420 37216
rect 18472 37204 18478 37256
rect 20346 37244 20352 37256
rect 20307 37216 20352 37244
rect 20346 37204 20352 37216
rect 20404 37244 20410 37256
rect 20824 37244 20852 37275
rect 21910 37272 21916 37284
rect 21968 37312 21974 37324
rect 22005 37315 22063 37321
rect 22005 37312 22017 37315
rect 21968 37284 22017 37312
rect 21968 37272 21974 37284
rect 22005 37281 22017 37284
rect 22051 37281 22063 37315
rect 22005 37275 22063 37281
rect 24765 37315 24823 37321
rect 24765 37281 24777 37315
rect 24811 37312 24823 37315
rect 24811 37284 25176 37312
rect 24811 37281 24823 37284
rect 24765 37275 24823 37281
rect 25148 37256 25176 37284
rect 22278 37244 22284 37256
rect 20404 37216 20852 37244
rect 22239 37216 22284 37244
rect 20404 37204 20410 37216
rect 22278 37204 22284 37216
rect 22336 37204 22342 37256
rect 23198 37204 23204 37256
rect 23256 37244 23262 37256
rect 23477 37247 23535 37253
rect 23477 37244 23489 37247
rect 23256 37216 23489 37244
rect 23256 37204 23262 37216
rect 23477 37213 23489 37216
rect 23523 37213 23535 37247
rect 23477 37207 23535 37213
rect 25130 37204 25136 37256
rect 25188 37244 25194 37256
rect 25317 37247 25375 37253
rect 25317 37244 25329 37247
rect 25188 37216 25329 37244
rect 25188 37204 25194 37216
rect 25317 37213 25329 37216
rect 25363 37213 25375 37247
rect 25317 37207 25375 37213
rect 26605 37247 26663 37253
rect 26605 37213 26617 37247
rect 26651 37244 26663 37247
rect 27154 37244 27160 37256
rect 26651 37216 27160 37244
rect 26651 37213 26663 37216
rect 26605 37207 26663 37213
rect 27154 37204 27160 37216
rect 27212 37204 27218 37256
rect 27338 37204 27344 37256
rect 27396 37244 27402 37256
rect 28445 37247 28503 37253
rect 28445 37244 28457 37247
rect 27396 37216 28457 37244
rect 27396 37204 27402 37216
rect 28445 37213 28457 37216
rect 28491 37213 28503 37247
rect 30374 37244 30380 37256
rect 30335 37216 30380 37244
rect 28445 37207 28503 37213
rect 30374 37204 30380 37216
rect 30432 37204 30438 37256
rect 30650 37204 30656 37256
rect 30708 37244 30714 37256
rect 32309 37247 32367 37253
rect 32309 37244 32321 37247
rect 30708 37216 32321 37244
rect 30708 37204 30714 37216
rect 32309 37213 32321 37216
rect 32355 37213 32367 37247
rect 33594 37244 33600 37256
rect 33555 37216 33600 37244
rect 32309 37207 32367 37213
rect 33594 37204 33600 37216
rect 33652 37204 33658 37256
rect 34790 37204 34796 37256
rect 34848 37244 34854 37256
rect 35529 37247 35587 37253
rect 35529 37244 35541 37247
rect 34848 37216 35541 37244
rect 34848 37204 34854 37216
rect 35529 37213 35541 37216
rect 35575 37213 35587 37247
rect 35529 37207 35587 37213
rect 36633 37247 36691 37253
rect 36633 37213 36645 37247
rect 36679 37213 36691 37247
rect 37461 37247 37519 37253
rect 37461 37244 37473 37247
rect 36633 37207 36691 37213
rect 36740 37216 37473 37244
rect 15562 37176 15568 37188
rect 10744 37148 15568 37176
rect 10744 37136 10750 37148
rect 15562 37136 15568 37148
rect 15620 37136 15626 37188
rect 26326 37136 26332 37188
rect 26384 37176 26390 37188
rect 36446 37176 36452 37188
rect 26384 37148 36452 37176
rect 26384 37136 26390 37148
rect 36446 37136 36452 37148
rect 36504 37176 36510 37188
rect 36648 37176 36676 37207
rect 36504 37148 36676 37176
rect 36504 37136 36510 37148
rect 1762 37108 1768 37120
rect 1723 37080 1768 37108
rect 1762 37068 1768 37080
rect 1820 37068 1826 37120
rect 2774 37068 2780 37120
rect 2832 37108 2838 37120
rect 2869 37111 2927 37117
rect 2869 37108 2881 37111
rect 2832 37080 2881 37108
rect 2832 37068 2838 37080
rect 2869 37077 2881 37080
rect 2915 37077 2927 37111
rect 2869 37071 2927 37077
rect 4614 37068 4620 37120
rect 4672 37108 4678 37120
rect 4709 37111 4767 37117
rect 4709 37108 4721 37111
rect 4672 37080 4721 37108
rect 4672 37068 4678 37080
rect 4709 37077 4721 37080
rect 4755 37077 4767 37111
rect 5442 37108 5448 37120
rect 5403 37080 5448 37108
rect 4709 37071 4767 37077
rect 5442 37068 5448 37080
rect 5500 37068 5506 37120
rect 7742 37068 7748 37120
rect 7800 37108 7806 37120
rect 7929 37111 7987 37117
rect 7929 37108 7941 37111
rect 7800 37080 7941 37108
rect 7800 37068 7806 37080
rect 7929 37077 7941 37080
rect 7975 37077 7987 37111
rect 7929 37071 7987 37077
rect 14826 37068 14832 37120
rect 14884 37108 14890 37120
rect 15013 37111 15071 37117
rect 15013 37108 15025 37111
rect 14884 37080 15025 37108
rect 14884 37068 14890 37080
rect 15013 37077 15025 37080
rect 15059 37077 15071 37111
rect 15013 37071 15071 37077
rect 16758 37068 16764 37120
rect 16816 37108 16822 37120
rect 16945 37111 17003 37117
rect 16945 37108 16957 37111
rect 16816 37080 16957 37108
rect 16816 37068 16822 37080
rect 16945 37077 16957 37080
rect 16991 37077 17003 37111
rect 16945 37071 17003 37077
rect 18046 37068 18052 37120
rect 18104 37108 18110 37120
rect 18233 37111 18291 37117
rect 18233 37108 18245 37111
rect 18104 37080 18245 37108
rect 18104 37068 18110 37080
rect 18233 37077 18245 37080
rect 18279 37077 18291 37111
rect 18233 37071 18291 37077
rect 19978 37068 19984 37120
rect 20036 37108 20042 37120
rect 20165 37111 20223 37117
rect 20165 37108 20177 37111
rect 20036 37080 20177 37108
rect 20036 37068 20042 37080
rect 20165 37077 20177 37080
rect 20211 37077 20223 37111
rect 25406 37108 25412 37120
rect 25367 37080 25412 37108
rect 20165 37071 20223 37077
rect 25406 37068 25412 37080
rect 25464 37068 25470 37120
rect 27062 37068 27068 37120
rect 27120 37108 27126 37120
rect 27341 37111 27399 37117
rect 27341 37108 27353 37111
rect 27120 37080 27353 37108
rect 27120 37068 27126 37080
rect 27341 37077 27353 37080
rect 27387 37077 27399 37111
rect 27341 37071 27399 37077
rect 28350 37068 28356 37120
rect 28408 37108 28414 37120
rect 28629 37111 28687 37117
rect 28629 37108 28641 37111
rect 28408 37080 28641 37108
rect 28408 37068 28414 37080
rect 28629 37077 28641 37080
rect 28675 37077 28687 37111
rect 28629 37071 28687 37077
rect 30282 37068 30288 37120
rect 30340 37108 30346 37120
rect 30561 37111 30619 37117
rect 30561 37108 30573 37111
rect 30340 37080 30573 37108
rect 30340 37068 30346 37080
rect 30561 37077 30573 37080
rect 30607 37077 30619 37111
rect 30561 37071 30619 37077
rect 32214 37068 32220 37120
rect 32272 37108 32278 37120
rect 32493 37111 32551 37117
rect 32493 37108 32505 37111
rect 32272 37080 32505 37108
rect 32272 37068 32278 37080
rect 32493 37077 32505 37080
rect 32539 37077 32551 37111
rect 32493 37071 32551 37077
rect 33502 37068 33508 37120
rect 33560 37108 33566 37120
rect 33781 37111 33839 37117
rect 33781 37108 33793 37111
rect 33560 37080 33793 37108
rect 33560 37068 33566 37080
rect 33781 37077 33793 37080
rect 33827 37077 33839 37111
rect 33781 37071 33839 37077
rect 34790 37068 34796 37120
rect 34848 37108 34854 37120
rect 34977 37111 35035 37117
rect 34977 37108 34989 37111
rect 34848 37080 34989 37108
rect 34848 37068 34854 37080
rect 34977 37077 34989 37080
rect 35023 37077 35035 37111
rect 34977 37071 35035 37077
rect 35434 37068 35440 37120
rect 35492 37108 35498 37120
rect 35713 37111 35771 37117
rect 35713 37108 35725 37111
rect 35492 37080 35725 37108
rect 35492 37068 35498 37080
rect 35713 37077 35725 37080
rect 35759 37077 35771 37111
rect 35713 37071 35771 37077
rect 36262 37068 36268 37120
rect 36320 37108 36326 37120
rect 36740 37108 36768 37216
rect 37461 37213 37473 37216
rect 37507 37213 37519 37247
rect 37461 37207 37519 37213
rect 36320 37080 36768 37108
rect 36320 37068 36326 37080
rect 37366 37068 37372 37120
rect 37424 37108 37430 37120
rect 37645 37111 37703 37117
rect 37645 37108 37657 37111
rect 37424 37080 37657 37108
rect 37424 37068 37430 37080
rect 37645 37077 37657 37080
rect 37691 37077 37703 37111
rect 37645 37071 37703 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 2409 36907 2467 36913
rect 2409 36873 2421 36907
rect 2455 36904 2467 36907
rect 2866 36904 2872 36916
rect 2455 36876 2872 36904
rect 2455 36873 2467 36876
rect 2409 36867 2467 36873
rect 2866 36864 2872 36876
rect 2924 36864 2930 36916
rect 6549 36907 6607 36913
rect 6549 36873 6561 36907
rect 6595 36873 6607 36907
rect 6549 36867 6607 36873
rect 1670 36836 1676 36848
rect 1631 36808 1676 36836
rect 1670 36796 1676 36808
rect 1728 36836 1734 36848
rect 3053 36839 3111 36845
rect 3053 36836 3065 36839
rect 1728 36808 3065 36836
rect 1728 36796 1734 36808
rect 3053 36805 3065 36808
rect 3099 36805 3111 36839
rect 3053 36799 3111 36805
rect 2593 36771 2651 36777
rect 2593 36737 2605 36771
rect 2639 36768 2651 36771
rect 6564 36768 6592 36867
rect 8110 36864 8116 36916
rect 8168 36904 8174 36916
rect 10505 36907 10563 36913
rect 10505 36904 10517 36907
rect 8168 36876 10517 36904
rect 8168 36864 8174 36876
rect 10505 36873 10517 36876
rect 10551 36873 10563 36907
rect 23198 36904 23204 36916
rect 23159 36876 23204 36904
rect 10505 36867 10563 36873
rect 23198 36864 23204 36876
rect 23256 36864 23262 36916
rect 27341 36907 27399 36913
rect 27341 36873 27353 36907
rect 27387 36904 27399 36907
rect 33594 36904 33600 36916
rect 27387 36876 33600 36904
rect 27387 36873 27399 36876
rect 27341 36867 27399 36873
rect 33594 36864 33600 36876
rect 33652 36864 33658 36916
rect 34977 36907 35035 36913
rect 34977 36873 34989 36907
rect 35023 36904 35035 36907
rect 36262 36904 36268 36916
rect 35023 36876 36268 36904
rect 35023 36873 35035 36876
rect 34977 36867 35035 36873
rect 36262 36864 36268 36876
rect 36320 36864 36326 36916
rect 36446 36904 36452 36916
rect 36407 36876 36452 36904
rect 36446 36864 36452 36876
rect 36504 36864 36510 36916
rect 38194 36904 38200 36916
rect 38155 36876 38200 36904
rect 38194 36864 38200 36876
rect 38252 36864 38258 36916
rect 2639 36740 6592 36768
rect 6733 36771 6791 36777
rect 2639 36737 2651 36740
rect 2593 36731 2651 36737
rect 6733 36737 6745 36771
rect 6779 36768 6791 36771
rect 10686 36768 10692 36780
rect 6779 36740 6914 36768
rect 10647 36740 10692 36768
rect 6779 36737 6791 36740
rect 6733 36731 6791 36737
rect 6886 36700 6914 36740
rect 10686 36728 10692 36740
rect 10744 36728 10750 36780
rect 11606 36728 11612 36780
rect 11664 36768 11670 36780
rect 11701 36771 11759 36777
rect 11701 36768 11713 36771
rect 11664 36740 11713 36768
rect 11664 36728 11670 36740
rect 11701 36737 11713 36740
rect 11747 36737 11759 36771
rect 11701 36731 11759 36737
rect 22278 36728 22284 36780
rect 22336 36768 22342 36780
rect 27157 36771 27215 36777
rect 27157 36768 27169 36771
rect 22336 36740 27169 36768
rect 22336 36728 22342 36740
rect 27157 36737 27169 36740
rect 27203 36737 27215 36771
rect 27157 36731 27215 36737
rect 34885 36771 34943 36777
rect 34885 36737 34897 36771
rect 34931 36768 34943 36771
rect 35526 36768 35532 36780
rect 34931 36740 35532 36768
rect 34931 36737 34943 36740
rect 34885 36731 34943 36737
rect 35526 36728 35532 36740
rect 35584 36728 35590 36780
rect 37274 36728 37280 36780
rect 37332 36768 37338 36780
rect 38013 36771 38071 36777
rect 38013 36768 38025 36771
rect 37332 36740 38025 36768
rect 37332 36728 37338 36740
rect 38013 36737 38025 36740
rect 38059 36737 38071 36771
rect 38013 36731 38071 36737
rect 11974 36700 11980 36712
rect 6886 36672 11980 36700
rect 11974 36660 11980 36672
rect 12032 36660 12038 36712
rect 1857 36635 1915 36641
rect 1857 36601 1869 36635
rect 1903 36632 1915 36635
rect 2130 36632 2136 36644
rect 1903 36604 2136 36632
rect 1903 36601 1915 36604
rect 1857 36595 1915 36601
rect 2130 36592 2136 36604
rect 2188 36592 2194 36644
rect 35526 36564 35532 36576
rect 35487 36536 35532 36564
rect 35526 36524 35532 36536
rect 35584 36524 35590 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 11606 36360 11612 36372
rect 11567 36332 11612 36360
rect 11606 36320 11612 36332
rect 11664 36320 11670 36372
rect 38197 36363 38255 36369
rect 38197 36329 38209 36363
rect 38243 36360 38255 36363
rect 38654 36360 38660 36372
rect 38243 36332 38660 36360
rect 38243 36329 38255 36332
rect 38197 36323 38255 36329
rect 38654 36320 38660 36332
rect 38712 36320 38718 36372
rect 37553 36295 37611 36301
rect 37553 36261 37565 36295
rect 37599 36261 37611 36295
rect 37553 36255 37611 36261
rect 1854 36156 1860 36168
rect 1815 36128 1860 36156
rect 1854 36116 1860 36128
rect 1912 36116 1918 36168
rect 37366 36156 37372 36168
rect 37327 36128 37372 36156
rect 37366 36116 37372 36128
rect 37424 36116 37430 36168
rect 37568 36156 37596 36255
rect 38013 36159 38071 36165
rect 38013 36156 38025 36159
rect 37568 36128 38025 36156
rect 38013 36125 38025 36128
rect 38059 36125 38071 36159
rect 38013 36119 38071 36125
rect 1670 36020 1676 36032
rect 1631 35992 1676 36020
rect 1670 35980 1676 35992
rect 1728 35980 1734 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 29549 35819 29607 35825
rect 29549 35785 29561 35819
rect 29595 35816 29607 35819
rect 30374 35816 30380 35828
rect 29595 35788 30380 35816
rect 29595 35785 29607 35788
rect 29549 35779 29607 35785
rect 30374 35776 30380 35788
rect 30432 35776 30438 35828
rect 28534 35640 28540 35692
rect 28592 35680 28598 35692
rect 29365 35683 29423 35689
rect 29365 35680 29377 35683
rect 28592 35652 29377 35680
rect 28592 35640 28598 35652
rect 29365 35649 29377 35652
rect 29411 35649 29423 35683
rect 29365 35643 29423 35649
rect 37366 35572 37372 35624
rect 37424 35612 37430 35624
rect 38013 35615 38071 35621
rect 38013 35612 38025 35615
rect 37424 35584 38025 35612
rect 37424 35572 37430 35584
rect 38013 35581 38025 35584
rect 38059 35581 38071 35615
rect 38286 35612 38292 35624
rect 38247 35584 38292 35612
rect 38013 35575 38071 35581
rect 38286 35572 38292 35584
rect 38344 35572 38350 35624
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 38286 35272 38292 35284
rect 38247 35244 38292 35272
rect 38286 35232 38292 35244
rect 38344 35232 38350 35284
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1854 34688 1860 34740
rect 1912 34728 1918 34740
rect 2409 34731 2467 34737
rect 2409 34728 2421 34731
rect 1912 34700 2421 34728
rect 1912 34688 1918 34700
rect 2409 34697 2421 34700
rect 2455 34697 2467 34731
rect 2409 34691 2467 34697
rect 1857 34595 1915 34601
rect 1857 34561 1869 34595
rect 1903 34592 1915 34595
rect 2038 34592 2044 34604
rect 1903 34564 2044 34592
rect 1903 34561 1915 34564
rect 1857 34555 1915 34561
rect 2038 34552 2044 34564
rect 2096 34552 2102 34604
rect 2501 34595 2559 34601
rect 2501 34561 2513 34595
rect 2547 34592 2559 34595
rect 2547 34564 3096 34592
rect 2547 34561 2559 34564
rect 2501 34555 2559 34561
rect 3068 34533 3096 34564
rect 3053 34527 3111 34533
rect 3053 34493 3065 34527
rect 3099 34524 3111 34527
rect 13078 34524 13084 34536
rect 3099 34496 13084 34524
rect 3099 34493 3111 34496
rect 3053 34487 3111 34493
rect 13078 34484 13084 34496
rect 13136 34484 13142 34536
rect 1670 34388 1676 34400
rect 1631 34360 1676 34388
rect 1670 34348 1676 34360
rect 1728 34348 1734 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 25682 33464 25688 33516
rect 25740 33504 25746 33516
rect 37461 33507 37519 33513
rect 37461 33504 37473 33507
rect 25740 33476 37473 33504
rect 25740 33464 25746 33476
rect 37461 33473 37473 33476
rect 37507 33504 37519 33507
rect 38013 33507 38071 33513
rect 38013 33504 38025 33507
rect 37507 33476 38025 33504
rect 37507 33473 37519 33476
rect 37461 33467 37519 33473
rect 38013 33473 38025 33476
rect 38059 33473 38071 33507
rect 38013 33467 38071 33473
rect 38194 33368 38200 33380
rect 38155 33340 38200 33368
rect 38194 33328 38200 33340
rect 38252 33328 38258 33380
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 27338 32552 27344 32564
rect 27299 32524 27344 32552
rect 27338 32512 27344 32524
rect 27396 32512 27402 32564
rect 1857 32419 1915 32425
rect 1857 32385 1869 32419
rect 1903 32416 1915 32419
rect 9122 32416 9128 32428
rect 1903 32388 9128 32416
rect 1903 32385 1915 32388
rect 1857 32379 1915 32385
rect 9122 32376 9128 32388
rect 9180 32376 9186 32428
rect 27157 32419 27215 32425
rect 27157 32385 27169 32419
rect 27203 32416 27215 32419
rect 27203 32388 27936 32416
rect 27203 32385 27215 32388
rect 27157 32379 27215 32385
rect 1670 32212 1676 32224
rect 1631 32184 1676 32212
rect 1670 32172 1676 32184
rect 1728 32172 1734 32224
rect 27908 32221 27936 32388
rect 28534 32308 28540 32360
rect 28592 32348 28598 32360
rect 38013 32351 38071 32357
rect 38013 32348 38025 32351
rect 28592 32320 38025 32348
rect 28592 32308 28598 32320
rect 38013 32317 38025 32320
rect 38059 32317 38071 32351
rect 38286 32348 38292 32360
rect 38247 32320 38292 32348
rect 38013 32311 38071 32317
rect 38286 32308 38292 32320
rect 38344 32308 38350 32360
rect 27893 32215 27951 32221
rect 27893 32181 27905 32215
rect 27939 32212 27951 32215
rect 28626 32212 28632 32224
rect 27939 32184 28632 32212
rect 27939 32181 27951 32184
rect 27893 32175 27951 32181
rect 28626 32172 28632 32184
rect 28684 32172 28690 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 38286 32008 38292 32020
rect 38247 31980 38292 32008
rect 38286 31968 38292 31980
rect 38344 31968 38350 32020
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 2498 30920 2504 30932
rect 2459 30892 2504 30920
rect 2498 30880 2504 30892
rect 2556 30880 2562 30932
rect 27341 30923 27399 30929
rect 27341 30889 27353 30923
rect 27387 30920 27399 30923
rect 30650 30920 30656 30932
rect 27387 30892 30656 30920
rect 27387 30889 27399 30892
rect 27341 30883 27399 30889
rect 30650 30880 30656 30892
rect 30708 30880 30714 30932
rect 1946 30676 1952 30728
rect 2004 30716 2010 30728
rect 2317 30719 2375 30725
rect 2317 30716 2329 30719
rect 2004 30688 2329 30716
rect 2004 30676 2010 30688
rect 2317 30685 2329 30688
rect 2363 30716 2375 30719
rect 2961 30719 3019 30725
rect 2961 30716 2973 30719
rect 2363 30688 2973 30716
rect 2363 30685 2375 30688
rect 2317 30679 2375 30685
rect 2961 30685 2973 30688
rect 3007 30685 3019 30719
rect 2961 30679 3019 30685
rect 26970 30676 26976 30728
rect 27028 30716 27034 30728
rect 27157 30719 27215 30725
rect 27157 30716 27169 30719
rect 27028 30688 27169 30716
rect 27028 30676 27034 30688
rect 27157 30685 27169 30688
rect 27203 30716 27215 30719
rect 27801 30719 27859 30725
rect 27801 30716 27813 30719
rect 27203 30688 27813 30716
rect 27203 30685 27215 30688
rect 27157 30679 27215 30685
rect 27801 30685 27813 30688
rect 27847 30685 27859 30719
rect 27801 30679 27859 30685
rect 1670 30648 1676 30660
rect 1631 30620 1676 30648
rect 1670 30608 1676 30620
rect 1728 30608 1734 30660
rect 1857 30651 1915 30657
rect 1857 30617 1869 30651
rect 1903 30648 1915 30651
rect 2222 30648 2228 30660
rect 1903 30620 2228 30648
rect 1903 30617 1915 30620
rect 1857 30611 1915 30617
rect 2222 30608 2228 30620
rect 2280 30608 2286 30660
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 1670 30376 1676 30388
rect 1631 30348 1676 30376
rect 1670 30336 1676 30348
rect 1728 30336 1734 30388
rect 30190 30240 30196 30252
rect 30151 30212 30196 30240
rect 30190 30200 30196 30212
rect 30248 30240 30254 30252
rect 30837 30243 30895 30249
rect 30837 30240 30849 30243
rect 30248 30212 30849 30240
rect 30248 30200 30254 30212
rect 30837 30209 30849 30212
rect 30883 30209 30895 30243
rect 30837 30203 30895 30209
rect 37553 30243 37611 30249
rect 37553 30209 37565 30243
rect 37599 30240 37611 30243
rect 38194 30240 38200 30252
rect 37599 30212 38200 30240
rect 37599 30209 37611 30212
rect 37553 30203 37611 30209
rect 38194 30200 38200 30212
rect 38252 30200 38258 30252
rect 30377 30107 30435 30113
rect 30377 30073 30389 30107
rect 30423 30104 30435 30107
rect 37274 30104 37280 30116
rect 30423 30076 37280 30104
rect 30423 30073 30435 30076
rect 30377 30067 30435 30073
rect 37274 30064 37280 30076
rect 37332 30064 37338 30116
rect 38102 30036 38108 30048
rect 38063 30008 38108 30036
rect 38102 29996 38108 30008
rect 38160 29996 38166 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 23109 29563 23167 29569
rect 23109 29529 23121 29563
rect 23155 29529 23167 29563
rect 23109 29523 23167 29529
rect 5442 29452 5448 29504
rect 5500 29492 5506 29504
rect 23017 29495 23075 29501
rect 23017 29492 23029 29495
rect 5500 29464 23029 29492
rect 5500 29452 5506 29464
rect 23017 29461 23029 29464
rect 23063 29461 23075 29495
rect 23124 29492 23152 29523
rect 23658 29492 23664 29504
rect 23124 29464 23664 29492
rect 23017 29455 23075 29461
rect 23658 29452 23664 29464
rect 23716 29452 23722 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 1578 29112 1584 29164
rect 1636 29152 1642 29164
rect 1673 29155 1731 29161
rect 1673 29152 1685 29155
rect 1636 29124 1685 29152
rect 1636 29112 1642 29124
rect 1673 29121 1685 29124
rect 1719 29121 1731 29155
rect 1673 29115 1731 29121
rect 1857 29019 1915 29025
rect 1857 28985 1869 29019
rect 1903 29016 1915 29019
rect 25590 29016 25596 29028
rect 1903 28988 25596 29016
rect 1903 28985 1915 28988
rect 1857 28979 1915 28985
rect 25590 28976 25596 28988
rect 25648 28976 25654 29028
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 18414 28704 18420 28756
rect 18472 28744 18478 28756
rect 19981 28747 20039 28753
rect 19981 28744 19993 28747
rect 18472 28716 19993 28744
rect 18472 28704 18478 28716
rect 19981 28713 19993 28716
rect 20027 28713 20039 28747
rect 19981 28707 20039 28713
rect 1578 28676 1584 28688
rect 1539 28648 1584 28676
rect 1578 28636 1584 28648
rect 1636 28636 1642 28688
rect 15562 28540 15568 28552
rect 15523 28512 15568 28540
rect 15562 28500 15568 28512
rect 15620 28500 15626 28552
rect 20073 28543 20131 28549
rect 20073 28509 20085 28543
rect 20119 28540 20131 28543
rect 20119 28512 20668 28540
rect 20119 28509 20131 28512
rect 20073 28503 20131 28509
rect 15654 28404 15660 28416
rect 15615 28376 15660 28404
rect 15654 28364 15660 28376
rect 15712 28364 15718 28416
rect 20640 28413 20668 28512
rect 20625 28407 20683 28413
rect 20625 28373 20637 28407
rect 20671 28404 20683 28407
rect 23106 28404 23112 28416
rect 20671 28376 23112 28404
rect 20671 28373 20683 28376
rect 20625 28367 20683 28373
rect 23106 28364 23112 28376
rect 23164 28364 23170 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 17126 28160 17132 28212
rect 17184 28200 17190 28212
rect 19245 28203 19303 28209
rect 19245 28200 19257 28203
rect 17184 28172 19257 28200
rect 17184 28160 17190 28172
rect 19245 28169 19257 28172
rect 19291 28169 19303 28203
rect 25590 28200 25596 28212
rect 25551 28172 25596 28200
rect 19245 28163 19303 28169
rect 25590 28160 25596 28172
rect 25648 28160 25654 28212
rect 26326 28200 26332 28212
rect 26287 28172 26332 28200
rect 26326 28160 26332 28172
rect 26384 28160 26390 28212
rect 15194 28092 15200 28144
rect 15252 28132 15258 28144
rect 18417 28135 18475 28141
rect 18417 28132 18429 28135
rect 15252 28104 18429 28132
rect 15252 28092 15258 28104
rect 18417 28101 18429 28104
rect 18463 28101 18475 28135
rect 18417 28095 18475 28101
rect 18506 28064 18512 28076
rect 18467 28036 18512 28064
rect 18506 28024 18512 28036
rect 18564 28024 18570 28076
rect 19337 28067 19395 28073
rect 19337 28033 19349 28067
rect 19383 28033 19395 28067
rect 19337 28027 19395 28033
rect 22189 28067 22247 28073
rect 22189 28033 22201 28067
rect 22235 28064 22247 28067
rect 22278 28064 22284 28076
rect 22235 28036 22284 28064
rect 22235 28033 22247 28036
rect 22189 28027 22247 28033
rect 19352 27996 19380 28027
rect 22278 28024 22284 28036
rect 22336 28024 22342 28076
rect 25608 28064 25636 28160
rect 26145 28067 26203 28073
rect 26145 28064 26157 28067
rect 25608 28036 26157 28064
rect 26145 28033 26157 28036
rect 26191 28033 26203 28067
rect 28534 28064 28540 28076
rect 28495 28036 28540 28064
rect 26145 28027 26203 28033
rect 28534 28024 28540 28036
rect 28592 28024 28598 28076
rect 37553 28067 37611 28073
rect 37553 28033 37565 28067
rect 37599 28064 37611 28067
rect 38194 28064 38200 28076
rect 37599 28036 38200 28064
rect 37599 28033 37611 28036
rect 37553 28027 37611 28033
rect 38194 28024 38200 28036
rect 38252 28024 38258 28076
rect 24762 27996 24768 28008
rect 19352 27968 24768 27996
rect 24762 27956 24768 27968
rect 24820 27956 24826 28008
rect 24854 27888 24860 27940
rect 24912 27928 24918 27940
rect 28445 27931 28503 27937
rect 28445 27928 28457 27931
rect 24912 27900 28457 27928
rect 24912 27888 24918 27900
rect 28445 27897 28457 27900
rect 28491 27897 28503 27931
rect 28445 27891 28503 27897
rect 37918 27888 37924 27940
rect 37976 27928 37982 27940
rect 38013 27931 38071 27937
rect 38013 27928 38025 27931
rect 37976 27900 38025 27928
rect 37976 27888 37982 27900
rect 38013 27897 38025 27900
rect 38059 27897 38071 27931
rect 38013 27891 38071 27897
rect 22097 27863 22155 27869
rect 22097 27829 22109 27863
rect 22143 27860 22155 27863
rect 22922 27860 22928 27872
rect 22143 27832 22928 27860
rect 22143 27829 22155 27832
rect 22097 27823 22155 27829
rect 22922 27820 22928 27832
rect 22980 27820 22986 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 11974 27412 11980 27464
rect 12032 27452 12038 27464
rect 14829 27455 14887 27461
rect 14829 27452 14841 27455
rect 12032 27424 14841 27452
rect 12032 27412 12038 27424
rect 14829 27421 14841 27424
rect 14875 27421 14887 27455
rect 14829 27415 14887 27421
rect 32401 27455 32459 27461
rect 32401 27421 32413 27455
rect 32447 27452 32459 27455
rect 37366 27452 37372 27464
rect 32447 27424 37372 27452
rect 32447 27421 32459 27424
rect 32401 27415 32459 27421
rect 37366 27412 37372 27424
rect 37424 27412 37430 27464
rect 14921 27319 14979 27325
rect 14921 27285 14933 27319
rect 14967 27316 14979 27319
rect 15562 27316 15568 27328
rect 14967 27288 15568 27316
rect 14967 27285 14979 27288
rect 14921 27279 14979 27285
rect 15562 27276 15568 27288
rect 15620 27276 15626 27328
rect 18506 27276 18512 27328
rect 18564 27316 18570 27328
rect 18693 27319 18751 27325
rect 18693 27316 18705 27319
rect 18564 27288 18705 27316
rect 18564 27276 18570 27288
rect 18693 27285 18705 27288
rect 18739 27316 18751 27319
rect 21450 27316 21456 27328
rect 18739 27288 21456 27316
rect 18739 27285 18751 27288
rect 18693 27279 18751 27285
rect 21450 27276 21456 27288
rect 21508 27276 21514 27328
rect 26418 27276 26424 27328
rect 26476 27316 26482 27328
rect 32309 27319 32367 27325
rect 32309 27316 32321 27319
rect 26476 27288 32321 27316
rect 26476 27276 26482 27288
rect 32309 27285 32321 27288
rect 32355 27285 32367 27319
rect 32309 27279 32367 27285
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 1857 26979 1915 26985
rect 1857 26945 1869 26979
rect 1903 26976 1915 26979
rect 6822 26976 6828 26988
rect 1903 26948 6828 26976
rect 1903 26945 1915 26948
rect 1857 26939 1915 26945
rect 6822 26936 6828 26948
rect 6880 26936 6886 26988
rect 23658 26868 23664 26920
rect 23716 26908 23722 26920
rect 38013 26911 38071 26917
rect 38013 26908 38025 26911
rect 23716 26880 38025 26908
rect 23716 26868 23722 26880
rect 38013 26877 38025 26880
rect 38059 26877 38071 26911
rect 38286 26908 38292 26920
rect 38247 26880 38292 26908
rect 38013 26871 38071 26877
rect 38286 26868 38292 26880
rect 38344 26868 38350 26920
rect 1670 26772 1676 26784
rect 1631 26744 1676 26772
rect 1670 26732 1676 26744
rect 1728 26732 1734 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 38286 26568 38292 26580
rect 38247 26540 38292 26568
rect 38286 26528 38292 26540
rect 38344 26528 38350 26580
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 2038 25440 2044 25492
rect 2096 25480 2102 25492
rect 7193 25483 7251 25489
rect 7193 25480 7205 25483
rect 2096 25452 7205 25480
rect 2096 25440 2102 25452
rect 7193 25449 7205 25452
rect 7239 25449 7251 25483
rect 9122 25480 9128 25492
rect 9083 25452 9128 25480
rect 7193 25443 7251 25449
rect 9122 25440 9128 25452
rect 9180 25440 9186 25492
rect 1578 25276 1584 25288
rect 1539 25248 1584 25276
rect 1578 25236 1584 25248
rect 1636 25236 1642 25288
rect 1857 25279 1915 25285
rect 1857 25245 1869 25279
rect 1903 25276 1915 25279
rect 1946 25276 1952 25288
rect 1903 25248 1952 25276
rect 1903 25245 1915 25248
rect 1857 25239 1915 25245
rect 1946 25236 1952 25248
rect 2004 25236 2010 25288
rect 7377 25279 7435 25285
rect 7377 25245 7389 25279
rect 7423 25276 7435 25279
rect 9309 25279 9367 25285
rect 7423 25248 7880 25276
rect 7423 25245 7435 25248
rect 7377 25239 7435 25245
rect 7852 25152 7880 25248
rect 9309 25245 9321 25279
rect 9355 25276 9367 25279
rect 9355 25248 9812 25276
rect 9355 25245 9367 25248
rect 9309 25239 9367 25245
rect 9784 25152 9812 25248
rect 7834 25140 7840 25152
rect 7795 25112 7840 25140
rect 7834 25100 7840 25112
rect 7892 25100 7898 25152
rect 9766 25140 9772 25152
rect 9727 25112 9772 25140
rect 9766 25100 9772 25112
rect 9824 25100 9830 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 1578 24936 1584 24948
rect 1539 24908 1584 24936
rect 1578 24896 1584 24908
rect 1636 24896 1642 24948
rect 37826 24692 37832 24744
rect 37884 24732 37890 24744
rect 38013 24735 38071 24741
rect 38013 24732 38025 24735
rect 37884 24704 38025 24732
rect 37884 24692 37890 24704
rect 38013 24701 38025 24704
rect 38059 24701 38071 24735
rect 38286 24732 38292 24744
rect 38247 24704 38292 24732
rect 38013 24695 38071 24701
rect 38286 24692 38292 24704
rect 38344 24692 38350 24744
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 38286 24392 38292 24404
rect 38247 24364 38292 24392
rect 38286 24352 38292 24364
rect 38344 24352 38350 24404
rect 20346 24148 20352 24200
rect 20404 24188 20410 24200
rect 27798 24188 27804 24200
rect 20404 24160 27804 24188
rect 20404 24148 20410 24160
rect 27798 24148 27804 24160
rect 27856 24148 27862 24200
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 1578 23644 1584 23656
rect 1539 23616 1584 23644
rect 1578 23604 1584 23616
rect 1636 23604 1642 23656
rect 1854 23644 1860 23656
rect 1815 23616 1860 23644
rect 1854 23604 1860 23616
rect 1912 23604 1918 23656
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 23658 23264 23664 23316
rect 23716 23304 23722 23316
rect 23845 23307 23903 23313
rect 23845 23304 23857 23307
rect 23716 23276 23857 23304
rect 23716 23264 23722 23276
rect 23845 23273 23857 23276
rect 23891 23273 23903 23307
rect 23845 23267 23903 23273
rect 1578 23236 1584 23248
rect 1539 23208 1584 23236
rect 1578 23196 1584 23208
rect 1636 23196 1642 23248
rect 23385 23103 23443 23109
rect 23385 23069 23397 23103
rect 23431 23100 23443 23103
rect 23658 23100 23664 23112
rect 23431 23072 23664 23100
rect 23431 23069 23443 23072
rect 23385 23063 23443 23069
rect 23658 23060 23664 23072
rect 23716 23060 23722 23112
rect 22830 22924 22836 22976
rect 22888 22964 22894 22976
rect 23293 22967 23351 22973
rect 23293 22964 23305 22967
rect 22888 22936 23305 22964
rect 22888 22924 22894 22936
rect 23293 22933 23305 22936
rect 23339 22933 23351 22967
rect 23293 22927 23351 22933
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 35986 22584 35992 22636
rect 36044 22624 36050 22636
rect 38013 22627 38071 22633
rect 38013 22624 38025 22627
rect 36044 22596 38025 22624
rect 36044 22584 36050 22596
rect 38013 22593 38025 22596
rect 38059 22593 38071 22627
rect 38013 22587 38071 22593
rect 38194 22488 38200 22500
rect 38155 22460 38200 22488
rect 38194 22448 38200 22460
rect 38252 22448 38258 22500
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 23569 22083 23627 22089
rect 23569 22049 23581 22083
rect 23615 22080 23627 22083
rect 25590 22080 25596 22092
rect 23615 22052 25596 22080
rect 23615 22049 23627 22052
rect 23569 22043 23627 22049
rect 23017 22015 23075 22021
rect 23017 21981 23029 22015
rect 23063 22012 23075 22015
rect 23584 22012 23612 22043
rect 25590 22040 25596 22052
rect 25648 22040 25654 22092
rect 23063 21984 23612 22012
rect 23063 21981 23075 21984
rect 23017 21975 23075 21981
rect 22646 21836 22652 21888
rect 22704 21876 22710 21888
rect 22925 21879 22983 21885
rect 22925 21876 22937 21879
rect 22704 21848 22937 21876
rect 22704 21836 22710 21848
rect 22925 21845 22937 21848
rect 22971 21845 22983 21879
rect 22925 21839 22983 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 6822 21632 6828 21684
rect 6880 21672 6886 21684
rect 6917 21675 6975 21681
rect 6917 21672 6929 21675
rect 6880 21644 6929 21672
rect 6880 21632 6886 21644
rect 6917 21641 6929 21644
rect 6963 21641 6975 21675
rect 25682 21672 25688 21684
rect 25643 21644 25688 21672
rect 6917 21635 6975 21641
rect 25682 21632 25688 21644
rect 25740 21632 25746 21684
rect 32769 21675 32827 21681
rect 32769 21641 32781 21675
rect 32815 21672 32827 21675
rect 35986 21672 35992 21684
rect 32815 21644 35992 21672
rect 32815 21641 32827 21644
rect 32769 21635 32827 21641
rect 35986 21632 35992 21644
rect 36044 21632 36050 21684
rect 1762 21496 1768 21548
rect 1820 21536 1826 21548
rect 1857 21539 1915 21545
rect 1857 21536 1869 21539
rect 1820 21508 1869 21536
rect 1820 21496 1826 21508
rect 1857 21505 1869 21508
rect 1903 21505 1915 21539
rect 1857 21499 1915 21505
rect 7101 21539 7159 21545
rect 7101 21505 7113 21539
rect 7147 21536 7159 21539
rect 25593 21539 25651 21545
rect 25593 21536 25605 21539
rect 7147 21508 7696 21536
rect 7147 21505 7159 21508
rect 7101 21499 7159 21505
rect 1670 21332 1676 21344
rect 1631 21304 1676 21332
rect 1670 21292 1676 21304
rect 1728 21292 1734 21344
rect 7668 21341 7696 21508
rect 24964 21508 25605 21536
rect 7653 21335 7711 21341
rect 7653 21301 7665 21335
rect 7699 21332 7711 21335
rect 13538 21332 13544 21344
rect 7699 21304 13544 21332
rect 7699 21301 7711 21304
rect 7653 21295 7711 21301
rect 13538 21292 13544 21304
rect 13596 21292 13602 21344
rect 21266 21292 21272 21344
rect 21324 21332 21330 21344
rect 24964 21341 24992 21508
rect 25593 21505 25605 21508
rect 25639 21505 25651 21539
rect 25593 21499 25651 21505
rect 30006 21496 30012 21548
rect 30064 21536 30070 21548
rect 32585 21539 32643 21545
rect 32585 21536 32597 21539
rect 30064 21508 32597 21536
rect 30064 21496 30070 21508
rect 32585 21505 32597 21508
rect 32631 21536 32643 21539
rect 33229 21539 33287 21545
rect 33229 21536 33241 21539
rect 32631 21508 33241 21536
rect 32631 21505 32643 21508
rect 32585 21499 32643 21505
rect 33229 21505 33241 21508
rect 33275 21505 33287 21539
rect 38010 21536 38016 21548
rect 37971 21508 38016 21536
rect 33229 21499 33287 21505
rect 38010 21496 38016 21508
rect 38068 21496 38074 21548
rect 24949 21335 25007 21341
rect 24949 21332 24961 21335
rect 21324 21304 24961 21332
rect 21324 21292 21330 21304
rect 24949 21301 24961 21304
rect 24995 21301 25007 21335
rect 38194 21332 38200 21344
rect 38155 21304 38200 21332
rect 24949 21295 25007 21301
rect 38194 21292 38200 21304
rect 38252 21292 38258 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 1762 21128 1768 21140
rect 1723 21100 1768 21128
rect 1762 21088 1768 21100
rect 1820 21088 1826 21140
rect 1946 20924 1952 20936
rect 1907 20896 1952 20924
rect 1946 20884 1952 20896
rect 2004 20884 2010 20936
rect 24765 20927 24823 20933
rect 24765 20893 24777 20927
rect 24811 20924 24823 20927
rect 24946 20924 24952 20936
rect 24811 20896 24952 20924
rect 24811 20893 24823 20896
rect 24765 20887 24823 20893
rect 24946 20884 24952 20896
rect 25004 20884 25010 20936
rect 13078 20748 13084 20800
rect 13136 20788 13142 20800
rect 20346 20788 20352 20800
rect 13136 20760 20352 20788
rect 13136 20748 13142 20760
rect 20346 20748 20352 20760
rect 20404 20748 20410 20800
rect 22002 20748 22008 20800
rect 22060 20788 22066 20800
rect 22097 20791 22155 20797
rect 22097 20788 22109 20791
rect 22060 20760 22109 20788
rect 22060 20748 22066 20760
rect 22097 20757 22109 20760
rect 22143 20757 22155 20791
rect 22097 20751 22155 20757
rect 24673 20791 24731 20797
rect 24673 20757 24685 20791
rect 24719 20788 24731 20791
rect 25130 20788 25136 20800
rect 24719 20760 25136 20788
rect 24719 20757 24731 20760
rect 24673 20751 24731 20757
rect 25130 20748 25136 20760
rect 25188 20748 25194 20800
rect 25406 20748 25412 20800
rect 25464 20788 25470 20800
rect 27522 20788 27528 20800
rect 25464 20760 27528 20788
rect 25464 20748 25470 20760
rect 27522 20748 27528 20760
rect 27580 20788 27586 20800
rect 30006 20788 30012 20800
rect 27580 20760 30012 20788
rect 27580 20748 27586 20760
rect 30006 20748 30012 20760
rect 30064 20748 30070 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 2222 20408 2228 20460
rect 2280 20448 2286 20460
rect 2280 20420 6914 20448
rect 2280 20408 2286 20420
rect 6886 20380 6914 20420
rect 22002 20408 22008 20460
rect 22060 20448 22066 20460
rect 22281 20451 22339 20457
rect 22281 20448 22293 20451
rect 22060 20420 22293 20448
rect 22060 20408 22066 20420
rect 22281 20417 22293 20420
rect 22327 20417 22339 20451
rect 22281 20411 22339 20417
rect 22925 20451 22983 20457
rect 22925 20417 22937 20451
rect 22971 20417 22983 20451
rect 22925 20411 22983 20417
rect 22940 20380 22968 20411
rect 23106 20408 23112 20460
rect 23164 20448 23170 20460
rect 24121 20451 24179 20457
rect 24121 20448 24133 20451
rect 23164 20420 24133 20448
rect 23164 20408 23170 20420
rect 24121 20417 24133 20420
rect 24167 20417 24179 20451
rect 24121 20411 24179 20417
rect 24765 20451 24823 20457
rect 24765 20417 24777 20451
rect 24811 20448 24823 20451
rect 24854 20448 24860 20460
rect 24811 20420 24860 20448
rect 24811 20417 24823 20420
rect 24765 20411 24823 20417
rect 24854 20408 24860 20420
rect 24912 20408 24918 20460
rect 24946 20408 24952 20460
rect 25004 20448 25010 20460
rect 25409 20451 25467 20457
rect 25409 20448 25421 20451
rect 25004 20420 25421 20448
rect 25004 20408 25010 20420
rect 25409 20417 25421 20420
rect 25455 20448 25467 20451
rect 26142 20448 26148 20460
rect 25455 20420 26148 20448
rect 25455 20417 25467 20420
rect 25409 20411 25467 20417
rect 26142 20408 26148 20420
rect 26200 20408 26206 20460
rect 6886 20352 22968 20380
rect 22370 20244 22376 20256
rect 22331 20216 22376 20244
rect 22370 20204 22376 20216
rect 22428 20204 22434 20256
rect 22940 20244 22968 20352
rect 24581 20383 24639 20389
rect 24581 20349 24593 20383
rect 24627 20380 24639 20383
rect 26050 20380 26056 20392
rect 24627 20352 26056 20380
rect 24627 20349 24639 20352
rect 24581 20343 24639 20349
rect 26050 20340 26056 20352
rect 26108 20340 26114 20392
rect 23109 20315 23167 20321
rect 23109 20281 23121 20315
rect 23155 20312 23167 20315
rect 38010 20312 38016 20324
rect 23155 20284 38016 20312
rect 23155 20281 23167 20284
rect 23109 20275 23167 20281
rect 38010 20272 38016 20284
rect 38068 20272 38074 20324
rect 23661 20247 23719 20253
rect 23661 20244 23673 20247
rect 22940 20216 23673 20244
rect 23661 20213 23673 20216
rect 23707 20244 23719 20247
rect 24854 20244 24860 20256
rect 23707 20216 24860 20244
rect 23707 20213 23719 20216
rect 23661 20207 23719 20213
rect 24854 20204 24860 20216
rect 24912 20204 24918 20256
rect 25222 20204 25228 20256
rect 25280 20244 25286 20256
rect 25317 20247 25375 20253
rect 25317 20244 25329 20247
rect 25280 20216 25329 20244
rect 25280 20204 25286 20216
rect 25317 20213 25329 20216
rect 25363 20213 25375 20247
rect 25317 20207 25375 20213
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 26050 20040 26056 20052
rect 26011 20012 26056 20040
rect 26050 20000 26056 20012
rect 26108 20000 26114 20052
rect 23106 19932 23112 19984
rect 23164 19972 23170 19984
rect 23164 19944 24072 19972
rect 23164 19932 23170 19944
rect 22370 19864 22376 19916
rect 22428 19904 22434 19916
rect 23569 19907 23627 19913
rect 23569 19904 23581 19907
rect 22428 19876 23581 19904
rect 22428 19864 22434 19876
rect 23569 19873 23581 19876
rect 23615 19873 23627 19907
rect 24044 19904 24072 19944
rect 24762 19932 24768 19984
rect 24820 19972 24826 19984
rect 24857 19975 24915 19981
rect 24857 19972 24869 19975
rect 24820 19944 24869 19972
rect 24820 19932 24826 19944
rect 24857 19941 24869 19944
rect 24903 19941 24915 19975
rect 24857 19935 24915 19941
rect 25409 19907 25467 19913
rect 25409 19904 25421 19907
rect 24044 19876 25421 19904
rect 23569 19867 23627 19873
rect 25409 19873 25421 19876
rect 25455 19873 25467 19907
rect 25409 19867 25467 19873
rect 21637 19839 21695 19845
rect 21637 19805 21649 19839
rect 21683 19836 21695 19839
rect 22281 19839 22339 19845
rect 22281 19836 22293 19839
rect 21683 19808 22293 19836
rect 21683 19805 21695 19808
rect 21637 19799 21695 19805
rect 22281 19805 22293 19808
rect 22327 19805 22339 19839
rect 23750 19836 23756 19848
rect 23711 19808 23756 19836
rect 22281 19799 22339 19805
rect 1670 19768 1676 19780
rect 1631 19740 1676 19768
rect 1670 19728 1676 19740
rect 1728 19728 1734 19780
rect 22296 19768 22324 19799
rect 23750 19796 23756 19808
rect 23808 19796 23814 19848
rect 26142 19836 26148 19848
rect 26103 19808 26148 19836
rect 26142 19796 26148 19808
rect 26200 19796 26206 19848
rect 25317 19771 25375 19777
rect 22296 19740 24808 19768
rect 1765 19703 1823 19709
rect 1765 19669 1777 19703
rect 1811 19700 1823 19703
rect 19426 19700 19432 19712
rect 1811 19672 19432 19700
rect 1811 19669 1823 19672
rect 1765 19663 1823 19669
rect 19426 19660 19432 19672
rect 19484 19660 19490 19712
rect 22186 19700 22192 19712
rect 22147 19672 22192 19700
rect 22186 19660 22192 19672
rect 22244 19660 22250 19712
rect 23106 19700 23112 19712
rect 23067 19672 23112 19700
rect 23106 19660 23112 19672
rect 23164 19660 23170 19712
rect 24026 19660 24032 19712
rect 24084 19700 24090 19712
rect 24670 19700 24676 19712
rect 24084 19672 24676 19700
rect 24084 19660 24090 19672
rect 24670 19660 24676 19672
rect 24728 19660 24734 19712
rect 24780 19700 24808 19740
rect 25317 19737 25329 19771
rect 25363 19768 25375 19771
rect 26602 19768 26608 19780
rect 25363 19740 26608 19768
rect 25363 19737 25375 19740
rect 25317 19731 25375 19737
rect 26602 19728 26608 19740
rect 26660 19728 26666 19780
rect 26326 19700 26332 19712
rect 24780 19672 26332 19700
rect 26326 19660 26332 19672
rect 26384 19660 26390 19712
rect 26694 19700 26700 19712
rect 26655 19672 26700 19700
rect 26694 19660 26700 19672
rect 26752 19660 26758 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 1670 19496 1676 19508
rect 1631 19468 1676 19496
rect 1670 19456 1676 19468
rect 1728 19456 1734 19508
rect 22094 19456 22100 19508
rect 22152 19496 22158 19508
rect 22649 19499 22707 19505
rect 22649 19496 22661 19499
rect 22152 19468 22661 19496
rect 22152 19456 22158 19468
rect 22649 19465 22661 19468
rect 22695 19496 22707 19499
rect 22695 19468 24164 19496
rect 22695 19465 22707 19468
rect 22649 19459 22707 19465
rect 24026 19428 24032 19440
rect 23987 19400 24032 19428
rect 24026 19388 24032 19400
rect 24084 19388 24090 19440
rect 24136 19437 24164 19468
rect 24121 19431 24179 19437
rect 24121 19397 24133 19431
rect 24167 19428 24179 19431
rect 24673 19431 24731 19437
rect 24673 19428 24685 19431
rect 24167 19400 24685 19428
rect 24167 19397 24179 19400
rect 24121 19391 24179 19397
rect 24673 19397 24685 19400
rect 24719 19397 24731 19431
rect 24673 19391 24731 19397
rect 1946 19320 1952 19372
rect 2004 19360 2010 19372
rect 9309 19363 9367 19369
rect 9309 19360 9321 19363
rect 2004 19332 9321 19360
rect 2004 19320 2010 19332
rect 9309 19329 9321 19332
rect 9355 19329 9367 19363
rect 9309 19323 9367 19329
rect 9401 19363 9459 19369
rect 9401 19329 9413 19363
rect 9447 19360 9459 19363
rect 16942 19360 16948 19372
rect 9447 19332 16948 19360
rect 9447 19329 9459 19332
rect 9401 19323 9459 19329
rect 16942 19320 16948 19332
rect 17000 19320 17006 19372
rect 20809 19363 20867 19369
rect 20809 19329 20821 19363
rect 20855 19360 20867 19363
rect 21269 19363 21327 19369
rect 21269 19360 21281 19363
rect 20855 19332 21281 19360
rect 20855 19329 20867 19332
rect 20809 19323 20867 19329
rect 21269 19329 21281 19332
rect 21315 19360 21327 19363
rect 21910 19360 21916 19372
rect 21315 19332 21916 19360
rect 21315 19329 21327 19332
rect 21269 19323 21327 19329
rect 21910 19320 21916 19332
rect 21968 19320 21974 19372
rect 22186 19360 22192 19372
rect 22147 19332 22192 19360
rect 22186 19320 22192 19332
rect 22244 19320 22250 19372
rect 24302 19320 24308 19372
rect 24360 19360 24366 19372
rect 25869 19363 25927 19369
rect 25869 19360 25881 19363
rect 24360 19332 25881 19360
rect 24360 19320 24366 19332
rect 25869 19329 25881 19332
rect 25915 19329 25927 19363
rect 25869 19323 25927 19329
rect 25961 19363 26019 19369
rect 25961 19329 25973 19363
rect 26007 19360 26019 19363
rect 26007 19332 26188 19360
rect 26007 19329 26019 19332
rect 25961 19323 26019 19329
rect 22005 19295 22063 19301
rect 22005 19261 22017 19295
rect 22051 19261 22063 19295
rect 22005 19255 22063 19261
rect 23845 19295 23903 19301
rect 23845 19261 23857 19295
rect 23891 19292 23903 19295
rect 24762 19292 24768 19304
rect 23891 19264 24768 19292
rect 23891 19261 23903 19264
rect 23845 19255 23903 19261
rect 21910 19184 21916 19236
rect 21968 19224 21974 19236
rect 22020 19224 22048 19255
rect 24762 19252 24768 19264
rect 24820 19252 24826 19304
rect 25130 19292 25136 19304
rect 25091 19264 25136 19292
rect 25130 19252 25136 19264
rect 25188 19252 25194 19304
rect 25317 19295 25375 19301
rect 25317 19261 25329 19295
rect 25363 19292 25375 19295
rect 25774 19292 25780 19304
rect 25363 19264 25780 19292
rect 25363 19261 25375 19264
rect 25317 19255 25375 19261
rect 25774 19252 25780 19264
rect 25832 19252 25838 19304
rect 26160 19292 26188 19332
rect 26234 19320 26240 19372
rect 26292 19360 26298 19372
rect 26513 19363 26571 19369
rect 26513 19360 26525 19363
rect 26292 19332 26525 19360
rect 26292 19320 26298 19332
rect 26513 19329 26525 19332
rect 26559 19329 26571 19363
rect 26513 19323 26571 19329
rect 26605 19363 26663 19369
rect 26605 19329 26617 19363
rect 26651 19360 26663 19363
rect 26694 19360 26700 19372
rect 26651 19332 26700 19360
rect 26651 19329 26663 19332
rect 26605 19323 26663 19329
rect 26694 19320 26700 19332
rect 26752 19360 26758 19372
rect 27154 19360 27160 19372
rect 26752 19332 27160 19360
rect 26752 19320 26758 19332
rect 27154 19320 27160 19332
rect 27212 19320 27218 19372
rect 33594 19320 33600 19372
rect 33652 19360 33658 19372
rect 38013 19363 38071 19369
rect 38013 19360 38025 19363
rect 33652 19332 38025 19360
rect 33652 19320 33658 19332
rect 38013 19329 38025 19332
rect 38059 19329 38071 19363
rect 38013 19323 38071 19329
rect 26326 19292 26332 19304
rect 26160 19264 26332 19292
rect 26326 19252 26332 19264
rect 26384 19292 26390 19304
rect 26384 19264 27292 19292
rect 26384 19252 26390 19264
rect 21968 19196 22048 19224
rect 21968 19184 21974 19196
rect 21358 19156 21364 19168
rect 21319 19128 21364 19156
rect 21358 19116 21364 19128
rect 21416 19116 21422 19168
rect 27264 19165 27292 19264
rect 27249 19159 27307 19165
rect 27249 19125 27261 19159
rect 27295 19156 27307 19159
rect 27338 19156 27344 19168
rect 27295 19128 27344 19156
rect 27295 19125 27307 19128
rect 27249 19119 27307 19125
rect 27338 19116 27344 19128
rect 27396 19116 27402 19168
rect 27614 19116 27620 19168
rect 27672 19156 27678 19168
rect 27709 19159 27767 19165
rect 27709 19156 27721 19159
rect 27672 19128 27721 19156
rect 27672 19116 27678 19128
rect 27709 19125 27721 19128
rect 27755 19125 27767 19159
rect 38194 19156 38200 19168
rect 38155 19128 38200 19156
rect 27709 19119 27767 19125
rect 38194 19116 38200 19128
rect 38252 19116 38258 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 19426 18912 19432 18964
rect 19484 18952 19490 18964
rect 19705 18955 19763 18961
rect 19705 18952 19717 18955
rect 19484 18924 19717 18952
rect 19484 18912 19490 18924
rect 19705 18921 19717 18924
rect 19751 18921 19763 18955
rect 19705 18915 19763 18921
rect 1854 18708 1860 18760
rect 1912 18748 1918 18760
rect 10137 18751 10195 18757
rect 10137 18748 10149 18751
rect 1912 18720 10149 18748
rect 1912 18708 1918 18720
rect 10137 18717 10149 18720
rect 10183 18748 10195 18751
rect 10781 18751 10839 18757
rect 10781 18748 10793 18751
rect 10183 18720 10793 18748
rect 10183 18717 10195 18720
rect 10137 18711 10195 18717
rect 10781 18717 10793 18720
rect 10827 18717 10839 18751
rect 19720 18748 19748 18915
rect 22094 18912 22100 18964
rect 22152 18952 22158 18964
rect 26970 18952 26976 18964
rect 22152 18924 22197 18952
rect 24504 18924 26976 18952
rect 22152 18912 22158 18924
rect 24504 18884 24532 18924
rect 26970 18912 26976 18924
rect 27028 18912 27034 18964
rect 20824 18856 24532 18884
rect 20824 18757 20852 18856
rect 24854 18844 24860 18896
rect 24912 18884 24918 18896
rect 24912 18856 26004 18884
rect 24912 18844 24918 18856
rect 21358 18776 21364 18828
rect 21416 18816 21422 18828
rect 21637 18819 21695 18825
rect 21637 18816 21649 18819
rect 21416 18788 21649 18816
rect 21416 18776 21422 18788
rect 21637 18785 21649 18788
rect 21683 18785 21695 18819
rect 22646 18816 22652 18828
rect 22607 18788 22652 18816
rect 21637 18779 21695 18785
rect 22646 18776 22652 18788
rect 22704 18776 22710 18828
rect 23750 18816 23756 18828
rect 23711 18788 23756 18816
rect 23750 18776 23756 18788
rect 23808 18776 23814 18828
rect 25133 18819 25191 18825
rect 25133 18785 25145 18819
rect 25179 18816 25191 18819
rect 25222 18816 25228 18828
rect 25179 18788 25228 18816
rect 25179 18785 25191 18788
rect 25133 18779 25191 18785
rect 25222 18776 25228 18788
rect 25280 18776 25286 18828
rect 25976 18816 26004 18856
rect 26050 18844 26056 18896
rect 26108 18884 26114 18896
rect 28261 18887 28319 18893
rect 28261 18884 28273 18887
rect 26108 18856 28273 18884
rect 26108 18844 26114 18856
rect 28261 18853 28273 18856
rect 28307 18884 28319 18887
rect 28307 18856 28994 18884
rect 28307 18853 28319 18856
rect 28261 18847 28319 18853
rect 27709 18819 27767 18825
rect 27709 18816 27721 18819
rect 25976 18788 27721 18816
rect 25976 18757 26004 18788
rect 27709 18785 27721 18788
rect 27755 18785 27767 18819
rect 28966 18816 28994 18856
rect 30190 18816 30196 18828
rect 28966 18788 30196 18816
rect 27709 18779 27767 18785
rect 30190 18776 30196 18788
rect 30248 18776 30254 18828
rect 20809 18751 20867 18757
rect 20809 18748 20821 18751
rect 19720 18720 20821 18748
rect 10781 18711 10839 18717
rect 20809 18717 20821 18720
rect 20855 18717 20867 18751
rect 20809 18711 20867 18717
rect 21453 18751 21511 18757
rect 21453 18717 21465 18751
rect 21499 18717 21511 18751
rect 25317 18751 25375 18757
rect 25317 18748 25329 18751
rect 21453 18711 21511 18717
rect 25148 18720 25329 18748
rect 10229 18683 10287 18689
rect 10229 18649 10241 18683
rect 10275 18680 10287 18683
rect 18322 18680 18328 18692
rect 10275 18652 18328 18680
rect 10275 18649 10287 18652
rect 10229 18643 10287 18649
rect 18322 18640 18328 18652
rect 18380 18640 18386 18692
rect 21468 18680 21496 18711
rect 25148 18692 25176 18720
rect 25317 18717 25329 18720
rect 25363 18748 25375 18751
rect 25869 18751 25927 18757
rect 25869 18748 25881 18751
rect 25363 18720 25881 18748
rect 25363 18717 25375 18720
rect 25317 18711 25375 18717
rect 25869 18717 25881 18720
rect 25915 18717 25927 18751
rect 25869 18711 25927 18717
rect 25961 18751 26019 18757
rect 25961 18717 25973 18751
rect 26007 18717 26019 18751
rect 25961 18711 26019 18717
rect 26605 18751 26663 18757
rect 26605 18717 26617 18751
rect 26651 18717 26663 18751
rect 27246 18748 27252 18760
rect 27159 18720 27252 18748
rect 26605 18711 26663 18717
rect 20272 18652 21496 18680
rect 20272 18624 20300 18652
rect 22002 18640 22008 18692
rect 22060 18680 22066 18692
rect 22462 18680 22468 18692
rect 22060 18652 22468 18680
rect 22060 18640 22066 18652
rect 22462 18640 22468 18652
rect 22520 18640 22526 18692
rect 22738 18640 22744 18692
rect 22796 18680 22802 18692
rect 23290 18680 23296 18692
rect 22796 18652 22841 18680
rect 23251 18652 23296 18680
rect 22796 18640 22802 18652
rect 23290 18640 23296 18652
rect 23348 18640 23354 18692
rect 24596 18652 25084 18680
rect 17494 18572 17500 18624
rect 17552 18612 17558 18624
rect 17589 18615 17647 18621
rect 17589 18612 17601 18615
rect 17552 18584 17601 18612
rect 17552 18572 17558 18584
rect 17589 18581 17601 18584
rect 17635 18581 17647 18615
rect 20254 18612 20260 18624
rect 20215 18584 20260 18612
rect 17589 18575 17647 18581
rect 20254 18572 20260 18584
rect 20312 18572 20318 18624
rect 20901 18615 20959 18621
rect 20901 18581 20913 18615
rect 20947 18612 20959 18615
rect 21910 18612 21916 18624
rect 20947 18584 21916 18612
rect 20947 18581 20959 18584
rect 20901 18575 20959 18581
rect 21910 18572 21916 18584
rect 21968 18572 21974 18624
rect 22480 18612 22508 18640
rect 24596 18612 24624 18652
rect 22480 18584 24624 18612
rect 24673 18615 24731 18621
rect 24673 18581 24685 18615
rect 24719 18612 24731 18615
rect 24946 18612 24952 18624
rect 24719 18584 24952 18612
rect 24719 18581 24731 18584
rect 24673 18575 24731 18581
rect 24946 18572 24952 18584
rect 25004 18572 25010 18624
rect 25056 18612 25084 18652
rect 25130 18640 25136 18692
rect 25188 18640 25194 18692
rect 26620 18680 26648 18711
rect 27246 18708 27252 18720
rect 27304 18748 27310 18760
rect 27304 18720 28948 18748
rect 27304 18708 27310 18720
rect 27614 18680 27620 18692
rect 25976 18652 27620 18680
rect 25976 18612 26004 18652
rect 27614 18640 27620 18652
rect 27672 18640 27678 18692
rect 26510 18612 26516 18624
rect 25056 18584 26004 18612
rect 26471 18584 26516 18612
rect 26510 18572 26516 18584
rect 26568 18572 26574 18624
rect 26694 18572 26700 18624
rect 26752 18612 26758 18624
rect 28920 18621 28948 18720
rect 27157 18615 27215 18621
rect 27157 18612 27169 18615
rect 26752 18584 27169 18612
rect 26752 18572 26758 18584
rect 27157 18581 27169 18584
rect 27203 18581 27215 18615
rect 27157 18575 27215 18581
rect 28905 18615 28963 18621
rect 28905 18581 28917 18615
rect 28951 18612 28963 18615
rect 29270 18612 29276 18624
rect 28951 18584 29276 18612
rect 28951 18581 28963 18584
rect 28905 18575 28963 18581
rect 29270 18572 29276 18584
rect 29328 18572 29334 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 2130 18368 2136 18420
rect 2188 18408 2194 18420
rect 2188 18380 24532 18408
rect 2188 18368 2194 18380
rect 17494 18340 17500 18352
rect 17455 18312 17500 18340
rect 17494 18300 17500 18312
rect 17552 18300 17558 18352
rect 17586 18300 17592 18352
rect 17644 18340 17650 18352
rect 19429 18343 19487 18349
rect 17644 18312 17689 18340
rect 17644 18300 17650 18312
rect 19429 18309 19441 18343
rect 19475 18340 19487 18343
rect 21361 18343 21419 18349
rect 19475 18312 21312 18340
rect 19475 18309 19487 18312
rect 19429 18303 19487 18309
rect 1857 18275 1915 18281
rect 1857 18241 1869 18275
rect 1903 18272 1915 18275
rect 4062 18272 4068 18284
rect 1903 18244 4068 18272
rect 1903 18241 1915 18244
rect 1857 18235 1915 18241
rect 4062 18232 4068 18244
rect 4120 18232 4126 18284
rect 18693 18275 18751 18281
rect 18693 18241 18705 18275
rect 18739 18272 18751 18275
rect 19444 18272 19472 18303
rect 20162 18272 20168 18284
rect 18739 18244 19472 18272
rect 19720 18244 20168 18272
rect 18739 18241 18751 18244
rect 18693 18235 18751 18241
rect 18138 18204 18144 18216
rect 18051 18176 18144 18204
rect 18138 18164 18144 18176
rect 18196 18204 18202 18216
rect 19720 18204 19748 18244
rect 20162 18232 20168 18244
rect 20220 18232 20226 18284
rect 21284 18281 21312 18312
rect 21361 18309 21373 18343
rect 21407 18340 21419 18343
rect 22557 18343 22615 18349
rect 22557 18340 22569 18343
rect 21407 18312 22569 18340
rect 21407 18309 21419 18312
rect 21361 18303 21419 18309
rect 22557 18309 22569 18312
rect 22603 18309 22615 18343
rect 22557 18303 22615 18309
rect 22646 18300 22652 18352
rect 22704 18340 22710 18352
rect 23382 18340 23388 18352
rect 22704 18312 22968 18340
rect 23343 18312 23388 18340
rect 22704 18300 22710 18312
rect 20441 18275 20499 18281
rect 20441 18241 20453 18275
rect 20487 18241 20499 18275
rect 20441 18235 20499 18241
rect 21269 18275 21327 18281
rect 21269 18241 21281 18275
rect 21315 18272 21327 18275
rect 21542 18272 21548 18284
rect 21315 18244 21548 18272
rect 21315 18241 21327 18244
rect 21269 18235 21327 18241
rect 19886 18204 19892 18216
rect 18196 18176 19748 18204
rect 19847 18176 19892 18204
rect 18196 18164 18202 18176
rect 19886 18164 19892 18176
rect 19944 18204 19950 18216
rect 20456 18204 20484 18235
rect 21542 18232 21548 18244
rect 21600 18232 21606 18284
rect 22646 18204 22652 18216
rect 19944 18176 20484 18204
rect 22607 18176 22652 18204
rect 19944 18164 19950 18176
rect 22646 18164 22652 18176
rect 22704 18204 22710 18216
rect 22830 18204 22836 18216
rect 22704 18176 22836 18204
rect 22704 18164 22710 18176
rect 22830 18164 22836 18176
rect 22888 18164 22894 18216
rect 22940 18204 22968 18312
rect 23382 18300 23388 18312
rect 23440 18300 23446 18352
rect 24504 18281 24532 18380
rect 27801 18343 27859 18349
rect 27801 18340 27813 18343
rect 25240 18312 27813 18340
rect 25240 18281 25268 18312
rect 27801 18309 27813 18312
rect 27847 18340 27859 18343
rect 28353 18343 28411 18349
rect 28353 18340 28365 18343
rect 27847 18312 28365 18340
rect 27847 18309 27859 18312
rect 27801 18303 27859 18309
rect 28353 18309 28365 18312
rect 28399 18309 28411 18343
rect 28353 18303 28411 18309
rect 24489 18275 24547 18281
rect 24489 18241 24501 18275
rect 24535 18272 24547 18275
rect 25225 18275 25283 18281
rect 25225 18272 25237 18275
rect 24535 18244 25237 18272
rect 24535 18241 24547 18244
rect 24489 18235 24547 18241
rect 25225 18241 25237 18244
rect 25271 18241 25283 18275
rect 25225 18235 25283 18241
rect 26421 18275 26479 18281
rect 26421 18241 26433 18275
rect 26467 18272 26479 18275
rect 26694 18272 26700 18284
rect 26467 18244 26700 18272
rect 26467 18241 26479 18244
rect 26421 18235 26479 18241
rect 26694 18232 26700 18244
rect 26752 18232 26758 18284
rect 23293 18207 23351 18213
rect 23293 18204 23305 18207
rect 22940 18176 23305 18204
rect 23293 18173 23305 18176
rect 23339 18173 23351 18207
rect 23293 18167 23351 18173
rect 23937 18207 23995 18213
rect 23937 18173 23949 18207
rect 23983 18204 23995 18207
rect 24026 18204 24032 18216
rect 23983 18176 24032 18204
rect 23983 18173 23995 18176
rect 23937 18167 23995 18173
rect 24026 18164 24032 18176
rect 24084 18164 24090 18216
rect 26605 18207 26663 18213
rect 26605 18173 26617 18207
rect 26651 18204 26663 18207
rect 27157 18207 27215 18213
rect 27157 18204 27169 18207
rect 26651 18176 27169 18204
rect 26651 18173 26663 18176
rect 26605 18167 26663 18173
rect 27157 18173 27169 18176
rect 27203 18173 27215 18207
rect 27157 18167 27215 18173
rect 18785 18139 18843 18145
rect 18785 18105 18797 18139
rect 18831 18136 18843 18139
rect 19978 18136 19984 18148
rect 18831 18108 19984 18136
rect 18831 18105 18843 18108
rect 18785 18099 18843 18105
rect 19978 18096 19984 18108
rect 20036 18096 20042 18148
rect 20162 18096 20168 18148
rect 20220 18136 20226 18148
rect 22097 18139 22155 18145
rect 22097 18136 22109 18139
rect 20220 18108 22109 18136
rect 20220 18096 20226 18108
rect 22097 18105 22109 18108
rect 22143 18105 22155 18139
rect 22097 18099 22155 18105
rect 25409 18139 25467 18145
rect 25409 18105 25421 18139
rect 25455 18136 25467 18139
rect 34422 18136 34428 18148
rect 25455 18108 34428 18136
rect 25455 18105 25467 18108
rect 25409 18099 25467 18105
rect 34422 18096 34428 18108
rect 34480 18096 34486 18148
rect 1670 18068 1676 18080
rect 1631 18040 1676 18068
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 17862 18028 17868 18080
rect 17920 18068 17926 18080
rect 19886 18068 19892 18080
rect 17920 18040 19892 18068
rect 17920 18028 17926 18040
rect 19886 18028 19892 18040
rect 19944 18028 19950 18080
rect 20533 18071 20591 18077
rect 20533 18037 20545 18071
rect 20579 18068 20591 18071
rect 20898 18068 20904 18080
rect 20579 18040 20904 18068
rect 20579 18037 20591 18040
rect 20533 18031 20591 18037
rect 20898 18028 20904 18040
rect 20956 18028 20962 18080
rect 24486 18068 24492 18080
rect 24447 18040 24492 18068
rect 24486 18028 24492 18040
rect 24544 18028 24550 18080
rect 25958 18068 25964 18080
rect 25919 18040 25964 18068
rect 25958 18028 25964 18040
rect 26016 18028 26022 18080
rect 28994 18068 29000 18080
rect 28955 18040 29000 18068
rect 28994 18028 29000 18040
rect 29052 18028 29058 18080
rect 29454 18068 29460 18080
rect 29415 18040 29460 18068
rect 29454 18028 29460 18040
rect 29512 18028 29518 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 17129 17867 17187 17873
rect 17129 17833 17141 17867
rect 17175 17864 17187 17867
rect 17586 17864 17592 17876
rect 17175 17836 17592 17864
rect 17175 17833 17187 17836
rect 17129 17827 17187 17833
rect 17586 17824 17592 17836
rect 17644 17824 17650 17876
rect 22465 17867 22523 17873
rect 22465 17833 22477 17867
rect 22511 17864 22523 17867
rect 22738 17864 22744 17876
rect 22511 17836 22744 17864
rect 22511 17833 22523 17836
rect 22465 17827 22523 17833
rect 22738 17824 22744 17836
rect 22796 17824 22802 17876
rect 23106 17824 23112 17876
rect 23164 17864 23170 17876
rect 23385 17867 23443 17873
rect 23385 17864 23397 17867
rect 23164 17836 23397 17864
rect 23164 17824 23170 17836
rect 23385 17833 23397 17836
rect 23431 17833 23443 17867
rect 23385 17827 23443 17833
rect 27522 17824 27528 17876
rect 27580 17864 27586 17876
rect 29733 17867 29791 17873
rect 29733 17864 29745 17867
rect 27580 17836 29745 17864
rect 27580 17824 27586 17836
rect 29733 17833 29745 17836
rect 29779 17833 29791 17867
rect 29733 17827 29791 17833
rect 15654 17756 15660 17808
rect 15712 17796 15718 17808
rect 19426 17796 19432 17808
rect 15712 17768 19432 17796
rect 15712 17756 15718 17768
rect 19426 17756 19432 17768
rect 19484 17796 19490 17808
rect 20254 17796 20260 17808
rect 19484 17768 20260 17796
rect 19484 17756 19490 17768
rect 20254 17756 20260 17768
rect 20312 17756 20318 17808
rect 24210 17796 24216 17808
rect 23952 17768 24216 17796
rect 17773 17731 17831 17737
rect 17773 17697 17785 17731
rect 17819 17728 17831 17731
rect 23952 17728 23980 17768
rect 24210 17756 24216 17768
rect 24268 17756 24274 17808
rect 17819 17700 23980 17728
rect 24029 17731 24087 17737
rect 17819 17697 17831 17700
rect 17773 17691 17831 17697
rect 24029 17697 24041 17731
rect 24075 17728 24087 17731
rect 24486 17728 24492 17740
rect 24075 17700 24492 17728
rect 24075 17697 24087 17700
rect 24029 17691 24087 17697
rect 16850 17620 16856 17672
rect 16908 17660 16914 17672
rect 17037 17663 17095 17669
rect 17037 17660 17049 17663
rect 16908 17632 17049 17660
rect 16908 17620 16914 17632
rect 17037 17629 17049 17632
rect 17083 17660 17095 17663
rect 17788 17660 17816 17691
rect 24486 17688 24492 17700
rect 24544 17688 24550 17740
rect 26786 17688 26792 17740
rect 26844 17728 26850 17740
rect 28721 17731 28779 17737
rect 28721 17728 28733 17731
rect 26844 17700 28733 17728
rect 26844 17688 26850 17700
rect 28721 17697 28733 17700
rect 28767 17697 28779 17731
rect 28721 17691 28779 17697
rect 20257 17663 20315 17669
rect 20257 17660 20269 17663
rect 17083 17632 17816 17660
rect 19306 17632 20269 17660
rect 17083 17629 17095 17632
rect 17037 17623 17095 17629
rect 16574 17552 16580 17604
rect 16632 17592 16638 17604
rect 18785 17595 18843 17601
rect 18785 17592 18797 17595
rect 16632 17564 18797 17592
rect 16632 17552 16638 17564
rect 18785 17561 18797 17564
rect 18831 17592 18843 17595
rect 19306 17592 19334 17632
rect 20257 17629 20269 17632
rect 20303 17660 20315 17663
rect 20438 17660 20444 17672
rect 20303 17632 20444 17660
rect 20303 17629 20315 17632
rect 20257 17623 20315 17629
rect 20438 17620 20444 17632
rect 20496 17620 20502 17672
rect 22373 17663 22431 17669
rect 22373 17660 22385 17663
rect 22066 17632 22385 17660
rect 20806 17592 20812 17604
rect 18831 17564 19334 17592
rect 20767 17564 20812 17592
rect 18831 17561 18843 17564
rect 18785 17555 18843 17561
rect 20806 17552 20812 17564
rect 20864 17552 20870 17604
rect 20898 17552 20904 17604
rect 20956 17592 20962 17604
rect 20956 17564 21001 17592
rect 20956 17552 20962 17564
rect 21082 17552 21088 17604
rect 21140 17592 21146 17604
rect 21453 17595 21511 17601
rect 21453 17592 21465 17595
rect 21140 17564 21465 17592
rect 21140 17552 21146 17564
rect 21453 17561 21465 17564
rect 21499 17561 21511 17595
rect 21453 17555 21511 17561
rect 21726 17552 21732 17604
rect 21784 17592 21790 17604
rect 21784 17564 21956 17592
rect 21784 17552 21790 17564
rect 18230 17524 18236 17536
rect 18191 17496 18236 17524
rect 18230 17484 18236 17496
rect 18288 17484 18294 17536
rect 19334 17484 19340 17536
rect 19392 17524 19398 17536
rect 19521 17527 19579 17533
rect 19521 17524 19533 17527
rect 19392 17496 19533 17524
rect 19392 17484 19398 17496
rect 19521 17493 19533 17496
rect 19567 17493 19579 17527
rect 20162 17524 20168 17536
rect 20123 17496 20168 17524
rect 19521 17487 19579 17493
rect 20162 17484 20168 17496
rect 20220 17484 20226 17536
rect 21928 17524 21956 17564
rect 22066 17524 22094 17632
rect 22373 17629 22385 17632
rect 22419 17629 22431 17663
rect 22373 17623 22431 17629
rect 23845 17663 23903 17669
rect 23845 17629 23857 17663
rect 23891 17660 23903 17663
rect 24302 17660 24308 17672
rect 23891 17632 24308 17660
rect 23891 17629 23903 17632
rect 23845 17623 23903 17629
rect 24302 17620 24308 17632
rect 24360 17620 24366 17672
rect 26050 17660 26056 17672
rect 26011 17632 26056 17660
rect 26050 17620 26056 17632
rect 26108 17620 26114 17672
rect 26878 17660 26884 17672
rect 26839 17632 26884 17660
rect 26878 17620 26884 17632
rect 26936 17620 26942 17672
rect 27522 17660 27528 17672
rect 27483 17632 27528 17660
rect 27522 17620 27528 17632
rect 27580 17620 27586 17672
rect 28166 17660 28172 17672
rect 28127 17632 28172 17660
rect 28166 17620 28172 17632
rect 28224 17620 28230 17672
rect 28813 17663 28871 17669
rect 28813 17629 28825 17663
rect 28859 17629 28871 17663
rect 28813 17623 28871 17629
rect 22646 17552 22652 17604
rect 22704 17592 22710 17604
rect 24949 17595 25007 17601
rect 24949 17592 24961 17595
rect 22704 17564 24961 17592
rect 22704 17552 22710 17564
rect 24949 17561 24961 17564
rect 24995 17561 25007 17595
rect 24949 17555 25007 17561
rect 25041 17595 25099 17601
rect 25041 17561 25053 17595
rect 25087 17561 25099 17595
rect 25590 17592 25596 17604
rect 25551 17564 25596 17592
rect 25041 17555 25099 17561
rect 21928 17496 22094 17524
rect 25056 17524 25084 17555
rect 25590 17552 25596 17564
rect 25648 17552 25654 17604
rect 26789 17595 26847 17601
rect 26789 17592 26801 17595
rect 25700 17564 26801 17592
rect 25700 17524 25728 17564
rect 26789 17561 26801 17564
rect 26835 17561 26847 17595
rect 26789 17555 26847 17561
rect 28718 17552 28724 17604
rect 28776 17592 28782 17604
rect 28828 17592 28856 17623
rect 28776 17564 28856 17592
rect 28776 17552 28782 17564
rect 25056 17496 25728 17524
rect 25774 17484 25780 17536
rect 25832 17524 25838 17536
rect 26145 17527 26203 17533
rect 26145 17524 26157 17527
rect 25832 17496 26157 17524
rect 25832 17484 25838 17496
rect 26145 17493 26157 17496
rect 26191 17524 26203 17527
rect 26326 17524 26332 17536
rect 26191 17496 26332 17524
rect 26191 17493 26203 17496
rect 26145 17487 26203 17493
rect 26326 17484 26332 17496
rect 26384 17484 26390 17536
rect 27430 17524 27436 17536
rect 27391 17496 27436 17524
rect 27430 17484 27436 17496
rect 27488 17484 27494 17536
rect 27522 17484 27528 17536
rect 27580 17524 27586 17536
rect 28077 17527 28135 17533
rect 28077 17524 28089 17527
rect 27580 17496 28089 17524
rect 27580 17484 27586 17496
rect 28077 17493 28089 17496
rect 28123 17493 28135 17527
rect 28077 17487 28135 17493
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 13078 17280 13084 17332
rect 13136 17320 13142 17332
rect 21634 17320 21640 17332
rect 13136 17292 21640 17320
rect 13136 17280 13142 17292
rect 21634 17280 21640 17292
rect 21692 17280 21698 17332
rect 21910 17280 21916 17332
rect 21968 17320 21974 17332
rect 23293 17323 23351 17329
rect 21968 17292 22140 17320
rect 21968 17280 21974 17292
rect 22112 17261 22140 17292
rect 23293 17289 23305 17323
rect 23339 17320 23351 17323
rect 23382 17320 23388 17332
rect 23339 17292 23388 17320
rect 23339 17289 23351 17292
rect 23293 17283 23351 17289
rect 23382 17280 23388 17292
rect 23440 17280 23446 17332
rect 25777 17323 25835 17329
rect 25777 17289 25789 17323
rect 25823 17320 25835 17323
rect 25958 17320 25964 17332
rect 25823 17292 25964 17320
rect 25823 17289 25835 17292
rect 25777 17283 25835 17289
rect 25958 17280 25964 17292
rect 26016 17280 26022 17332
rect 30282 17320 30288 17332
rect 27080 17292 30288 17320
rect 19521 17255 19579 17261
rect 19521 17221 19533 17255
rect 19567 17252 19579 17255
rect 22097 17255 22155 17261
rect 19567 17224 21312 17252
rect 19567 17221 19579 17224
rect 19521 17215 19579 17221
rect 1578 17144 1584 17196
rect 1636 17184 1642 17196
rect 11698 17184 11704 17196
rect 1636 17156 11704 17184
rect 1636 17144 1642 17156
rect 11698 17144 11704 17156
rect 11756 17144 11762 17196
rect 16301 17187 16359 17193
rect 16301 17153 16313 17187
rect 16347 17184 16359 17187
rect 16850 17184 16856 17196
rect 16347 17156 16856 17184
rect 16347 17153 16359 17156
rect 16301 17147 16359 17153
rect 16850 17144 16856 17156
rect 16908 17144 16914 17196
rect 19536 17184 19564 17215
rect 21284 17196 21312 17224
rect 22097 17221 22109 17255
rect 22143 17221 22155 17255
rect 22097 17215 22155 17221
rect 22186 17212 22192 17264
rect 22244 17252 22250 17264
rect 22741 17255 22799 17261
rect 22244 17224 22289 17252
rect 22244 17212 22250 17224
rect 22741 17221 22753 17255
rect 22787 17252 22799 17255
rect 24578 17252 24584 17264
rect 22787 17224 24584 17252
rect 22787 17221 22799 17224
rect 22741 17215 22799 17221
rect 24578 17212 24584 17224
rect 24636 17212 24642 17264
rect 24857 17255 24915 17261
rect 24857 17221 24869 17255
rect 24903 17252 24915 17255
rect 27080 17252 27108 17292
rect 30282 17280 30288 17292
rect 30340 17280 30346 17332
rect 28994 17252 29000 17264
rect 24903 17224 27108 17252
rect 27172 17224 29000 17252
rect 24903 17221 24915 17224
rect 24857 17215 24915 17221
rect 17604 17156 19564 17184
rect 19981 17187 20039 17193
rect 8294 17076 8300 17128
rect 8352 17116 8358 17128
rect 17604 17116 17632 17156
rect 19981 17153 19993 17187
rect 20027 17153 20039 17187
rect 19981 17147 20039 17153
rect 8352 17088 17632 17116
rect 8352 17076 8358 17088
rect 17678 17076 17684 17128
rect 17736 17116 17742 17128
rect 18969 17119 19027 17125
rect 18969 17116 18981 17119
rect 17736 17088 18981 17116
rect 17736 17076 17742 17088
rect 18969 17085 18981 17088
rect 19015 17116 19027 17119
rect 19996 17116 20024 17147
rect 20530 17144 20536 17196
rect 20588 17184 20594 17196
rect 20625 17187 20683 17193
rect 20625 17184 20637 17187
rect 20588 17156 20637 17184
rect 20588 17144 20594 17156
rect 20625 17153 20637 17156
rect 20671 17184 20683 17187
rect 20671 17156 21220 17184
rect 20671 17153 20683 17156
rect 20625 17147 20683 17153
rect 20990 17116 20996 17128
rect 19015 17088 20996 17116
rect 19015 17085 19027 17088
rect 18969 17079 19027 17085
rect 20990 17076 20996 17088
rect 21048 17076 21054 17128
rect 21192 17116 21220 17156
rect 21266 17144 21272 17196
rect 21324 17184 21330 17196
rect 23201 17187 23259 17193
rect 21324 17156 21369 17184
rect 21324 17144 21330 17156
rect 23201 17153 23213 17187
rect 23247 17153 23259 17187
rect 26234 17184 26240 17196
rect 26195 17156 26240 17184
rect 23201 17147 23259 17153
rect 21726 17116 21732 17128
rect 21192 17088 21732 17116
rect 21726 17076 21732 17088
rect 21784 17076 21790 17128
rect 21818 17076 21824 17128
rect 21876 17116 21882 17128
rect 23216 17116 23244 17147
rect 26234 17144 26240 17156
rect 26292 17144 26298 17196
rect 26418 17184 26424 17196
rect 26379 17156 26424 17184
rect 26418 17144 26424 17156
rect 26476 17144 26482 17196
rect 26510 17144 26516 17196
rect 26568 17184 26574 17196
rect 26878 17184 26884 17196
rect 26568 17156 26884 17184
rect 26568 17144 26574 17156
rect 26878 17144 26884 17156
rect 26936 17184 26942 17196
rect 27172 17193 27200 17224
rect 28994 17212 29000 17224
rect 29052 17252 29058 17264
rect 29641 17255 29699 17261
rect 29641 17252 29653 17255
rect 29052 17224 29653 17252
rect 29052 17212 29058 17224
rect 29641 17221 29653 17224
rect 29687 17221 29699 17255
rect 29641 17215 29699 17221
rect 27157 17187 27215 17193
rect 27157 17184 27169 17187
rect 26936 17156 27169 17184
rect 26936 17144 26942 17156
rect 27157 17153 27169 17156
rect 27203 17153 27215 17187
rect 27157 17147 27215 17153
rect 27985 17187 28043 17193
rect 27985 17153 27997 17187
rect 28031 17153 28043 17187
rect 27985 17147 28043 17153
rect 21876 17088 23244 17116
rect 21876 17076 21882 17088
rect 16666 17008 16672 17060
rect 16724 17048 16730 17060
rect 17770 17048 17776 17060
rect 16724 17020 17776 17048
rect 16724 17008 16730 17020
rect 17770 17008 17776 17020
rect 17828 17008 17834 17060
rect 20073 17051 20131 17057
rect 20073 17017 20085 17051
rect 20119 17048 20131 17051
rect 23216 17048 23244 17088
rect 24673 17119 24731 17125
rect 24673 17085 24685 17119
rect 24719 17116 24731 17119
rect 24762 17116 24768 17128
rect 24719 17088 24768 17116
rect 24719 17085 24731 17088
rect 24673 17079 24731 17085
rect 24762 17076 24768 17088
rect 24820 17076 24826 17128
rect 24946 17116 24952 17128
rect 24907 17088 24952 17116
rect 24946 17076 24952 17088
rect 25004 17076 25010 17128
rect 25498 17076 25504 17128
rect 25556 17116 25562 17128
rect 27522 17116 27528 17128
rect 25556 17088 27528 17116
rect 25556 17076 25562 17088
rect 27522 17076 27528 17088
rect 27580 17076 27586 17128
rect 28000 17116 28028 17147
rect 28074 17144 28080 17196
rect 28132 17184 28138 17196
rect 28626 17184 28632 17196
rect 28132 17156 28632 17184
rect 28132 17144 28138 17156
rect 28626 17144 28632 17156
rect 28684 17184 28690 17196
rect 28902 17184 28908 17196
rect 28684 17156 28908 17184
rect 28684 17144 28690 17156
rect 28902 17144 28908 17156
rect 28960 17144 28966 17196
rect 28718 17116 28724 17128
rect 28000 17088 28724 17116
rect 28718 17076 28724 17088
rect 28776 17076 28782 17128
rect 30006 17076 30012 17128
rect 30064 17116 30070 17128
rect 38013 17119 38071 17125
rect 38013 17116 38025 17119
rect 30064 17088 38025 17116
rect 30064 17076 30070 17088
rect 38013 17085 38025 17088
rect 38059 17085 38071 17119
rect 38286 17116 38292 17128
rect 38247 17088 38292 17116
rect 38013 17079 38071 17085
rect 38286 17076 38292 17088
rect 38344 17076 38350 17128
rect 28166 17048 28172 17060
rect 20119 17020 23152 17048
rect 23216 17020 28172 17048
rect 20119 17017 20131 17020
rect 20073 17011 20131 17017
rect 16945 16983 17003 16989
rect 16945 16949 16957 16983
rect 16991 16980 17003 16983
rect 17402 16980 17408 16992
rect 16991 16952 17408 16980
rect 16991 16949 17003 16952
rect 16945 16943 17003 16949
rect 17402 16940 17408 16952
rect 17460 16940 17466 16992
rect 18046 16940 18052 16992
rect 18104 16980 18110 16992
rect 18325 16983 18383 16989
rect 18325 16980 18337 16983
rect 18104 16952 18337 16980
rect 18104 16940 18110 16952
rect 18325 16949 18337 16952
rect 18371 16949 18383 16983
rect 18325 16943 18383 16949
rect 19334 16940 19340 16992
rect 19392 16980 19398 16992
rect 20530 16980 20536 16992
rect 19392 16952 20536 16980
rect 19392 16940 19398 16952
rect 20530 16940 20536 16952
rect 20588 16940 20594 16992
rect 20714 16980 20720 16992
rect 20675 16952 20720 16980
rect 20714 16940 20720 16952
rect 20772 16940 20778 16992
rect 21361 16983 21419 16989
rect 21361 16949 21373 16983
rect 21407 16980 21419 16983
rect 22554 16980 22560 16992
rect 21407 16952 22560 16980
rect 21407 16949 21419 16952
rect 21361 16943 21419 16949
rect 22554 16940 22560 16952
rect 22612 16940 22618 16992
rect 23124 16980 23152 17020
rect 28166 17008 28172 17020
rect 28224 17048 28230 17060
rect 29089 17051 29147 17057
rect 29089 17048 29101 17051
rect 28224 17020 29101 17048
rect 28224 17008 28230 17020
rect 29089 17017 29101 17020
rect 29135 17048 29147 17051
rect 29454 17048 29460 17060
rect 29135 17020 29460 17048
rect 29135 17017 29147 17020
rect 29089 17011 29147 17017
rect 29454 17008 29460 17020
rect 29512 17008 29518 17060
rect 23474 16980 23480 16992
rect 23124 16952 23480 16980
rect 23474 16940 23480 16952
rect 23532 16940 23538 16992
rect 24302 16940 24308 16992
rect 24360 16980 24366 16992
rect 24762 16980 24768 16992
rect 24360 16952 24768 16980
rect 24360 16940 24366 16952
rect 24762 16940 24768 16952
rect 24820 16940 24826 16992
rect 24854 16940 24860 16992
rect 24912 16980 24918 16992
rect 26786 16980 26792 16992
rect 24912 16952 26792 16980
rect 24912 16940 24918 16952
rect 26786 16940 26792 16952
rect 26844 16940 26850 16992
rect 27249 16983 27307 16989
rect 27249 16949 27261 16983
rect 27295 16980 27307 16983
rect 27338 16980 27344 16992
rect 27295 16952 27344 16980
rect 27295 16949 27307 16952
rect 27249 16943 27307 16949
rect 27338 16940 27344 16952
rect 27396 16940 27402 16992
rect 27890 16980 27896 16992
rect 27851 16952 27896 16980
rect 27890 16940 27896 16952
rect 27948 16940 27954 16992
rect 27982 16940 27988 16992
rect 28040 16980 28046 16992
rect 28537 16983 28595 16989
rect 28537 16980 28549 16983
rect 28040 16952 28549 16980
rect 28040 16940 28046 16952
rect 28537 16949 28549 16952
rect 28583 16949 28595 16983
rect 28537 16943 28595 16949
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 15654 16736 15660 16788
rect 15712 16776 15718 16788
rect 17037 16779 17095 16785
rect 17037 16776 17049 16779
rect 15712 16748 17049 16776
rect 15712 16736 15718 16748
rect 17037 16745 17049 16748
rect 17083 16745 17095 16779
rect 17678 16776 17684 16788
rect 17639 16748 17684 16776
rect 17037 16739 17095 16745
rect 17678 16736 17684 16748
rect 17736 16736 17742 16788
rect 21542 16776 21548 16788
rect 21503 16748 21548 16776
rect 21542 16736 21548 16748
rect 21600 16736 21606 16788
rect 21634 16736 21640 16788
rect 21692 16776 21698 16788
rect 22189 16779 22247 16785
rect 22189 16776 22201 16779
rect 21692 16748 22201 16776
rect 21692 16736 21698 16748
rect 22189 16745 22201 16748
rect 22235 16745 22247 16779
rect 22189 16739 22247 16745
rect 24762 16736 24768 16788
rect 24820 16776 24826 16788
rect 38286 16776 38292 16788
rect 24820 16748 28764 16776
rect 38247 16748 38292 16776
rect 24820 16736 24826 16748
rect 11698 16668 11704 16720
rect 11756 16708 11762 16720
rect 18141 16711 18199 16717
rect 18141 16708 18153 16711
rect 11756 16680 18153 16708
rect 11756 16668 11762 16680
rect 18141 16677 18153 16680
rect 18187 16708 18199 16711
rect 18230 16708 18236 16720
rect 18187 16680 18236 16708
rect 18187 16677 18199 16680
rect 18141 16671 18199 16677
rect 18230 16668 18236 16680
rect 18288 16708 18294 16720
rect 19334 16708 19340 16720
rect 18288 16680 19340 16708
rect 18288 16668 18294 16680
rect 19334 16668 19340 16680
rect 19392 16668 19398 16720
rect 22278 16708 22284 16720
rect 20916 16680 22284 16708
rect 17770 16600 17776 16652
rect 17828 16640 17834 16652
rect 19429 16643 19487 16649
rect 19429 16640 19441 16643
rect 17828 16612 17908 16640
rect 17828 16600 17834 16612
rect 17880 16572 17908 16612
rect 19306 16612 19441 16640
rect 18693 16575 18751 16581
rect 18693 16572 18705 16575
rect 17880 16544 18705 16572
rect 18693 16541 18705 16544
rect 18739 16541 18751 16575
rect 18693 16535 18751 16541
rect 17218 16464 17224 16516
rect 17276 16504 17282 16516
rect 19306 16504 19334 16612
rect 19429 16609 19441 16612
rect 19475 16609 19487 16643
rect 19429 16603 19487 16609
rect 20916 16581 20944 16680
rect 22278 16668 22284 16680
rect 22336 16708 22342 16720
rect 22833 16711 22891 16717
rect 22833 16708 22845 16711
rect 22336 16680 22845 16708
rect 22336 16668 22342 16680
rect 22833 16677 22845 16680
rect 22879 16677 22891 16711
rect 22833 16671 22891 16677
rect 24118 16668 24124 16720
rect 24176 16708 24182 16720
rect 24176 16680 24992 16708
rect 24176 16668 24182 16680
rect 20990 16600 20996 16652
rect 21048 16640 21054 16652
rect 23566 16640 23572 16652
rect 21048 16612 22324 16640
rect 23527 16612 23572 16640
rect 21048 16600 21054 16612
rect 20901 16575 20959 16581
rect 20901 16541 20913 16575
rect 20947 16541 20959 16575
rect 20901 16535 20959 16541
rect 19978 16504 19984 16516
rect 17276 16476 19334 16504
rect 19939 16476 19984 16504
rect 17276 16464 17282 16476
rect 19978 16464 19984 16476
rect 20036 16464 20042 16516
rect 20073 16507 20131 16513
rect 20073 16473 20085 16507
rect 20119 16473 20131 16507
rect 20073 16467 20131 16473
rect 20993 16507 21051 16513
rect 20993 16473 21005 16507
rect 21039 16504 21051 16507
rect 22186 16504 22192 16516
rect 21039 16476 22192 16504
rect 21039 16473 21051 16476
rect 20993 16467 21051 16473
rect 18782 16436 18788 16448
rect 18743 16408 18788 16436
rect 18782 16396 18788 16408
rect 18840 16396 18846 16448
rect 20088 16436 20116 16467
rect 22186 16464 22192 16476
rect 22244 16464 22250 16516
rect 22296 16513 22324 16612
rect 23566 16600 23572 16612
rect 23624 16600 23630 16652
rect 23750 16600 23756 16652
rect 23808 16640 23814 16652
rect 24964 16649 24992 16680
rect 24673 16643 24731 16649
rect 24673 16640 24685 16643
rect 23808 16612 24685 16640
rect 23808 16600 23814 16612
rect 24673 16609 24685 16612
rect 24719 16609 24731 16643
rect 24673 16603 24731 16609
rect 24949 16643 25007 16649
rect 24949 16609 24961 16643
rect 24995 16609 25007 16643
rect 24949 16603 25007 16609
rect 25958 16600 25964 16652
rect 26016 16640 26022 16652
rect 26789 16643 26847 16649
rect 26789 16640 26801 16643
rect 26016 16612 26801 16640
rect 26016 16600 26022 16612
rect 26789 16609 26801 16612
rect 26835 16640 26847 16643
rect 27341 16643 27399 16649
rect 27341 16640 27353 16643
rect 26835 16612 27353 16640
rect 26835 16609 26847 16612
rect 26789 16603 26847 16609
rect 27341 16609 27353 16612
rect 27387 16609 27399 16643
rect 27341 16603 27399 16609
rect 27801 16643 27859 16649
rect 27801 16609 27813 16643
rect 27847 16640 27859 16643
rect 28537 16643 28595 16649
rect 28537 16640 28549 16643
rect 27847 16612 28549 16640
rect 27847 16609 27859 16612
rect 27801 16603 27859 16609
rect 28537 16609 28549 16612
rect 28583 16609 28595 16643
rect 28736 16640 28764 16748
rect 38286 16736 38292 16748
rect 38344 16736 38350 16788
rect 28902 16668 28908 16720
rect 28960 16708 28966 16720
rect 29089 16711 29147 16717
rect 29089 16708 29101 16711
rect 28960 16680 29101 16708
rect 28960 16668 28966 16680
rect 29089 16677 29101 16680
rect 29135 16677 29147 16711
rect 29089 16671 29147 16677
rect 29733 16643 29791 16649
rect 29733 16640 29745 16643
rect 28537 16603 28595 16609
rect 28644 16612 29745 16640
rect 23385 16575 23443 16581
rect 23385 16541 23397 16575
rect 23431 16572 23443 16575
rect 23658 16572 23664 16584
rect 23431 16544 23664 16572
rect 23431 16541 23443 16544
rect 23385 16535 23443 16541
rect 23658 16532 23664 16544
rect 23716 16532 23722 16584
rect 27982 16572 27988 16584
rect 27943 16544 27988 16572
rect 27982 16532 27988 16544
rect 28040 16532 28046 16584
rect 28644 16581 28672 16612
rect 29733 16609 29745 16612
rect 29779 16609 29791 16643
rect 29733 16603 29791 16609
rect 28629 16575 28687 16581
rect 28629 16541 28641 16575
rect 28675 16541 28687 16575
rect 28629 16535 28687 16541
rect 22281 16507 22339 16513
rect 22281 16473 22293 16507
rect 22327 16504 22339 16507
rect 24765 16507 24823 16513
rect 22327 16476 24624 16504
rect 22327 16473 22339 16476
rect 22281 16467 22339 16473
rect 20806 16436 20812 16448
rect 20088 16408 20812 16436
rect 20806 16396 20812 16408
rect 20864 16436 20870 16448
rect 22922 16436 22928 16448
rect 20864 16408 22928 16436
rect 20864 16396 20870 16408
rect 22922 16396 22928 16408
rect 22980 16436 22986 16448
rect 23750 16436 23756 16448
rect 22980 16408 23756 16436
rect 22980 16396 22986 16408
rect 23750 16396 23756 16408
rect 23808 16396 23814 16448
rect 24029 16439 24087 16445
rect 24029 16405 24041 16439
rect 24075 16436 24087 16439
rect 24394 16436 24400 16448
rect 24075 16408 24400 16436
rect 24075 16405 24087 16408
rect 24029 16399 24087 16405
rect 24394 16396 24400 16408
rect 24452 16396 24458 16448
rect 24596 16436 24624 16476
rect 24765 16473 24777 16507
rect 24811 16504 24823 16507
rect 24854 16504 24860 16516
rect 24811 16476 24860 16504
rect 24811 16473 24823 16476
rect 24765 16467 24823 16473
rect 24854 16464 24860 16476
rect 24912 16464 24918 16516
rect 25774 16504 25780 16516
rect 25735 16476 25780 16504
rect 25774 16464 25780 16476
rect 25832 16464 25838 16516
rect 26694 16504 26700 16516
rect 26655 16476 26700 16504
rect 26694 16464 26700 16476
rect 26752 16464 26758 16516
rect 37918 16504 37924 16516
rect 26804 16476 37924 16504
rect 26804 16436 26832 16476
rect 37918 16464 37924 16476
rect 37976 16464 37982 16516
rect 24596 16408 26832 16436
rect 27246 16396 27252 16448
rect 27304 16436 27310 16448
rect 29178 16436 29184 16448
rect 27304 16408 29184 16436
rect 27304 16396 27310 16408
rect 29178 16396 29184 16408
rect 29236 16436 29242 16448
rect 30285 16439 30343 16445
rect 30285 16436 30297 16439
rect 29236 16408 30297 16436
rect 29236 16396 29242 16408
rect 30285 16405 30297 16408
rect 30331 16405 30343 16439
rect 30285 16399 30343 16405
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 18138 16232 18144 16244
rect 17604 16204 18144 16232
rect 17604 16173 17632 16204
rect 18138 16192 18144 16204
rect 18196 16192 18202 16244
rect 20622 16232 20628 16244
rect 18248 16204 20628 16232
rect 15105 16167 15163 16173
rect 15105 16133 15117 16167
rect 15151 16164 15163 16167
rect 17037 16167 17095 16173
rect 17037 16164 17049 16167
rect 15151 16136 17049 16164
rect 15151 16133 15163 16136
rect 15105 16127 15163 16133
rect 17037 16133 17049 16136
rect 17083 16133 17095 16167
rect 17037 16127 17095 16133
rect 17589 16167 17647 16173
rect 17589 16133 17601 16167
rect 17635 16133 17647 16167
rect 17589 16127 17647 16133
rect 18046 16124 18052 16176
rect 18104 16164 18110 16176
rect 18248 16164 18276 16204
rect 20622 16192 20628 16204
rect 20680 16192 20686 16244
rect 24394 16192 24400 16244
rect 24452 16232 24458 16244
rect 24762 16232 24768 16244
rect 24452 16204 24768 16232
rect 24452 16192 24458 16204
rect 24762 16192 24768 16204
rect 24820 16192 24826 16244
rect 26234 16232 26240 16244
rect 24872 16204 26240 16232
rect 18104 16136 18276 16164
rect 18325 16167 18383 16173
rect 18104 16124 18110 16136
rect 18325 16133 18337 16167
rect 18371 16164 18383 16167
rect 20162 16164 20168 16176
rect 18371 16136 20168 16164
rect 18371 16133 18383 16136
rect 18325 16127 18383 16133
rect 20162 16124 20168 16136
rect 20220 16124 20226 16176
rect 20349 16167 20407 16173
rect 20349 16133 20361 16167
rect 20395 16164 20407 16167
rect 22649 16167 22707 16173
rect 22649 16164 22661 16167
rect 20395 16136 22661 16164
rect 20395 16133 20407 16136
rect 20349 16127 20407 16133
rect 22649 16133 22661 16136
rect 22695 16133 22707 16167
rect 22649 16127 22707 16133
rect 23201 16167 23259 16173
rect 23201 16133 23213 16167
rect 23247 16164 23259 16167
rect 23290 16164 23296 16176
rect 23247 16136 23296 16164
rect 23247 16133 23259 16136
rect 23201 16127 23259 16133
rect 23290 16124 23296 16136
rect 23348 16124 23354 16176
rect 23842 16164 23848 16176
rect 23803 16136 23848 16164
rect 23842 16124 23848 16136
rect 23900 16124 23906 16176
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16096 1915 16099
rect 1903 16068 2452 16096
rect 1903 16065 1915 16068
rect 1857 16059 1915 16065
rect 2424 15904 2452 16068
rect 14734 16056 14740 16108
rect 14792 16096 14798 16108
rect 15013 16099 15071 16105
rect 15013 16096 15025 16099
rect 14792 16068 15025 16096
rect 14792 16056 14798 16068
rect 15013 16065 15025 16068
rect 15059 16065 15071 16099
rect 15013 16059 15071 16065
rect 19334 16056 19340 16108
rect 19392 16096 19398 16108
rect 19521 16099 19579 16105
rect 19521 16096 19533 16099
rect 19392 16068 19533 16096
rect 19392 16056 19398 16068
rect 19521 16065 19533 16068
rect 19567 16096 19579 16099
rect 19794 16096 19800 16108
rect 19567 16068 19800 16096
rect 19567 16065 19579 16068
rect 19521 16059 19579 16065
rect 19794 16056 19800 16068
rect 19852 16056 19858 16108
rect 19978 16056 19984 16108
rect 20036 16096 20042 16108
rect 20257 16099 20315 16105
rect 20257 16096 20269 16099
rect 20036 16068 20269 16096
rect 20036 16056 20042 16068
rect 20257 16065 20269 16068
rect 20303 16065 20315 16099
rect 20257 16059 20315 16065
rect 21085 16099 21143 16105
rect 21085 16065 21097 16099
rect 21131 16096 21143 16099
rect 21634 16096 21640 16108
rect 21131 16068 21640 16096
rect 21131 16065 21143 16068
rect 21085 16059 21143 16065
rect 21634 16056 21640 16068
rect 21692 16056 21698 16108
rect 16942 16028 16948 16040
rect 16903 16000 16948 16028
rect 16942 15988 16948 16000
rect 17000 15988 17006 16040
rect 18233 16031 18291 16037
rect 18233 15997 18245 16031
rect 18279 16028 18291 16031
rect 18690 16028 18696 16040
rect 18279 16000 18696 16028
rect 18279 15997 18291 16000
rect 18233 15991 18291 15997
rect 18690 15988 18696 16000
rect 18748 16028 18754 16040
rect 19429 16031 19487 16037
rect 19429 16028 19441 16031
rect 18748 16000 19441 16028
rect 18748 15988 18754 16000
rect 19429 15997 19441 16000
rect 19475 15997 19487 16031
rect 22554 16028 22560 16040
rect 22515 16000 22560 16028
rect 19429 15991 19487 15997
rect 22554 15988 22560 16000
rect 22612 16028 22618 16040
rect 23753 16031 23811 16037
rect 23753 16028 23765 16031
rect 22612 16000 23765 16028
rect 22612 15988 22618 16000
rect 23753 15997 23765 16000
rect 23799 15997 23811 16031
rect 24026 16028 24032 16040
rect 23987 16000 24032 16028
rect 23753 15991 23811 15997
rect 24026 15988 24032 16000
rect 24084 16028 24090 16040
rect 24872 16037 24900 16204
rect 26234 16192 26240 16204
rect 26292 16192 26298 16244
rect 26694 16192 26700 16244
rect 26752 16232 26758 16244
rect 28442 16232 28448 16244
rect 26752 16204 28448 16232
rect 26752 16192 26758 16204
rect 28442 16192 28448 16204
rect 28500 16192 28506 16244
rect 25406 16164 25412 16176
rect 25367 16136 25412 16164
rect 25406 16124 25412 16136
rect 25464 16124 25470 16176
rect 27338 16164 27344 16176
rect 27299 16136 27344 16164
rect 27338 16124 27344 16136
rect 27396 16124 27402 16176
rect 28552 16136 29868 16164
rect 28552 16105 28580 16136
rect 28537 16099 28595 16105
rect 28537 16065 28549 16099
rect 28583 16065 28595 16099
rect 29178 16096 29184 16108
rect 29139 16068 29184 16096
rect 28537 16059 28595 16065
rect 29178 16056 29184 16068
rect 29236 16056 29242 16108
rect 29840 16105 29868 16136
rect 29825 16099 29883 16105
rect 29825 16065 29837 16099
rect 29871 16096 29883 16099
rect 30469 16099 30527 16105
rect 30469 16096 30481 16099
rect 29871 16068 30481 16096
rect 29871 16065 29883 16068
rect 29825 16059 29883 16065
rect 30469 16065 30481 16068
rect 30515 16096 30527 16099
rect 30742 16096 30748 16108
rect 30515 16068 30748 16096
rect 30515 16065 30527 16068
rect 30469 16059 30527 16065
rect 30742 16056 30748 16068
rect 30800 16056 30806 16108
rect 38010 16096 38016 16108
rect 37971 16068 38016 16096
rect 38010 16056 38016 16068
rect 38068 16056 38074 16108
rect 24857 16031 24915 16037
rect 24857 16028 24869 16031
rect 24084 16000 24869 16028
rect 24084 15988 24090 16000
rect 24857 15997 24869 16000
rect 24903 15997 24915 16031
rect 24857 15991 24915 15997
rect 25501 16031 25559 16037
rect 25501 15997 25513 16031
rect 25547 16028 25559 16031
rect 26053 16031 26111 16037
rect 26053 16028 26065 16031
rect 25547 16000 26065 16028
rect 25547 15997 25559 16000
rect 25501 15991 25559 15997
rect 26053 15997 26065 16000
rect 26099 15997 26111 16031
rect 26053 15991 26111 15997
rect 26786 15988 26792 16040
rect 26844 16028 26850 16040
rect 27249 16031 27307 16037
rect 27249 16028 27261 16031
rect 26844 16000 27261 16028
rect 26844 15988 26850 16000
rect 27249 15997 27261 16000
rect 27295 16028 27307 16031
rect 27430 16028 27436 16040
rect 27295 16000 27436 16028
rect 27295 15997 27307 16000
rect 27249 15991 27307 15997
rect 27430 15988 27436 16000
rect 27488 15988 27494 16040
rect 27522 15988 27528 16040
rect 27580 16028 27586 16040
rect 29089 16031 29147 16037
rect 29089 16028 29101 16031
rect 27580 16000 27625 16028
rect 27724 16000 29101 16028
rect 27580 15988 27586 16000
rect 18785 15963 18843 15969
rect 18785 15929 18797 15963
rect 18831 15960 18843 15963
rect 18966 15960 18972 15972
rect 18831 15932 18972 15960
rect 18831 15929 18843 15932
rect 18785 15923 18843 15929
rect 18966 15920 18972 15932
rect 19024 15960 19030 15972
rect 20806 15960 20812 15972
rect 19024 15932 20812 15960
rect 19024 15920 19030 15932
rect 20806 15920 20812 15932
rect 20864 15960 20870 15972
rect 21082 15960 21088 15972
rect 20864 15932 21088 15960
rect 20864 15920 20870 15932
rect 21082 15920 21088 15932
rect 21140 15920 21146 15972
rect 25682 15920 25688 15972
rect 25740 15960 25746 15972
rect 27724 15960 27752 16000
rect 29089 15997 29101 16000
rect 29135 15997 29147 16031
rect 29089 15991 29147 15997
rect 25740 15932 27752 15960
rect 27816 15932 28580 15960
rect 25740 15920 25746 15932
rect 1670 15892 1676 15904
rect 1631 15864 1676 15892
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 2406 15892 2412 15904
rect 2367 15864 2412 15892
rect 2406 15852 2412 15864
rect 2464 15852 2470 15904
rect 16022 15852 16028 15904
rect 16080 15892 16086 15904
rect 16209 15895 16267 15901
rect 16209 15892 16221 15895
rect 16080 15864 16221 15892
rect 16080 15852 16086 15864
rect 16209 15861 16221 15864
rect 16255 15861 16267 15895
rect 16209 15855 16267 15861
rect 17770 15852 17776 15904
rect 17828 15892 17834 15904
rect 20530 15892 20536 15904
rect 17828 15864 20536 15892
rect 17828 15852 17834 15864
rect 20530 15852 20536 15864
rect 20588 15852 20594 15904
rect 20898 15892 20904 15904
rect 20859 15864 20904 15892
rect 20898 15852 20904 15864
rect 20956 15852 20962 15904
rect 25958 15852 25964 15904
rect 26016 15892 26022 15904
rect 27816 15892 27844 15932
rect 26016 15864 27844 15892
rect 26016 15852 26022 15864
rect 28166 15852 28172 15904
rect 28224 15892 28230 15904
rect 28445 15895 28503 15901
rect 28445 15892 28457 15895
rect 28224 15864 28457 15892
rect 28224 15852 28230 15864
rect 28445 15861 28457 15864
rect 28491 15861 28503 15895
rect 28552 15892 28580 15932
rect 28718 15920 28724 15972
rect 28776 15960 28782 15972
rect 29733 15963 29791 15969
rect 29733 15960 29745 15963
rect 28776 15932 29745 15960
rect 28776 15920 28782 15932
rect 29733 15929 29745 15932
rect 29779 15929 29791 15963
rect 29733 15923 29791 15929
rect 28810 15892 28816 15904
rect 28552 15864 28816 15892
rect 28445 15855 28503 15861
rect 28810 15852 28816 15864
rect 28868 15852 28874 15904
rect 29362 15852 29368 15904
rect 29420 15892 29426 15904
rect 30377 15895 30435 15901
rect 30377 15892 30389 15895
rect 29420 15864 30389 15892
rect 29420 15852 29426 15864
rect 30377 15861 30389 15864
rect 30423 15861 30435 15895
rect 38194 15892 38200 15904
rect 38155 15864 38200 15892
rect 30377 15855 30435 15861
rect 38194 15852 38200 15864
rect 38252 15852 38258 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 22281 15691 22339 15697
rect 22281 15657 22293 15691
rect 22327 15688 22339 15691
rect 23842 15688 23848 15700
rect 22327 15660 23848 15688
rect 22327 15657 22339 15660
rect 22281 15651 22339 15657
rect 23842 15648 23848 15660
rect 23900 15648 23906 15700
rect 25406 15648 25412 15700
rect 25464 15688 25470 15700
rect 28721 15691 28779 15697
rect 28721 15688 28733 15691
rect 25464 15660 28733 15688
rect 25464 15648 25470 15660
rect 28721 15657 28733 15660
rect 28767 15657 28779 15691
rect 28721 15651 28779 15657
rect 28810 15648 28816 15700
rect 28868 15688 28874 15700
rect 31297 15691 31355 15697
rect 31297 15688 31309 15691
rect 28868 15660 31309 15688
rect 28868 15648 28874 15660
rect 31297 15657 31309 15660
rect 31343 15657 31355 15691
rect 33594 15688 33600 15700
rect 33555 15660 33600 15688
rect 31297 15651 31355 15657
rect 33594 15648 33600 15660
rect 33652 15648 33658 15700
rect 38010 15688 38016 15700
rect 37971 15660 38016 15688
rect 38010 15648 38016 15660
rect 38068 15648 38074 15700
rect 2406 15580 2412 15632
rect 2464 15620 2470 15632
rect 20898 15620 20904 15632
rect 2464 15592 20904 15620
rect 2464 15580 2470 15592
rect 20898 15580 20904 15592
rect 20956 15580 20962 15632
rect 21450 15580 21456 15632
rect 21508 15620 21514 15632
rect 21910 15620 21916 15632
rect 21508 15592 21916 15620
rect 21508 15580 21514 15592
rect 21910 15580 21916 15592
rect 21968 15580 21974 15632
rect 23106 15620 23112 15632
rect 23067 15592 23112 15620
rect 23106 15580 23112 15592
rect 23164 15580 23170 15632
rect 24673 15623 24731 15629
rect 24673 15589 24685 15623
rect 24719 15620 24731 15623
rect 28534 15620 28540 15632
rect 24719 15592 28540 15620
rect 24719 15589 24731 15592
rect 24673 15583 24731 15589
rect 17218 15552 17224 15564
rect 17179 15524 17224 15552
rect 17218 15512 17224 15524
rect 17276 15512 17282 15564
rect 17497 15555 17555 15561
rect 17497 15521 17509 15555
rect 17543 15552 17555 15555
rect 18690 15552 18696 15564
rect 17543 15524 18696 15552
rect 17543 15521 17555 15524
rect 17497 15515 17555 15521
rect 18690 15512 18696 15524
rect 18748 15512 18754 15564
rect 19518 15552 19524 15564
rect 19479 15524 19524 15552
rect 19518 15512 19524 15524
rect 19576 15512 19582 15564
rect 19794 15512 19800 15564
rect 19852 15552 19858 15564
rect 19852 15524 21496 15552
rect 19852 15512 19858 15524
rect 20622 15484 20628 15496
rect 20583 15456 20628 15484
rect 20622 15444 20628 15456
rect 20680 15444 20686 15496
rect 21468 15493 21496 15524
rect 21634 15512 21640 15564
rect 21692 15552 21698 15564
rect 24688 15552 24716 15583
rect 28534 15580 28540 15592
rect 28592 15580 28598 15632
rect 31662 15620 31668 15632
rect 28644 15592 31668 15620
rect 21692 15524 24716 15552
rect 26329 15555 26387 15561
rect 21692 15512 21698 15524
rect 26329 15521 26341 15555
rect 26375 15552 26387 15555
rect 26418 15552 26424 15564
rect 26375 15524 26424 15552
rect 26375 15521 26387 15524
rect 26329 15515 26387 15521
rect 26418 15512 26424 15524
rect 26476 15512 26482 15564
rect 26513 15555 26571 15561
rect 26513 15521 26525 15555
rect 26559 15552 26571 15555
rect 27890 15552 27896 15564
rect 26559 15524 27896 15552
rect 26559 15521 26571 15524
rect 26513 15515 26571 15521
rect 27890 15512 27896 15524
rect 27948 15512 27954 15564
rect 21453 15487 21511 15493
rect 21453 15453 21465 15487
rect 21499 15453 21511 15487
rect 22186 15484 22192 15496
rect 22147 15456 22192 15484
rect 21453 15447 21511 15453
rect 22186 15444 22192 15456
rect 22244 15444 22250 15496
rect 23290 15484 23296 15496
rect 23251 15456 23296 15484
rect 23290 15444 23296 15456
rect 23348 15444 23354 15496
rect 23477 15487 23535 15493
rect 23477 15453 23489 15487
rect 23523 15484 23535 15487
rect 23658 15484 23664 15496
rect 23523 15456 23664 15484
rect 23523 15453 23535 15456
rect 23477 15447 23535 15453
rect 23658 15444 23664 15456
rect 23716 15444 23722 15496
rect 28169 15487 28227 15493
rect 28169 15453 28181 15487
rect 28215 15484 28227 15487
rect 28258 15484 28264 15496
rect 28215 15456 28264 15484
rect 28215 15453 28227 15456
rect 28169 15447 28227 15453
rect 28258 15444 28264 15456
rect 28316 15444 28322 15496
rect 28644 15484 28672 15592
rect 31662 15580 31668 15592
rect 31720 15580 31726 15632
rect 29086 15512 29092 15564
rect 29144 15552 29150 15564
rect 30469 15555 30527 15561
rect 30469 15552 30481 15555
rect 29144 15524 30481 15552
rect 29144 15512 29150 15524
rect 30469 15521 30481 15524
rect 30515 15521 30527 15555
rect 30469 15515 30527 15521
rect 31726 15524 35894 15552
rect 28460 15456 28672 15484
rect 28813 15487 28871 15493
rect 16025 15419 16083 15425
rect 16025 15416 16037 15419
rect 6886 15388 16037 15416
rect 1946 15308 1952 15360
rect 2004 15348 2010 15360
rect 6886 15348 6914 15388
rect 16025 15385 16037 15388
rect 16071 15385 16083 15419
rect 16206 15416 16212 15428
rect 16167 15388 16212 15416
rect 16025 15379 16083 15385
rect 16206 15376 16212 15388
rect 16264 15376 16270 15428
rect 17402 15416 17408 15428
rect 17363 15388 17408 15416
rect 17402 15376 17408 15388
rect 17460 15376 17466 15428
rect 17770 15376 17776 15428
rect 17828 15416 17834 15428
rect 18049 15419 18107 15425
rect 18049 15416 18061 15419
rect 17828 15388 18061 15416
rect 17828 15376 17834 15388
rect 18049 15385 18061 15388
rect 18095 15385 18107 15419
rect 18598 15416 18604 15428
rect 18559 15388 18604 15416
rect 18049 15379 18107 15385
rect 18598 15376 18604 15388
rect 18656 15376 18662 15428
rect 18874 15376 18880 15428
rect 18932 15416 18938 15428
rect 19518 15416 19524 15428
rect 18932 15388 19524 15416
rect 18932 15376 18938 15388
rect 19518 15376 19524 15388
rect 19576 15376 19582 15428
rect 19613 15419 19671 15425
rect 19613 15385 19625 15419
rect 19659 15385 19671 15419
rect 19613 15379 19671 15385
rect 2004 15320 6914 15348
rect 15565 15351 15623 15357
rect 2004 15308 2010 15320
rect 15565 15317 15577 15351
rect 15611 15348 15623 15351
rect 16224 15348 16252 15376
rect 15611 15320 16252 15348
rect 15611 15317 15623 15320
rect 15565 15311 15623 15317
rect 18782 15308 18788 15360
rect 18840 15348 18846 15360
rect 19628 15348 19656 15379
rect 19702 15376 19708 15428
rect 19760 15416 19766 15428
rect 20165 15419 20223 15425
rect 20165 15416 20177 15419
rect 19760 15388 20177 15416
rect 19760 15376 19766 15388
rect 20165 15385 20177 15388
rect 20211 15385 20223 15419
rect 25222 15416 25228 15428
rect 25183 15388 25228 15416
rect 20165 15379 20223 15385
rect 25222 15376 25228 15388
rect 25280 15376 25286 15428
rect 25317 15419 25375 15425
rect 25317 15385 25329 15419
rect 25363 15416 25375 15419
rect 25406 15416 25412 15428
rect 25363 15388 25412 15416
rect 25363 15385 25375 15388
rect 25317 15379 25375 15385
rect 25406 15376 25412 15388
rect 25464 15376 25470 15428
rect 25866 15416 25872 15428
rect 25827 15388 25872 15416
rect 25866 15376 25872 15388
rect 25924 15376 25930 15428
rect 27522 15416 27528 15428
rect 27483 15388 27528 15416
rect 27522 15376 27528 15388
rect 27580 15376 27586 15428
rect 27617 15419 27675 15425
rect 27617 15385 27629 15419
rect 27663 15416 27675 15419
rect 28460 15416 28488 15456
rect 28813 15453 28825 15487
rect 28859 15484 28871 15487
rect 29822 15484 29828 15496
rect 28859 15456 29828 15484
rect 28859 15453 28871 15456
rect 28813 15447 28871 15453
rect 29822 15444 29828 15456
rect 29880 15444 29886 15496
rect 29914 15444 29920 15496
rect 29972 15484 29978 15496
rect 30377 15487 30435 15493
rect 30377 15484 30389 15487
rect 29972 15456 30389 15484
rect 29972 15444 29978 15456
rect 30377 15453 30389 15456
rect 30423 15453 30435 15487
rect 30377 15447 30435 15453
rect 31389 15487 31447 15493
rect 31389 15453 31401 15487
rect 31435 15484 31447 15487
rect 31726 15484 31754 15524
rect 33502 15484 33508 15496
rect 31435 15456 31754 15484
rect 33463 15456 33508 15484
rect 31435 15453 31447 15456
rect 31389 15447 31447 15453
rect 33502 15444 33508 15456
rect 33560 15444 33566 15496
rect 35866 15484 35894 15524
rect 37826 15484 37832 15496
rect 35866 15456 37832 15484
rect 37826 15444 37832 15456
rect 37884 15444 37890 15496
rect 27663 15388 28488 15416
rect 27663 15385 27675 15388
rect 27617 15379 27675 15385
rect 28534 15376 28540 15428
rect 28592 15416 28598 15428
rect 37734 15416 37740 15428
rect 28592 15388 37740 15416
rect 28592 15376 28598 15388
rect 37734 15376 37740 15388
rect 37792 15376 37798 15428
rect 18840 15320 19656 15348
rect 20717 15351 20775 15357
rect 18840 15308 18846 15320
rect 20717 15317 20729 15351
rect 20763 15348 20775 15351
rect 21082 15348 21088 15360
rect 20763 15320 21088 15348
rect 20763 15317 20775 15320
rect 20717 15311 20775 15317
rect 21082 15308 21088 15320
rect 21140 15308 21146 15360
rect 21266 15348 21272 15360
rect 21227 15320 21272 15348
rect 21266 15308 21272 15320
rect 21324 15308 21330 15360
rect 21726 15308 21732 15360
rect 21784 15348 21790 15360
rect 22370 15348 22376 15360
rect 21784 15320 22376 15348
rect 21784 15308 21790 15320
rect 22370 15308 22376 15320
rect 22428 15348 22434 15360
rect 23937 15351 23995 15357
rect 23937 15348 23949 15351
rect 22428 15320 23949 15348
rect 22428 15308 22434 15320
rect 23937 15317 23949 15320
rect 23983 15317 23995 15351
rect 26970 15348 26976 15360
rect 26931 15320 26976 15348
rect 23937 15311 23995 15317
rect 26970 15308 26976 15320
rect 27028 15308 27034 15360
rect 27246 15308 27252 15360
rect 27304 15348 27310 15360
rect 29825 15351 29883 15357
rect 29825 15348 29837 15351
rect 27304 15320 29837 15348
rect 27304 15308 27310 15320
rect 29825 15317 29837 15320
rect 29871 15317 29883 15351
rect 29825 15311 29883 15317
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 16022 15104 16028 15156
rect 16080 15144 16086 15156
rect 16080 15116 17908 15144
rect 16080 15104 16086 15116
rect 16206 15036 16212 15088
rect 16264 15076 16270 15088
rect 17221 15079 17279 15085
rect 17221 15076 17233 15079
rect 16264 15048 17233 15076
rect 16264 15036 16270 15048
rect 17221 15045 17233 15048
rect 17267 15045 17279 15079
rect 17221 15039 17279 15045
rect 14734 15008 14740 15020
rect 14695 14980 14740 15008
rect 14734 14968 14740 14980
rect 14792 14968 14798 15020
rect 16117 15011 16175 15017
rect 16117 14977 16129 15011
rect 16163 15006 16175 15011
rect 17880 15008 17908 15116
rect 18598 15104 18604 15156
rect 18656 15144 18662 15156
rect 18693 15147 18751 15153
rect 18693 15144 18705 15147
rect 18656 15116 18705 15144
rect 18656 15104 18662 15116
rect 18693 15113 18705 15116
rect 18739 15113 18751 15147
rect 18693 15107 18751 15113
rect 18800 15116 19564 15144
rect 17954 15036 17960 15088
rect 18012 15076 18018 15088
rect 18800 15076 18828 15116
rect 18012 15048 18828 15076
rect 18012 15036 18018 15048
rect 19150 15036 19156 15088
rect 19208 15076 19214 15088
rect 19429 15079 19487 15085
rect 19429 15076 19441 15079
rect 19208 15048 19441 15076
rect 19208 15036 19214 15048
rect 19429 15045 19441 15048
rect 19475 15045 19487 15079
rect 19536 15076 19564 15116
rect 20070 15104 20076 15156
rect 20128 15144 20134 15156
rect 22186 15144 22192 15156
rect 20128 15116 22192 15144
rect 20128 15104 20134 15116
rect 22186 15104 22192 15116
rect 22244 15144 22250 15156
rect 22646 15144 22652 15156
rect 22244 15116 22652 15144
rect 22244 15104 22250 15116
rect 22646 15104 22652 15116
rect 22704 15104 22710 15156
rect 28166 15144 28172 15156
rect 24596 15116 28172 15144
rect 20346 15076 20352 15088
rect 19536 15048 20208 15076
rect 20307 15048 20352 15076
rect 19429 15039 19487 15045
rect 18785 15011 18843 15017
rect 18785 15008 18797 15011
rect 16224 15006 16896 15008
rect 16163 14980 16896 15006
rect 17880 14980 18797 15008
rect 16163 14978 16252 14980
rect 16163 14977 16175 14978
rect 16117 14971 16175 14977
rect 15565 14943 15623 14949
rect 15565 14909 15577 14943
rect 15611 14940 15623 14943
rect 16574 14940 16580 14952
rect 15611 14912 16580 14940
rect 15611 14909 15623 14912
rect 15565 14903 15623 14909
rect 16574 14900 16580 14912
rect 16632 14900 16638 14952
rect 14645 14875 14703 14881
rect 14645 14841 14657 14875
rect 14691 14872 14703 14875
rect 15746 14872 15752 14884
rect 14691 14844 15752 14872
rect 14691 14841 14703 14844
rect 14645 14835 14703 14841
rect 15746 14832 15752 14844
rect 15804 14832 15810 14884
rect 16758 14832 16764 14884
rect 16816 14872 16822 14884
rect 16868 14872 16896 14980
rect 18785 14977 18797 14980
rect 18831 15008 18843 15011
rect 19058 15008 19064 15020
rect 18831 14980 19064 15008
rect 18831 14977 18843 14980
rect 18785 14971 18843 14977
rect 19058 14968 19064 14980
rect 19116 14968 19122 15020
rect 20180 15008 20208 15048
rect 20346 15036 20352 15048
rect 20404 15076 20410 15088
rect 20530 15076 20536 15088
rect 20404 15048 20536 15076
rect 20404 15036 20410 15048
rect 20530 15036 20536 15048
rect 20588 15036 20594 15088
rect 20714 15036 20720 15088
rect 20772 15076 20778 15088
rect 23385 15079 23443 15085
rect 23385 15076 23397 15079
rect 20772 15048 23397 15076
rect 20772 15036 20778 15048
rect 23385 15045 23397 15048
rect 23431 15045 23443 15079
rect 23385 15039 23443 15045
rect 23474 15036 23480 15088
rect 23532 15076 23538 15088
rect 24596 15085 24624 15116
rect 28166 15104 28172 15116
rect 28224 15104 28230 15156
rect 28368 15116 28994 15144
rect 24581 15079 24639 15085
rect 23532 15048 23577 15076
rect 23532 15036 23538 15048
rect 24581 15045 24593 15079
rect 24627 15045 24639 15079
rect 24581 15039 24639 15045
rect 24946 15036 24952 15088
rect 25004 15076 25010 15088
rect 25225 15079 25283 15085
rect 25225 15076 25237 15079
rect 25004 15048 25237 15076
rect 25004 15036 25010 15048
rect 25225 15045 25237 15048
rect 25271 15045 25283 15079
rect 25225 15039 25283 15045
rect 25590 15036 25596 15088
rect 25648 15076 25654 15088
rect 27433 15079 27491 15085
rect 27433 15076 27445 15079
rect 25648 15048 27445 15076
rect 25648 15036 25654 15048
rect 27433 15045 27445 15048
rect 27479 15045 27491 15079
rect 27433 15039 27491 15045
rect 27525 15079 27583 15085
rect 27525 15045 27537 15079
rect 27571 15076 27583 15079
rect 28368 15076 28396 15116
rect 27571 15048 28396 15076
rect 28966 15076 28994 15116
rect 29454 15104 29460 15156
rect 29512 15144 29518 15156
rect 30745 15147 30803 15153
rect 30745 15144 30757 15147
rect 29512 15116 30757 15144
rect 29512 15104 29518 15116
rect 30745 15113 30757 15116
rect 30791 15113 30803 15147
rect 30745 15107 30803 15113
rect 31754 15076 31760 15088
rect 28966 15048 31760 15076
rect 27571 15045 27583 15048
rect 27525 15039 27583 15045
rect 31754 15036 31760 15048
rect 31812 15036 31818 15088
rect 20180 14980 21220 15008
rect 16942 14900 16948 14952
rect 17000 14940 17006 14952
rect 17129 14943 17187 14949
rect 17129 14940 17141 14943
rect 17000 14912 17141 14940
rect 17000 14900 17006 14912
rect 17129 14909 17141 14912
rect 17175 14909 17187 14943
rect 17129 14903 17187 14909
rect 17402 14900 17408 14952
rect 17460 14940 17466 14952
rect 18046 14940 18052 14952
rect 17460 14912 18052 14940
rect 17460 14900 17466 14912
rect 18046 14900 18052 14912
rect 18104 14900 18110 14952
rect 18138 14900 18144 14952
rect 18196 14940 18202 14952
rect 19337 14943 19395 14949
rect 19337 14940 19349 14943
rect 18196 14912 19349 14940
rect 18196 14900 18202 14912
rect 19337 14909 19349 14912
rect 19383 14909 19395 14943
rect 19337 14903 19395 14909
rect 20990 14900 20996 14952
rect 21048 14940 21054 14952
rect 21085 14943 21143 14949
rect 21085 14940 21097 14943
rect 21048 14912 21097 14940
rect 21048 14900 21054 14912
rect 21085 14909 21097 14912
rect 21131 14909 21143 14943
rect 21192 14940 21220 14980
rect 22094 14968 22100 15020
rect 22152 15008 22158 15020
rect 22189 15011 22247 15017
rect 22189 15008 22201 15011
rect 22152 14980 22201 15008
rect 22152 14968 22158 14980
rect 22189 14977 22201 14980
rect 22235 14977 22247 15011
rect 22189 14971 22247 14977
rect 24854 14968 24860 15020
rect 24912 15008 24918 15020
rect 25682 15008 25688 15020
rect 24912 14980 25544 15008
rect 25643 14980 25688 15008
rect 24912 14968 24918 14980
rect 24673 14943 24731 14949
rect 21192 14912 23428 14940
rect 21085 14903 21143 14909
rect 17586 14872 17592 14884
rect 16816 14844 17592 14872
rect 16816 14832 16822 14844
rect 17586 14832 17592 14844
rect 17644 14832 17650 14884
rect 17681 14875 17739 14881
rect 17681 14841 17693 14875
rect 17727 14872 17739 14875
rect 21174 14872 21180 14884
rect 17727 14844 21180 14872
rect 17727 14841 17739 14844
rect 17681 14835 17739 14841
rect 21174 14832 21180 14844
rect 21232 14872 21238 14884
rect 21726 14872 21732 14884
rect 21232 14844 21732 14872
rect 21232 14832 21238 14844
rect 21726 14832 21732 14844
rect 21784 14832 21790 14884
rect 22922 14872 22928 14884
rect 22883 14844 22928 14872
rect 22922 14832 22928 14844
rect 22980 14832 22986 14884
rect 23400 14872 23428 14912
rect 23584 14912 24256 14940
rect 23584 14872 23612 14912
rect 24118 14872 24124 14884
rect 23400 14844 23612 14872
rect 24079 14844 24124 14872
rect 24118 14832 24124 14844
rect 24176 14832 24182 14884
rect 24228 14872 24256 14912
rect 24673 14909 24685 14943
rect 24719 14940 24731 14943
rect 25038 14940 25044 14952
rect 24719 14912 25044 14940
rect 24719 14909 24731 14912
rect 24673 14903 24731 14909
rect 25038 14900 25044 14912
rect 25096 14900 25102 14952
rect 25516 14940 25544 14980
rect 25682 14968 25688 14980
rect 25740 14968 25746 15020
rect 26513 15011 26571 15017
rect 26513 14977 26525 15011
rect 26559 15008 26571 15011
rect 26694 15008 26700 15020
rect 26559 14980 26700 15008
rect 26559 14977 26571 14980
rect 26513 14971 26571 14977
rect 26694 14968 26700 14980
rect 26752 14968 26758 15020
rect 28077 15011 28135 15017
rect 28077 14977 28089 15011
rect 28123 15008 28135 15011
rect 28258 15008 28264 15020
rect 28123 14980 28264 15008
rect 28123 14977 28135 14980
rect 28077 14971 28135 14977
rect 28258 14968 28264 14980
rect 28316 14968 28322 15020
rect 28350 14968 28356 15020
rect 28408 15008 28414 15020
rect 28537 15011 28595 15017
rect 28537 15008 28549 15011
rect 28408 14980 28549 15008
rect 28408 14968 28414 14980
rect 28537 14977 28549 14980
rect 28583 14977 28595 15011
rect 28718 15008 28724 15020
rect 28679 14980 28724 15008
rect 28537 14971 28595 14977
rect 28718 14968 28724 14980
rect 28776 14968 28782 15020
rect 28810 14968 28816 15020
rect 28868 15014 28874 15020
rect 28868 15008 29040 15014
rect 31386 15008 31392 15020
rect 28868 14986 30420 15008
rect 28868 14968 28874 14986
rect 29012 14980 30420 14986
rect 31347 14980 31392 15008
rect 25869 14943 25927 14949
rect 25869 14940 25881 14943
rect 25516 14912 25881 14940
rect 25869 14909 25881 14912
rect 25915 14909 25927 14943
rect 25869 14903 25927 14909
rect 26050 14900 26056 14952
rect 26108 14940 26114 14952
rect 27246 14940 27252 14952
rect 26108 14912 27252 14940
rect 26108 14900 26114 14912
rect 27246 14900 27252 14912
rect 27304 14900 27310 14952
rect 30101 14943 30159 14949
rect 30101 14909 30113 14943
rect 30147 14909 30159 14943
rect 30101 14903 30159 14909
rect 26329 14875 26387 14881
rect 26329 14872 26341 14875
rect 24228 14844 26341 14872
rect 26329 14841 26341 14844
rect 26375 14841 26387 14875
rect 26329 14835 26387 14841
rect 26878 14832 26884 14884
rect 26936 14872 26942 14884
rect 26936 14844 28488 14872
rect 26936 14832 26942 14844
rect 16209 14807 16267 14813
rect 16209 14773 16221 14807
rect 16255 14804 16267 14807
rect 19242 14804 19248 14816
rect 16255 14776 19248 14804
rect 16255 14773 16267 14776
rect 16209 14767 16267 14773
rect 19242 14764 19248 14776
rect 19300 14764 19306 14816
rect 22281 14807 22339 14813
rect 22281 14773 22293 14807
rect 22327 14804 22339 14807
rect 23566 14804 23572 14816
rect 22327 14776 23572 14804
rect 22327 14773 22339 14776
rect 22281 14767 22339 14773
rect 23566 14764 23572 14776
rect 23624 14764 23630 14816
rect 23750 14764 23756 14816
rect 23808 14804 23814 14816
rect 26418 14804 26424 14816
rect 23808 14776 26424 14804
rect 23808 14764 23814 14776
rect 26418 14764 26424 14776
rect 26476 14804 26482 14816
rect 28350 14804 28356 14816
rect 26476 14776 28356 14804
rect 26476 14764 26482 14776
rect 28350 14764 28356 14776
rect 28408 14764 28414 14816
rect 28460 14804 28488 14844
rect 28810 14832 28816 14884
rect 28868 14872 28874 14884
rect 29546 14872 29552 14884
rect 28868 14844 29552 14872
rect 28868 14832 28874 14844
rect 29546 14832 29552 14844
rect 29604 14832 29610 14884
rect 30116 14872 30144 14903
rect 30190 14900 30196 14952
rect 30248 14940 30254 14952
rect 30285 14943 30343 14949
rect 30285 14940 30297 14943
rect 30248 14912 30297 14940
rect 30248 14900 30254 14912
rect 30285 14909 30297 14912
rect 30331 14909 30343 14943
rect 30392 14940 30420 14980
rect 31386 14968 31392 14980
rect 31444 14968 31450 15020
rect 31294 14940 31300 14952
rect 30392 14912 31300 14940
rect 30285 14903 30343 14909
rect 31294 14900 31300 14912
rect 31352 14900 31358 14952
rect 31481 14875 31539 14881
rect 31481 14872 31493 14875
rect 30116 14844 31493 14872
rect 31481 14841 31493 14844
rect 31527 14841 31539 14875
rect 31481 14835 31539 14841
rect 28997 14807 29055 14813
rect 28997 14804 29009 14807
rect 28460 14776 29009 14804
rect 28997 14773 29009 14776
rect 29043 14804 29055 14807
rect 29638 14804 29644 14816
rect 29043 14776 29644 14804
rect 29043 14773 29055 14776
rect 28997 14767 29055 14773
rect 29638 14764 29644 14776
rect 29696 14764 29702 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 4062 14560 4068 14612
rect 4120 14600 4126 14612
rect 9217 14603 9275 14609
rect 9217 14600 9229 14603
rect 4120 14572 9229 14600
rect 4120 14560 4126 14572
rect 9217 14569 9229 14572
rect 9263 14569 9275 14603
rect 9217 14563 9275 14569
rect 13998 14560 14004 14612
rect 14056 14600 14062 14612
rect 15105 14603 15163 14609
rect 15105 14600 15117 14603
rect 14056 14572 15117 14600
rect 14056 14560 14062 14572
rect 15105 14569 15117 14572
rect 15151 14600 15163 14603
rect 17494 14600 17500 14612
rect 15151 14572 17500 14600
rect 15151 14569 15163 14572
rect 15105 14563 15163 14569
rect 17494 14560 17500 14572
rect 17552 14600 17558 14612
rect 22094 14600 22100 14612
rect 17552 14572 22100 14600
rect 17552 14560 17558 14572
rect 22094 14560 22100 14572
rect 22152 14560 22158 14612
rect 22189 14603 22247 14609
rect 22189 14569 22201 14603
rect 22235 14600 22247 14603
rect 23290 14600 23296 14612
rect 22235 14572 23296 14600
rect 22235 14569 22247 14572
rect 22189 14563 22247 14569
rect 23290 14560 23296 14572
rect 23348 14560 23354 14612
rect 23658 14560 23664 14612
rect 23716 14600 23722 14612
rect 25682 14600 25688 14612
rect 23716 14572 25688 14600
rect 23716 14560 23722 14572
rect 25682 14560 25688 14572
rect 25740 14600 25746 14612
rect 28810 14600 28816 14612
rect 25740 14572 28816 14600
rect 25740 14560 25746 14572
rect 28810 14560 28816 14572
rect 28868 14560 28874 14612
rect 28902 14560 28908 14612
rect 28960 14600 28966 14612
rect 30469 14603 30527 14609
rect 30469 14600 30481 14603
rect 28960 14572 30481 14600
rect 28960 14560 28966 14572
rect 30469 14569 30481 14572
rect 30515 14569 30527 14603
rect 31754 14600 31760 14612
rect 31715 14572 31760 14600
rect 30469 14563 30527 14569
rect 31754 14560 31760 14572
rect 31812 14560 31818 14612
rect 32306 14600 32312 14612
rect 32267 14572 32312 14600
rect 32306 14560 32312 14572
rect 32364 14600 32370 14612
rect 38102 14600 38108 14612
rect 32364 14572 38108 14600
rect 32364 14560 32370 14572
rect 38102 14560 38108 14572
rect 38160 14560 38166 14612
rect 13725 14535 13783 14541
rect 13725 14501 13737 14535
rect 13771 14532 13783 14535
rect 16114 14532 16120 14544
rect 13771 14504 16120 14532
rect 13771 14501 13783 14504
rect 13725 14495 13783 14501
rect 16114 14492 16120 14504
rect 16172 14492 16178 14544
rect 16209 14535 16267 14541
rect 16209 14501 16221 14535
rect 16255 14532 16267 14535
rect 17218 14532 17224 14544
rect 16255 14504 17224 14532
rect 16255 14501 16267 14504
rect 16209 14495 16267 14501
rect 17218 14492 17224 14504
rect 17276 14492 17282 14544
rect 20622 14532 20628 14544
rect 17512 14504 20628 14532
rect 14553 14467 14611 14473
rect 14553 14433 14565 14467
rect 14599 14464 14611 14467
rect 17512 14464 17540 14504
rect 20622 14492 20628 14504
rect 20680 14492 20686 14544
rect 23106 14532 23112 14544
rect 23067 14504 23112 14532
rect 23106 14492 23112 14504
rect 23164 14492 23170 14544
rect 23934 14492 23940 14544
rect 23992 14532 23998 14544
rect 26786 14532 26792 14544
rect 23992 14504 26792 14532
rect 23992 14492 23998 14504
rect 26786 14492 26792 14504
rect 26844 14492 26850 14544
rect 26970 14492 26976 14544
rect 27028 14532 27034 14544
rect 27893 14535 27951 14541
rect 27893 14532 27905 14535
rect 27028 14504 27905 14532
rect 27028 14492 27034 14504
rect 27893 14501 27905 14504
rect 27939 14501 27951 14535
rect 29362 14532 29368 14544
rect 27893 14495 27951 14501
rect 28276 14504 29368 14532
rect 14599 14436 17540 14464
rect 14599 14433 14611 14436
rect 14553 14427 14611 14433
rect 1578 14396 1584 14408
rect 1539 14368 1584 14396
rect 1578 14356 1584 14368
rect 1636 14356 1642 14408
rect 1857 14399 1915 14405
rect 1857 14365 1869 14399
rect 1903 14396 1915 14399
rect 5534 14396 5540 14408
rect 1903 14368 5540 14396
rect 1903 14365 1915 14368
rect 1857 14359 1915 14365
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 9309 14399 9367 14405
rect 9309 14365 9321 14399
rect 9355 14396 9367 14399
rect 14090 14396 14096 14408
rect 9355 14368 14096 14396
rect 9355 14365 9367 14368
rect 9309 14359 9367 14365
rect 14090 14356 14096 14368
rect 14148 14356 14154 14408
rect 16853 14399 16911 14405
rect 16853 14365 16865 14399
rect 16899 14396 16911 14399
rect 17034 14396 17040 14408
rect 16899 14368 17040 14396
rect 16899 14365 16911 14368
rect 16853 14359 16911 14365
rect 15657 14331 15715 14337
rect 15657 14328 15669 14331
rect 13740 14300 15669 14328
rect 13740 14272 13768 14300
rect 15657 14297 15669 14300
rect 15703 14297 15715 14331
rect 15657 14291 15715 14297
rect 13722 14220 13728 14272
rect 13780 14220 13786 14272
rect 15672 14260 15700 14291
rect 15746 14288 15752 14340
rect 15804 14328 15810 14340
rect 15804 14300 15849 14328
rect 15804 14288 15810 14300
rect 16114 14288 16120 14340
rect 16172 14328 16178 14340
rect 16868 14328 16896 14359
rect 17034 14356 17040 14368
rect 17092 14396 17098 14408
rect 17402 14396 17408 14408
rect 17092 14368 17408 14396
rect 17092 14356 17098 14368
rect 17402 14356 17408 14368
rect 17460 14356 17466 14408
rect 17512 14405 17540 14436
rect 17586 14424 17592 14476
rect 17644 14464 17650 14476
rect 19978 14464 19984 14476
rect 17644 14436 19984 14464
rect 17644 14424 17650 14436
rect 19978 14424 19984 14436
rect 20036 14424 20042 14476
rect 23566 14464 23572 14476
rect 20824 14436 21956 14464
rect 23527 14436 23572 14464
rect 17497 14399 17555 14405
rect 17497 14365 17509 14399
rect 17543 14365 17555 14399
rect 17497 14359 17555 14365
rect 19429 14399 19487 14405
rect 19429 14365 19441 14399
rect 19475 14396 19487 14399
rect 20070 14396 20076 14408
rect 19475 14368 20076 14396
rect 19475 14365 19487 14368
rect 19429 14359 19487 14365
rect 20070 14356 20076 14368
rect 20128 14356 20134 14408
rect 20257 14399 20315 14405
rect 20257 14365 20269 14399
rect 20303 14365 20315 14399
rect 20257 14359 20315 14365
rect 16172 14300 16896 14328
rect 16945 14331 17003 14337
rect 16172 14288 16178 14300
rect 16945 14297 16957 14331
rect 16991 14328 17003 14331
rect 18046 14328 18052 14340
rect 16991 14300 18052 14328
rect 16991 14297 17003 14300
rect 16945 14291 17003 14297
rect 18046 14288 18052 14300
rect 18104 14288 18110 14340
rect 18230 14328 18236 14340
rect 18191 14300 18236 14328
rect 18230 14288 18236 14300
rect 18288 14288 18294 14340
rect 18325 14331 18383 14337
rect 18325 14297 18337 14331
rect 18371 14297 18383 14331
rect 18874 14328 18880 14340
rect 18835 14300 18880 14328
rect 18325 14291 18383 14297
rect 17402 14260 17408 14272
rect 15672 14232 17408 14260
rect 17402 14220 17408 14232
rect 17460 14220 17466 14272
rect 17586 14260 17592 14272
rect 17547 14232 17592 14260
rect 17586 14220 17592 14232
rect 17644 14220 17650 14272
rect 18340 14260 18368 14291
rect 18874 14288 18880 14300
rect 18932 14288 18938 14340
rect 20165 14331 20223 14337
rect 20165 14328 20177 14331
rect 18984 14300 20177 14328
rect 18984 14260 19012 14300
rect 20165 14297 20177 14300
rect 20211 14297 20223 14331
rect 20272 14328 20300 14359
rect 20824 14328 20852 14436
rect 21928 14396 21956 14436
rect 23566 14424 23572 14436
rect 23624 14424 23630 14476
rect 24302 14464 24308 14476
rect 23676 14436 24308 14464
rect 22002 14396 22008 14408
rect 21928 14368 22008 14396
rect 22002 14356 22008 14368
rect 22060 14356 22066 14408
rect 22094 14356 22100 14408
rect 22152 14396 22158 14408
rect 23676 14396 23704 14436
rect 24302 14424 24308 14436
rect 24360 14424 24366 14476
rect 25225 14467 25283 14473
rect 25225 14433 25237 14467
rect 25271 14464 25283 14467
rect 25406 14464 25412 14476
rect 25271 14436 25412 14464
rect 25271 14433 25283 14436
rect 25225 14427 25283 14433
rect 25406 14424 25412 14436
rect 25464 14464 25470 14476
rect 25958 14464 25964 14476
rect 25464 14436 25964 14464
rect 25464 14424 25470 14436
rect 25958 14424 25964 14436
rect 26016 14424 26022 14476
rect 26234 14424 26240 14476
rect 26292 14464 26298 14476
rect 26421 14467 26479 14473
rect 26421 14464 26433 14467
rect 26292 14436 26433 14464
rect 26292 14424 26298 14436
rect 26421 14433 26433 14436
rect 26467 14433 26479 14467
rect 26421 14427 26479 14433
rect 22152 14368 23704 14396
rect 22152 14356 22158 14368
rect 23750 14356 23756 14408
rect 23808 14396 23814 14408
rect 24578 14396 24584 14408
rect 23808 14368 23853 14396
rect 24539 14368 24584 14396
rect 23808 14356 23814 14368
rect 24578 14356 24584 14368
rect 24636 14356 24642 14408
rect 25498 14356 25504 14408
rect 25556 14396 25562 14408
rect 25777 14399 25835 14405
rect 25777 14396 25789 14399
rect 25556 14368 25789 14396
rect 25556 14356 25562 14368
rect 25777 14365 25789 14368
rect 25823 14365 25835 14399
rect 28276 14396 28304 14504
rect 29362 14492 29368 14504
rect 29420 14492 29426 14544
rect 29454 14492 29460 14544
rect 29512 14532 29518 14544
rect 29512 14504 31248 14532
rect 29512 14492 29518 14504
rect 28902 14424 28908 14476
rect 28960 14464 28966 14476
rect 31113 14467 31171 14473
rect 31113 14464 31125 14467
rect 28960 14436 31125 14464
rect 28960 14424 28966 14436
rect 31113 14433 31125 14436
rect 31159 14433 31171 14467
rect 31113 14427 31171 14433
rect 28353 14399 28411 14405
rect 28353 14396 28365 14399
rect 28276 14368 28365 14396
rect 25777 14359 25835 14365
rect 28353 14365 28365 14368
rect 28399 14365 28411 14399
rect 28353 14359 28411 14365
rect 28442 14356 28448 14408
rect 28500 14396 28506 14408
rect 28539 14399 28597 14405
rect 28539 14396 28551 14399
rect 28500 14368 28551 14396
rect 28500 14356 28506 14368
rect 28539 14365 28551 14368
rect 28585 14365 28597 14399
rect 29178 14396 29184 14408
rect 29139 14368 29184 14396
rect 28539 14359 28597 14365
rect 29178 14356 29184 14368
rect 29236 14356 29242 14408
rect 29362 14356 29368 14408
rect 29420 14396 29426 14408
rect 29917 14399 29975 14405
rect 29917 14396 29929 14399
rect 29420 14368 29929 14396
rect 29420 14356 29426 14368
rect 29917 14365 29929 14368
rect 29963 14396 29975 14399
rect 29963 14368 30052 14396
rect 29963 14365 29975 14368
rect 29917 14359 29975 14365
rect 20990 14328 20996 14340
rect 20272 14300 20852 14328
rect 20951 14300 20996 14328
rect 20165 14291 20223 14297
rect 20990 14288 20996 14300
rect 21048 14288 21054 14340
rect 21082 14288 21088 14340
rect 21140 14328 21146 14340
rect 21637 14331 21695 14337
rect 21140 14300 21185 14328
rect 21140 14288 21146 14300
rect 21637 14297 21649 14331
rect 21683 14297 21695 14331
rect 21637 14291 21695 14297
rect 18340 14232 19012 14260
rect 19521 14263 19579 14269
rect 19521 14229 19533 14263
rect 19567 14260 19579 14263
rect 20070 14260 20076 14272
rect 19567 14232 20076 14260
rect 19567 14229 19579 14232
rect 19521 14223 19579 14229
rect 20070 14220 20076 14232
rect 20128 14220 20134 14272
rect 21652 14260 21680 14291
rect 21726 14288 21732 14340
rect 21784 14328 21790 14340
rect 25133 14331 25191 14337
rect 21784 14300 23727 14328
rect 21784 14288 21790 14300
rect 22094 14260 22100 14272
rect 21652 14232 22100 14260
rect 22094 14220 22100 14232
rect 22152 14260 22158 14272
rect 23198 14260 23204 14272
rect 22152 14232 23204 14260
rect 22152 14220 22158 14232
rect 23198 14220 23204 14232
rect 23256 14220 23262 14272
rect 23699 14260 23727 14300
rect 25133 14297 25145 14331
rect 25179 14328 25191 14331
rect 26513 14331 26571 14337
rect 25179 14300 26464 14328
rect 25179 14297 25191 14300
rect 25133 14291 25191 14297
rect 25590 14260 25596 14272
rect 23699 14232 25596 14260
rect 25590 14220 25596 14232
rect 25648 14220 25654 14272
rect 26436 14260 26464 14300
rect 26513 14297 26525 14331
rect 26559 14328 26571 14331
rect 27246 14328 27252 14340
rect 26559 14300 27252 14328
rect 26559 14297 26571 14300
rect 26513 14291 26571 14297
rect 27246 14288 27252 14300
rect 27304 14288 27310 14340
rect 27430 14328 27436 14340
rect 27391 14300 27436 14328
rect 27430 14288 27436 14300
rect 27488 14288 27494 14340
rect 29825 14331 29883 14337
rect 29825 14328 29837 14331
rect 27540 14300 29837 14328
rect 27540 14260 27568 14300
rect 29825 14297 29837 14300
rect 29871 14297 29883 14331
rect 30024 14328 30052 14368
rect 30098 14356 30104 14408
rect 30156 14396 30162 14408
rect 30377 14399 30435 14405
rect 30377 14396 30389 14399
rect 30156 14368 30389 14396
rect 30156 14356 30162 14368
rect 30377 14365 30389 14368
rect 30423 14365 30435 14399
rect 30377 14359 30435 14365
rect 31021 14399 31079 14405
rect 31021 14365 31033 14399
rect 31067 14396 31079 14399
rect 31220 14396 31248 14504
rect 31067 14368 31248 14396
rect 31849 14399 31907 14405
rect 31067 14365 31079 14368
rect 31021 14359 31079 14365
rect 31849 14365 31861 14399
rect 31895 14396 31907 14399
rect 32030 14396 32036 14408
rect 31895 14368 32036 14396
rect 31895 14365 31907 14368
rect 31849 14359 31907 14365
rect 32030 14356 32036 14368
rect 32088 14356 32094 14408
rect 31570 14328 31576 14340
rect 30024 14300 31576 14328
rect 29825 14291 29883 14297
rect 31570 14288 31576 14300
rect 31628 14328 31634 14340
rect 32861 14331 32919 14337
rect 32861 14328 32873 14331
rect 31628 14300 32873 14328
rect 31628 14288 31634 14300
rect 32861 14297 32873 14300
rect 32907 14297 32919 14331
rect 32861 14291 32919 14297
rect 26436 14232 27568 14260
rect 27614 14220 27620 14272
rect 27672 14260 27678 14272
rect 28994 14260 29000 14272
rect 27672 14232 29000 14260
rect 27672 14220 27678 14232
rect 28994 14220 29000 14232
rect 29052 14220 29058 14272
rect 29089 14263 29147 14269
rect 29089 14229 29101 14263
rect 29135 14260 29147 14263
rect 29546 14260 29552 14272
rect 29135 14232 29552 14260
rect 29135 14229 29147 14232
rect 29089 14223 29147 14229
rect 29546 14220 29552 14232
rect 29604 14220 29610 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 1578 14056 1584 14068
rect 1539 14028 1584 14056
rect 1578 14016 1584 14028
rect 1636 14016 1642 14068
rect 13998 14056 14004 14068
rect 13959 14028 14004 14056
rect 13998 14016 14004 14028
rect 14056 14016 14062 14068
rect 14553 14059 14611 14065
rect 14553 14025 14565 14059
rect 14599 14056 14611 14059
rect 16022 14056 16028 14068
rect 14599 14028 16028 14056
rect 14599 14025 14611 14028
rect 14553 14019 14611 14025
rect 16022 14016 16028 14028
rect 16080 14016 16086 14068
rect 16206 14056 16212 14068
rect 16167 14028 16212 14056
rect 16206 14016 16212 14028
rect 16264 14016 16270 14068
rect 16298 14016 16304 14068
rect 16356 14056 16362 14068
rect 19978 14056 19984 14068
rect 16356 14028 19984 14056
rect 16356 14016 16362 14028
rect 19978 14016 19984 14028
rect 20036 14016 20042 14068
rect 20070 14016 20076 14068
rect 20128 14056 20134 14068
rect 20128 14028 20944 14056
rect 20128 14016 20134 14028
rect 13449 13991 13507 13997
rect 13449 13957 13461 13991
rect 13495 13988 13507 13991
rect 16390 13988 16396 14000
rect 13495 13960 16396 13988
rect 13495 13957 13507 13960
rect 13449 13951 13507 13957
rect 16390 13948 16396 13960
rect 16448 13948 16454 14000
rect 17589 13991 17647 13997
rect 17589 13957 17601 13991
rect 17635 13988 17647 13991
rect 18325 13991 18383 13997
rect 18325 13988 18337 13991
rect 17635 13960 18337 13988
rect 17635 13957 17647 13960
rect 17589 13951 17647 13957
rect 18325 13957 18337 13960
rect 18371 13957 18383 13991
rect 18325 13951 18383 13957
rect 18877 13991 18935 13997
rect 18877 13957 18889 13991
rect 18923 13988 18935 13991
rect 18966 13988 18972 14000
rect 18923 13960 18972 13988
rect 18923 13957 18935 13960
rect 18877 13951 18935 13957
rect 18966 13948 18972 13960
rect 19024 13948 19030 14000
rect 20257 13991 20315 13997
rect 20257 13957 20269 13991
rect 20303 13988 20315 13991
rect 20806 13988 20812 14000
rect 20303 13960 20812 13988
rect 20303 13957 20315 13960
rect 20257 13951 20315 13957
rect 20806 13948 20812 13960
rect 20864 13948 20870 14000
rect 20916 13997 20944 14028
rect 23474 14016 23480 14068
rect 23532 14056 23538 14068
rect 25222 14056 25228 14068
rect 23532 14028 25228 14056
rect 23532 14016 23538 14028
rect 20901 13991 20959 13997
rect 20901 13957 20913 13991
rect 20947 13957 20959 13991
rect 23842 13988 23848 14000
rect 23803 13960 23848 13988
rect 20901 13951 20959 13957
rect 23842 13948 23848 13960
rect 23900 13948 23906 14000
rect 23952 13997 23980 14028
rect 25222 14016 25228 14028
rect 25280 14016 25286 14068
rect 26329 14059 26387 14065
rect 26329 14025 26341 14059
rect 26375 14056 26387 14059
rect 26878 14056 26884 14068
rect 26375 14028 26884 14056
rect 26375 14025 26387 14028
rect 26329 14019 26387 14025
rect 26878 14016 26884 14028
rect 26936 14016 26942 14068
rect 26970 14016 26976 14068
rect 27028 14056 27034 14068
rect 27157 14059 27215 14065
rect 27157 14056 27169 14059
rect 27028 14028 27169 14056
rect 27028 14016 27034 14028
rect 27157 14025 27169 14028
rect 27203 14025 27215 14059
rect 27157 14019 27215 14025
rect 28258 14016 28264 14068
rect 28316 14016 28322 14068
rect 32401 14059 32459 14065
rect 32401 14056 32413 14059
rect 28460 14028 32413 14056
rect 23937 13991 23995 13997
rect 23937 13957 23949 13991
rect 23983 13957 23995 13991
rect 23937 13951 23995 13957
rect 25041 13991 25099 13997
rect 25041 13957 25053 13991
rect 25087 13988 25099 13991
rect 28166 13988 28172 14000
rect 25087 13960 28172 13988
rect 25087 13957 25099 13960
rect 25041 13951 25099 13957
rect 28166 13948 28172 13960
rect 28224 13948 28230 14000
rect 28276 13988 28304 14016
rect 28460 13997 28488 14028
rect 32401 14025 32413 14028
rect 32447 14025 32459 14059
rect 32401 14019 32459 14025
rect 37366 14016 37372 14068
rect 37424 14056 37430 14068
rect 38105 14059 38163 14065
rect 38105 14056 38117 14059
rect 37424 14028 38117 14056
rect 37424 14016 37430 14028
rect 38105 14025 38117 14028
rect 38151 14025 38163 14059
rect 38105 14019 38163 14025
rect 28353 13991 28411 13997
rect 28353 13988 28365 13991
rect 28276 13960 28365 13988
rect 28353 13957 28365 13960
rect 28399 13957 28411 13991
rect 28353 13951 28411 13957
rect 28445 13991 28503 13997
rect 28445 13957 28457 13991
rect 28491 13957 28503 13991
rect 28445 13951 28503 13957
rect 28534 13948 28540 14000
rect 28592 13988 28598 14000
rect 28718 13988 28724 14000
rect 28592 13960 28724 13988
rect 28592 13948 28598 13960
rect 28718 13948 28724 13960
rect 28776 13948 28782 14000
rect 29454 13948 29460 14000
rect 29512 13988 29518 14000
rect 31202 13988 31208 14000
rect 29512 13960 29868 13988
rect 31163 13960 31208 13988
rect 29512 13948 29518 13960
rect 29840 13932 29868 13960
rect 31202 13948 31208 13960
rect 31260 13948 31266 14000
rect 13722 13880 13728 13932
rect 13780 13920 13786 13932
rect 16117 13923 16175 13929
rect 16117 13920 16129 13923
rect 13780 13892 16129 13920
rect 13780 13880 13786 13892
rect 16117 13889 16129 13892
rect 16163 13889 16175 13923
rect 16117 13883 16175 13889
rect 16574 13880 16580 13932
rect 16632 13920 16638 13932
rect 17037 13923 17095 13929
rect 17037 13920 17049 13923
rect 16632 13892 17049 13920
rect 16632 13880 16638 13892
rect 17037 13889 17049 13892
rect 17083 13920 17095 13923
rect 17126 13920 17132 13932
rect 17083 13892 17132 13920
rect 17083 13889 17095 13892
rect 17037 13883 17095 13889
rect 17126 13880 17132 13892
rect 17184 13880 17190 13932
rect 17494 13920 17500 13932
rect 17455 13892 17500 13920
rect 17494 13880 17500 13892
rect 17552 13880 17558 13932
rect 19058 13880 19064 13932
rect 19116 13920 19122 13932
rect 19429 13923 19487 13929
rect 19429 13920 19441 13923
rect 19116 13892 19441 13920
rect 19116 13880 19122 13892
rect 19429 13889 19441 13892
rect 19475 13920 19487 13923
rect 20622 13920 20628 13932
rect 19475 13892 20628 13920
rect 19475 13889 19487 13892
rect 19429 13883 19487 13889
rect 20622 13880 20628 13892
rect 20680 13880 20686 13932
rect 21634 13880 21640 13932
rect 21692 13920 21698 13932
rect 22005 13923 22063 13929
rect 22005 13920 22017 13923
rect 21692 13892 22017 13920
rect 21692 13880 21698 13892
rect 22005 13889 22017 13892
rect 22051 13889 22063 13923
rect 22005 13883 22063 13889
rect 22833 13923 22891 13929
rect 22833 13889 22845 13923
rect 22879 13920 22891 13923
rect 23290 13920 23296 13932
rect 22879 13892 23296 13920
rect 22879 13889 22891 13892
rect 22833 13883 22891 13889
rect 23290 13880 23296 13892
rect 23348 13880 23354 13932
rect 25314 13880 25320 13932
rect 25372 13920 25378 13932
rect 27801 13923 27859 13929
rect 25372 13892 27752 13920
rect 25372 13880 25378 13892
rect 15105 13855 15163 13861
rect 15105 13821 15117 13855
rect 15151 13852 15163 13855
rect 16298 13852 16304 13864
rect 15151 13824 16304 13852
rect 15151 13821 15163 13824
rect 15105 13815 15163 13821
rect 16298 13812 16304 13824
rect 16356 13812 16362 13864
rect 16942 13852 16948 13864
rect 16903 13824 16948 13852
rect 16942 13812 16948 13824
rect 17000 13812 17006 13864
rect 17402 13812 17408 13864
rect 17460 13852 17466 13864
rect 18233 13855 18291 13861
rect 18233 13852 18245 13855
rect 17460 13824 18245 13852
rect 17460 13812 17466 13824
rect 18233 13821 18245 13824
rect 18279 13852 18291 13855
rect 19334 13852 19340 13864
rect 18279 13824 19340 13852
rect 18279 13821 18291 13824
rect 18233 13815 18291 13821
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 19521 13855 19579 13861
rect 19521 13821 19533 13855
rect 19567 13852 19579 13855
rect 20809 13855 20867 13861
rect 19567 13824 20760 13852
rect 19567 13821 19579 13824
rect 19521 13815 19579 13821
rect 10870 13744 10876 13796
rect 10928 13784 10934 13796
rect 17954 13784 17960 13796
rect 10928 13756 17960 13784
rect 10928 13744 10934 13756
rect 17954 13744 17960 13756
rect 18012 13744 18018 13796
rect 20732 13784 20760 13824
rect 20809 13821 20821 13855
rect 20855 13852 20867 13855
rect 22097 13855 22155 13861
rect 20855 13824 21036 13852
rect 20855 13821 20867 13824
rect 20809 13815 20867 13821
rect 20898 13784 20904 13796
rect 20732 13756 20904 13784
rect 20898 13744 20904 13756
rect 20956 13744 20962 13796
rect 15562 13716 15568 13728
rect 15523 13688 15568 13716
rect 15562 13676 15568 13688
rect 15620 13676 15626 13728
rect 15746 13676 15752 13728
rect 15804 13716 15810 13728
rect 19426 13716 19432 13728
rect 15804 13688 19432 13716
rect 15804 13676 15810 13688
rect 19426 13676 19432 13688
rect 19484 13676 19490 13728
rect 19518 13676 19524 13728
rect 19576 13716 19582 13728
rect 21008 13716 21036 13824
rect 22097 13821 22109 13855
rect 22143 13852 22155 13855
rect 23474 13852 23480 13864
rect 22143 13824 23480 13852
rect 22143 13821 22155 13824
rect 22097 13815 22155 13821
rect 23474 13812 23480 13824
rect 23532 13812 23538 13864
rect 23661 13855 23719 13861
rect 23661 13821 23673 13855
rect 23707 13852 23719 13855
rect 23750 13852 23756 13864
rect 23707 13824 23756 13852
rect 23707 13821 23719 13824
rect 23661 13815 23719 13821
rect 23750 13812 23756 13824
rect 23808 13852 23814 13864
rect 24489 13855 24547 13861
rect 24489 13852 24501 13855
rect 23808 13824 23888 13852
rect 23808 13812 23814 13824
rect 21361 13787 21419 13793
rect 21361 13753 21373 13787
rect 21407 13784 21419 13787
rect 23382 13784 23388 13796
rect 21407 13756 23388 13784
rect 21407 13753 21419 13756
rect 21361 13747 21419 13753
rect 23382 13744 23388 13756
rect 23440 13744 23446 13796
rect 23860 13784 23888 13824
rect 24044 13824 24501 13852
rect 24044 13784 24072 13824
rect 24489 13821 24501 13824
rect 24535 13821 24547 13855
rect 25130 13852 25136 13864
rect 25043 13824 25136 13852
rect 24489 13815 24547 13821
rect 25130 13812 25136 13824
rect 25188 13852 25194 13864
rect 25406 13852 25412 13864
rect 25188 13824 25412 13852
rect 25188 13812 25194 13824
rect 25406 13812 25412 13824
rect 25464 13812 25470 13864
rect 25682 13852 25688 13864
rect 25643 13824 25688 13852
rect 25682 13812 25688 13824
rect 25740 13812 25746 13864
rect 25869 13855 25927 13861
rect 25869 13821 25881 13855
rect 25915 13852 25927 13855
rect 26050 13852 26056 13864
rect 25915 13824 26056 13852
rect 25915 13821 25927 13824
rect 25869 13815 25927 13821
rect 26050 13812 26056 13824
rect 26108 13812 26114 13864
rect 26602 13812 26608 13864
rect 26660 13852 26666 13864
rect 27154 13852 27160 13864
rect 26660 13824 27160 13852
rect 26660 13812 26666 13824
rect 27154 13812 27160 13824
rect 27212 13812 27218 13864
rect 27614 13852 27620 13864
rect 27575 13824 27620 13852
rect 27614 13812 27620 13824
rect 27672 13812 27678 13864
rect 27724 13852 27752 13892
rect 27801 13889 27813 13923
rect 27847 13920 27859 13923
rect 27982 13920 27988 13932
rect 27847 13892 27988 13920
rect 27847 13889 27859 13892
rect 27801 13883 27859 13889
rect 27982 13880 27988 13892
rect 28040 13880 28046 13932
rect 29641 13923 29699 13929
rect 29641 13889 29653 13923
rect 29687 13889 29699 13923
rect 29641 13883 29699 13889
rect 29178 13852 29184 13864
rect 27724 13824 29184 13852
rect 29178 13812 29184 13824
rect 29236 13812 29242 13864
rect 28166 13784 28172 13796
rect 23860 13756 24072 13784
rect 26528 13756 28172 13784
rect 22738 13716 22744 13728
rect 19576 13688 21036 13716
rect 22699 13688 22744 13716
rect 19576 13676 19582 13688
rect 22738 13676 22744 13688
rect 22796 13676 22802 13728
rect 24854 13676 24860 13728
rect 24912 13716 24918 13728
rect 26528 13716 26556 13756
rect 28166 13744 28172 13756
rect 28224 13744 28230 13796
rect 28902 13784 28908 13796
rect 28863 13756 28908 13784
rect 28902 13744 28908 13756
rect 28960 13744 28966 13796
rect 28994 13744 29000 13796
rect 29052 13784 29058 13796
rect 29656 13784 29684 13883
rect 29822 13880 29828 13932
rect 29880 13920 29886 13932
rect 30101 13923 30159 13929
rect 30101 13920 30113 13923
rect 29880 13892 30113 13920
rect 29880 13880 29886 13892
rect 30101 13889 30113 13892
rect 30147 13889 30159 13923
rect 30101 13883 30159 13889
rect 32493 13923 32551 13929
rect 32493 13889 32505 13923
rect 32539 13920 32551 13923
rect 32582 13920 32588 13932
rect 32539 13892 32588 13920
rect 32539 13889 32551 13892
rect 32493 13883 32551 13889
rect 32582 13880 32588 13892
rect 32640 13880 32646 13932
rect 37553 13923 37611 13929
rect 37553 13889 37565 13923
rect 37599 13920 37611 13923
rect 38286 13920 38292 13932
rect 37599 13892 38292 13920
rect 37599 13889 37611 13892
rect 37553 13883 37611 13889
rect 38286 13880 38292 13892
rect 38344 13880 38350 13932
rect 29914 13812 29920 13864
rect 29972 13852 29978 13864
rect 30193 13855 30251 13861
rect 30193 13852 30205 13855
rect 29972 13824 30205 13852
rect 29972 13812 29978 13824
rect 30193 13821 30205 13824
rect 30239 13821 30251 13855
rect 31110 13852 31116 13864
rect 31071 13824 31116 13852
rect 30193 13815 30251 13821
rect 31110 13812 31116 13824
rect 31168 13812 31174 13864
rect 32953 13855 33011 13861
rect 32953 13852 32965 13855
rect 31220 13824 32965 13852
rect 31220 13784 31248 13824
rect 32953 13821 32965 13824
rect 32999 13821 33011 13855
rect 32953 13815 33011 13821
rect 29052 13756 31248 13784
rect 29052 13744 29058 13756
rect 31294 13744 31300 13796
rect 31352 13784 31358 13796
rect 31665 13787 31723 13793
rect 31665 13784 31677 13787
rect 31352 13756 31677 13784
rect 31352 13744 31358 13756
rect 31665 13753 31677 13756
rect 31711 13753 31723 13787
rect 31665 13747 31723 13753
rect 31754 13744 31760 13796
rect 31812 13784 31818 13796
rect 35526 13784 35532 13796
rect 31812 13756 35532 13784
rect 31812 13744 31818 13756
rect 35526 13744 35532 13756
rect 35584 13744 35590 13796
rect 24912 13688 26556 13716
rect 24912 13676 24918 13688
rect 27246 13676 27252 13728
rect 27304 13716 27310 13728
rect 29549 13719 29607 13725
rect 29549 13716 29561 13719
rect 27304 13688 29561 13716
rect 27304 13676 27310 13688
rect 29549 13685 29561 13688
rect 29595 13685 29607 13719
rect 29549 13679 29607 13685
rect 29730 13676 29736 13728
rect 29788 13716 29794 13728
rect 30190 13716 30196 13728
rect 29788 13688 30196 13716
rect 29788 13676 29794 13688
rect 30190 13676 30196 13688
rect 30248 13676 30254 13728
rect 30466 13676 30472 13728
rect 30524 13716 30530 13728
rect 33502 13716 33508 13728
rect 30524 13688 33508 13716
rect 30524 13676 30530 13688
rect 33502 13676 33508 13688
rect 33560 13676 33566 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 13722 13512 13728 13524
rect 13683 13484 13728 13512
rect 13722 13472 13728 13484
rect 13780 13472 13786 13524
rect 14737 13515 14795 13521
rect 14737 13481 14749 13515
rect 14783 13512 14795 13515
rect 15654 13512 15660 13524
rect 14783 13484 15660 13512
rect 14783 13481 14795 13484
rect 14737 13475 14795 13481
rect 15654 13472 15660 13484
rect 15712 13512 15718 13524
rect 15712 13484 18644 13512
rect 15712 13472 15718 13484
rect 15933 13447 15991 13453
rect 15933 13413 15945 13447
rect 15979 13444 15991 13447
rect 18506 13444 18512 13456
rect 15979 13416 18512 13444
rect 15979 13413 15991 13416
rect 15933 13407 15991 13413
rect 18506 13404 18512 13416
rect 18564 13404 18570 13456
rect 2314 13336 2320 13388
rect 2372 13376 2378 13388
rect 10870 13376 10876 13388
rect 2372 13348 10876 13376
rect 2372 13336 2378 13348
rect 10870 13336 10876 13348
rect 10928 13336 10934 13388
rect 12621 13379 12679 13385
rect 12621 13345 12633 13379
rect 12667 13376 12679 13379
rect 15746 13376 15752 13388
rect 12667 13348 15752 13376
rect 12667 13345 12679 13348
rect 12621 13339 12679 13345
rect 15746 13336 15752 13348
rect 15804 13336 15810 13388
rect 17494 13336 17500 13388
rect 17552 13376 17558 13388
rect 17957 13379 18015 13385
rect 17957 13376 17969 13379
rect 17552 13348 17969 13376
rect 17552 13336 17558 13348
rect 17957 13345 17969 13348
rect 18003 13376 18015 13379
rect 18230 13376 18236 13388
rect 18003 13348 18236 13376
rect 18003 13345 18015 13348
rect 17957 13339 18015 13345
rect 18230 13336 18236 13348
rect 18288 13336 18294 13388
rect 18616 13376 18644 13484
rect 21450 13472 21456 13524
rect 21508 13512 21514 13524
rect 24118 13512 24124 13524
rect 21508 13484 24124 13512
rect 21508 13472 21514 13484
rect 24118 13472 24124 13484
rect 24176 13472 24182 13524
rect 27154 13512 27160 13524
rect 24964 13484 27160 13512
rect 18782 13404 18788 13456
rect 18840 13444 18846 13456
rect 20073 13447 20131 13453
rect 20073 13444 20085 13447
rect 18840 13416 20085 13444
rect 18840 13404 18846 13416
rect 20073 13413 20085 13416
rect 20119 13444 20131 13447
rect 22922 13444 22928 13456
rect 20119 13416 22928 13444
rect 20119 13413 20131 13416
rect 20073 13407 20131 13413
rect 22922 13404 22928 13416
rect 22980 13404 22986 13456
rect 23014 13404 23020 13456
rect 23072 13444 23078 13456
rect 23072 13416 24900 13444
rect 23072 13404 23078 13416
rect 19518 13376 19524 13388
rect 18616 13348 19524 13376
rect 19518 13336 19524 13348
rect 19576 13336 19582 13388
rect 20806 13376 20812 13388
rect 20767 13348 20812 13376
rect 20806 13336 20812 13348
rect 20864 13336 20870 13388
rect 21174 13376 21180 13388
rect 21135 13348 21180 13376
rect 21174 13336 21180 13348
rect 21232 13336 21238 13388
rect 21910 13336 21916 13388
rect 21968 13376 21974 13388
rect 22281 13379 22339 13385
rect 22281 13376 22293 13379
rect 21968 13348 22293 13376
rect 21968 13336 21974 13348
rect 22281 13345 22293 13348
rect 22327 13345 22339 13379
rect 22281 13339 22339 13345
rect 23106 13336 23112 13388
rect 23164 13376 23170 13388
rect 23290 13376 23296 13388
rect 23164 13348 23296 13376
rect 23164 13336 23170 13348
rect 23290 13336 23296 13348
rect 23348 13336 23354 13388
rect 24872 13385 24900 13416
rect 24857 13379 24915 13385
rect 24857 13345 24869 13379
rect 24903 13345 24915 13379
rect 24857 13339 24915 13345
rect 13354 13268 13360 13320
rect 13412 13308 13418 13320
rect 15197 13311 15255 13317
rect 15197 13308 15209 13311
rect 13412 13280 15209 13308
rect 13412 13268 13418 13280
rect 15197 13277 15209 13280
rect 15243 13277 15255 13311
rect 15764 13308 15792 13336
rect 15841 13311 15899 13317
rect 15841 13308 15853 13311
rect 15764 13280 15853 13308
rect 15197 13271 15255 13277
rect 15841 13277 15853 13280
rect 15887 13277 15899 13311
rect 15841 13271 15899 13277
rect 16485 13311 16543 13317
rect 16485 13277 16497 13311
rect 16531 13277 16543 13311
rect 16485 13271 16543 13277
rect 16577 13311 16635 13317
rect 16577 13277 16589 13311
rect 16623 13308 16635 13311
rect 17678 13308 17684 13320
rect 16623 13280 17684 13308
rect 16623 13277 16635 13280
rect 16577 13271 16635 13277
rect 13173 13243 13231 13249
rect 13173 13209 13185 13243
rect 13219 13240 13231 13243
rect 13814 13240 13820 13252
rect 13219 13212 13820 13240
rect 13219 13209 13231 13212
rect 13173 13203 13231 13209
rect 13814 13200 13820 13212
rect 13872 13240 13878 13252
rect 16500 13240 16528 13271
rect 17678 13268 17684 13280
rect 17736 13268 17742 13320
rect 24029 13311 24087 13317
rect 24029 13277 24041 13311
rect 24075 13308 24087 13311
rect 24964 13308 24992 13484
rect 27154 13472 27160 13484
rect 27212 13472 27218 13524
rect 28902 13472 28908 13524
rect 28960 13512 28966 13524
rect 30466 13512 30472 13524
rect 28960 13484 30472 13512
rect 28960 13472 28966 13484
rect 30466 13472 30472 13484
rect 30524 13472 30530 13524
rect 30558 13472 30564 13524
rect 30616 13512 30622 13524
rect 31021 13515 31079 13521
rect 31021 13512 31033 13515
rect 30616 13484 31033 13512
rect 30616 13472 30622 13484
rect 31021 13481 31033 13484
rect 31067 13481 31079 13515
rect 31662 13512 31668 13524
rect 31623 13484 31668 13512
rect 31021 13475 31079 13481
rect 31662 13472 31668 13484
rect 31720 13472 31726 13524
rect 25406 13404 25412 13456
rect 25464 13444 25470 13456
rect 25464 13416 27476 13444
rect 25464 13404 25470 13416
rect 25774 13336 25780 13388
rect 25832 13376 25838 13388
rect 27246 13376 27252 13388
rect 25832 13348 27252 13376
rect 25832 13336 25838 13348
rect 27246 13336 27252 13348
rect 27304 13336 27310 13388
rect 24075 13280 24992 13308
rect 27448 13308 27476 13416
rect 28166 13404 28172 13456
rect 28224 13444 28230 13456
rect 29730 13444 29736 13456
rect 28224 13416 29736 13444
rect 28224 13404 28230 13416
rect 29730 13404 29736 13416
rect 29788 13404 29794 13456
rect 29822 13404 29828 13456
rect 29880 13444 29886 13456
rect 31754 13444 31760 13456
rect 29880 13416 31760 13444
rect 29880 13404 29886 13416
rect 31754 13404 31760 13416
rect 31812 13404 31818 13456
rect 27614 13336 27620 13388
rect 27672 13376 27678 13388
rect 28994 13376 29000 13388
rect 27672 13348 29000 13376
rect 27672 13336 27678 13348
rect 28994 13336 29000 13348
rect 29052 13336 29058 13388
rect 32953 13379 33011 13385
rect 32953 13376 32965 13379
rect 29104 13348 32965 13376
rect 27448 13280 27752 13308
rect 24075 13277 24087 13280
rect 24029 13271 24087 13277
rect 17310 13240 17316 13252
rect 13872 13212 16528 13240
rect 17271 13212 17316 13240
rect 13872 13200 13878 13212
rect 17310 13200 17316 13212
rect 17368 13200 17374 13252
rect 18046 13200 18052 13252
rect 18104 13240 18110 13252
rect 18104 13212 18149 13240
rect 18104 13200 18110 13212
rect 18322 13200 18328 13252
rect 18380 13240 18386 13252
rect 18601 13243 18659 13249
rect 18601 13240 18613 13243
rect 18380 13212 18613 13240
rect 18380 13200 18386 13212
rect 18601 13209 18613 13212
rect 18647 13240 18659 13243
rect 18782 13240 18788 13252
rect 18647 13212 18788 13240
rect 18647 13209 18659 13212
rect 18601 13203 18659 13209
rect 18782 13200 18788 13212
rect 18840 13200 18846 13252
rect 19613 13243 19671 13249
rect 19613 13209 19625 13243
rect 19659 13209 19671 13243
rect 20898 13240 20904 13252
rect 20859 13212 20904 13240
rect 19613 13203 19671 13209
rect 15289 13175 15347 13181
rect 15289 13141 15301 13175
rect 15335 13172 15347 13175
rect 15838 13172 15844 13184
rect 15335 13144 15844 13172
rect 15335 13141 15347 13144
rect 15289 13135 15347 13141
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 17218 13172 17224 13184
rect 17179 13144 17224 13172
rect 17218 13132 17224 13144
rect 17276 13132 17282 13184
rect 19242 13132 19248 13184
rect 19300 13172 19306 13184
rect 19628 13172 19656 13203
rect 20898 13200 20904 13212
rect 20956 13200 20962 13252
rect 23198 13240 23204 13252
rect 23159 13212 23204 13240
rect 23198 13200 23204 13212
rect 23256 13200 23262 13252
rect 25682 13240 25688 13252
rect 25643 13212 25688 13240
rect 25682 13200 25688 13212
rect 25740 13200 25746 13252
rect 25777 13243 25835 13249
rect 25777 13209 25789 13243
rect 25823 13240 25835 13243
rect 25958 13240 25964 13252
rect 25823 13212 25964 13240
rect 25823 13209 25835 13212
rect 25777 13203 25835 13209
rect 25958 13200 25964 13212
rect 26016 13200 26022 13252
rect 26605 13243 26663 13249
rect 26605 13209 26617 13243
rect 26651 13209 26663 13243
rect 26605 13203 26663 13209
rect 26697 13243 26755 13249
rect 26697 13209 26709 13243
rect 26743 13209 26755 13243
rect 26697 13203 26755 13209
rect 19300 13144 19656 13172
rect 19300 13132 19306 13144
rect 21174 13132 21180 13184
rect 21232 13172 21238 13184
rect 23937 13175 23995 13181
rect 23937 13172 23949 13175
rect 21232 13144 23949 13172
rect 21232 13132 21238 13144
rect 23937 13141 23949 13144
rect 23983 13141 23995 13175
rect 23937 13135 23995 13141
rect 24762 13132 24768 13184
rect 24820 13172 24826 13184
rect 25866 13172 25872 13184
rect 24820 13144 25872 13172
rect 24820 13132 24826 13144
rect 25866 13132 25872 13144
rect 25924 13172 25930 13184
rect 26620 13172 26648 13203
rect 25924 13144 26648 13172
rect 26712 13172 26740 13203
rect 27522 13200 27528 13252
rect 27580 13240 27586 13252
rect 27617 13243 27675 13249
rect 27617 13240 27629 13243
rect 27580 13212 27629 13240
rect 27580 13200 27586 13212
rect 27617 13209 27629 13212
rect 27663 13209 27675 13243
rect 27724 13240 27752 13280
rect 28169 13243 28227 13249
rect 28169 13240 28181 13243
rect 27724 13212 28181 13240
rect 27617 13203 27675 13209
rect 28169 13209 28181 13212
rect 28215 13209 28227 13243
rect 28169 13203 28227 13209
rect 28261 13243 28319 13249
rect 28261 13209 28273 13243
rect 28307 13240 28319 13243
rect 29104 13240 29132 13348
rect 32953 13345 32965 13348
rect 32999 13345 33011 13379
rect 32953 13339 33011 13345
rect 30466 13268 30472 13320
rect 30524 13308 30530 13320
rect 30524 13280 30569 13308
rect 30524 13268 30530 13280
rect 31018 13268 31024 13320
rect 31076 13308 31082 13320
rect 31113 13311 31171 13317
rect 31113 13308 31125 13311
rect 31076 13280 31125 13308
rect 31076 13268 31082 13280
rect 31113 13277 31125 13280
rect 31159 13277 31171 13311
rect 31113 13271 31171 13277
rect 31757 13311 31815 13317
rect 31757 13277 31769 13311
rect 31803 13308 31815 13311
rect 32122 13308 32128 13320
rect 31803 13280 32128 13308
rect 31803 13277 31815 13280
rect 31757 13271 31815 13277
rect 32122 13268 32128 13280
rect 32180 13268 32186 13320
rect 32217 13311 32275 13317
rect 32217 13277 32229 13311
rect 32263 13308 32275 13311
rect 32858 13308 32864 13320
rect 32263 13280 32444 13308
rect 32819 13280 32864 13308
rect 32263 13277 32275 13280
rect 32217 13271 32275 13277
rect 28307 13212 29132 13240
rect 28307 13209 28319 13212
rect 28261 13203 28319 13209
rect 29178 13200 29184 13252
rect 29236 13240 29242 13252
rect 29236 13212 29281 13240
rect 29236 13200 29242 13212
rect 29638 13200 29644 13252
rect 29696 13240 29702 13252
rect 29825 13243 29883 13249
rect 29825 13240 29837 13243
rect 29696 13212 29837 13240
rect 29696 13200 29702 13212
rect 29825 13209 29837 13212
rect 29871 13209 29883 13243
rect 29825 13203 29883 13209
rect 29917 13243 29975 13249
rect 29917 13209 29929 13243
rect 29963 13240 29975 13243
rect 30282 13240 30288 13252
rect 29963 13212 30288 13240
rect 29963 13209 29975 13212
rect 29917 13203 29975 13209
rect 30282 13200 30288 13212
rect 30340 13200 30346 13252
rect 32309 13243 32367 13249
rect 32309 13240 32321 13243
rect 30576 13212 32321 13240
rect 30576 13172 30604 13212
rect 32309 13209 32321 13212
rect 32355 13209 32367 13243
rect 32309 13203 32367 13209
rect 26712 13144 30604 13172
rect 25924 13132 25930 13144
rect 31386 13132 31392 13184
rect 31444 13172 31450 13184
rect 32416 13172 32444 13280
rect 32858 13268 32864 13280
rect 32916 13268 32922 13320
rect 31444 13144 32444 13172
rect 31444 13132 31450 13144
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 13354 12968 13360 12980
rect 13315 12940 13360 12968
rect 13354 12928 13360 12940
rect 13412 12928 13418 12980
rect 14458 12968 14464 12980
rect 14371 12940 14464 12968
rect 14458 12928 14464 12940
rect 14516 12968 14522 12980
rect 17310 12968 17316 12980
rect 14516 12940 17316 12968
rect 14516 12928 14522 12940
rect 17310 12928 17316 12940
rect 17368 12928 17374 12980
rect 17862 12968 17868 12980
rect 17512 12940 17868 12968
rect 12805 12903 12863 12909
rect 12805 12869 12817 12903
rect 12851 12900 12863 12903
rect 15654 12900 15660 12912
rect 12851 12872 15660 12900
rect 12851 12869 12863 12872
rect 12805 12863 12863 12869
rect 15654 12860 15660 12872
rect 15712 12860 15718 12912
rect 15749 12903 15807 12909
rect 15749 12869 15761 12903
rect 15795 12900 15807 12903
rect 15838 12900 15844 12912
rect 15795 12872 15844 12900
rect 15795 12869 15807 12872
rect 15749 12863 15807 12869
rect 15838 12860 15844 12872
rect 15896 12860 15902 12912
rect 16022 12860 16028 12912
rect 16080 12900 16086 12912
rect 16301 12903 16359 12909
rect 16301 12900 16313 12903
rect 16080 12872 16313 12900
rect 16080 12860 16086 12872
rect 16301 12869 16313 12872
rect 16347 12869 16359 12903
rect 17512 12900 17540 12940
rect 17862 12928 17868 12940
rect 17920 12928 17926 12980
rect 22738 12968 22744 12980
rect 20916 12940 22744 12968
rect 16301 12863 16359 12869
rect 17144 12872 17540 12900
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12832 1915 12835
rect 4062 12832 4068 12844
rect 1903 12804 4068 12832
rect 1903 12801 1915 12804
rect 1857 12795 1915 12801
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 14918 12832 14924 12844
rect 14879 12804 14924 12832
rect 14918 12792 14924 12804
rect 14976 12792 14982 12844
rect 17144 12841 17172 12872
rect 17586 12860 17592 12912
rect 17644 12900 17650 12912
rect 17957 12903 18015 12909
rect 17957 12900 17969 12903
rect 17644 12872 17969 12900
rect 17644 12860 17650 12872
rect 17957 12869 17969 12872
rect 18003 12869 18015 12903
rect 19153 12903 19211 12909
rect 19153 12900 19165 12903
rect 17957 12863 18015 12869
rect 18524 12872 19165 12900
rect 17129 12835 17187 12841
rect 17129 12832 17141 12835
rect 16960 12804 17141 12832
rect 16960 12764 16988 12804
rect 17129 12801 17141 12804
rect 17175 12801 17187 12835
rect 17129 12795 17187 12801
rect 15672 12752 15884 12764
rect 16132 12752 16988 12764
rect 15672 12736 16988 12752
rect 13909 12699 13967 12705
rect 13909 12665 13921 12699
rect 13955 12696 13967 12699
rect 15672 12696 15700 12736
rect 15856 12724 16160 12736
rect 17034 12724 17040 12776
rect 17092 12764 17098 12776
rect 17310 12764 17316 12776
rect 17092 12736 17316 12764
rect 17092 12724 17098 12736
rect 17310 12724 17316 12736
rect 17368 12724 17374 12776
rect 17862 12764 17868 12776
rect 17823 12736 17868 12764
rect 17862 12724 17868 12736
rect 17920 12724 17926 12776
rect 18524 12764 18552 12872
rect 19153 12869 19165 12872
rect 19199 12869 19211 12903
rect 19153 12863 19211 12869
rect 19334 12860 19340 12912
rect 19392 12900 19398 12912
rect 20916 12909 20944 12940
rect 22738 12928 22744 12940
rect 22796 12928 22802 12980
rect 23198 12928 23204 12980
rect 23256 12968 23262 12980
rect 24857 12971 24915 12977
rect 24857 12968 24869 12971
rect 23256 12940 24869 12968
rect 23256 12928 23262 12940
rect 24857 12937 24869 12940
rect 24903 12937 24915 12971
rect 30101 12971 30159 12977
rect 30101 12968 30113 12971
rect 24857 12931 24915 12937
rect 26067 12940 30113 12968
rect 20809 12903 20867 12909
rect 20809 12900 20821 12903
rect 19392 12872 20821 12900
rect 19392 12860 19398 12872
rect 20809 12869 20821 12872
rect 20855 12869 20867 12903
rect 20809 12863 20867 12869
rect 20901 12903 20959 12909
rect 20901 12869 20913 12903
rect 20947 12869 20959 12903
rect 21450 12900 21456 12912
rect 21411 12872 21456 12900
rect 20901 12863 20959 12869
rect 21450 12860 21456 12872
rect 21508 12860 21514 12912
rect 22189 12903 22247 12909
rect 22189 12900 22201 12903
rect 21560 12872 22201 12900
rect 19058 12764 19064 12776
rect 17972 12736 18552 12764
rect 19019 12736 19064 12764
rect 13955 12668 15700 12696
rect 13955 12665 13967 12668
rect 13909 12659 13967 12665
rect 15746 12656 15752 12708
rect 15804 12696 15810 12708
rect 17972 12696 18000 12736
rect 19058 12724 19064 12736
rect 19116 12724 19122 12776
rect 20073 12767 20131 12773
rect 20073 12733 20085 12767
rect 20119 12764 20131 12767
rect 20162 12764 20168 12776
rect 20119 12736 20168 12764
rect 20119 12733 20131 12736
rect 20073 12727 20131 12733
rect 20162 12724 20168 12736
rect 20220 12764 20226 12776
rect 20530 12764 20536 12776
rect 20220 12736 20536 12764
rect 20220 12724 20226 12736
rect 20530 12724 20536 12736
rect 20588 12724 20594 12776
rect 15804 12668 18000 12696
rect 18417 12699 18475 12705
rect 15804 12656 15810 12668
rect 18417 12665 18429 12699
rect 18463 12696 18475 12699
rect 18874 12696 18880 12708
rect 18463 12668 18880 12696
rect 18463 12665 18475 12668
rect 18417 12659 18475 12665
rect 18874 12656 18880 12668
rect 18932 12696 18938 12708
rect 18932 12668 20208 12696
rect 18932 12656 18938 12668
rect 1670 12628 1676 12640
rect 1631 12600 1676 12628
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 15013 12631 15071 12637
rect 15013 12597 15025 12631
rect 15059 12628 15071 12631
rect 16482 12628 16488 12640
rect 15059 12600 16488 12628
rect 15059 12597 15071 12600
rect 15013 12591 15071 12597
rect 16482 12588 16488 12600
rect 16540 12588 16546 12640
rect 17221 12631 17279 12637
rect 17221 12597 17233 12631
rect 17267 12628 17279 12631
rect 20070 12628 20076 12640
rect 17267 12600 20076 12628
rect 17267 12597 17279 12600
rect 17221 12591 17279 12597
rect 20070 12588 20076 12600
rect 20128 12588 20134 12640
rect 20180 12628 20208 12668
rect 20254 12656 20260 12708
rect 20312 12696 20318 12708
rect 21560 12696 21588 12872
rect 22189 12869 22201 12872
rect 22235 12869 22247 12903
rect 22189 12863 22247 12869
rect 23474 12860 23480 12912
rect 23532 12900 23538 12912
rect 23661 12903 23719 12909
rect 23661 12900 23673 12903
rect 23532 12872 23673 12900
rect 23532 12860 23538 12872
rect 23661 12869 23673 12872
rect 23707 12869 23719 12903
rect 23661 12863 23719 12869
rect 23753 12903 23811 12909
rect 23753 12869 23765 12903
rect 23799 12900 23811 12903
rect 25314 12900 25320 12912
rect 23799 12872 25320 12900
rect 23799 12869 23811 12872
rect 23753 12863 23811 12869
rect 25314 12860 25320 12872
rect 25372 12860 25378 12912
rect 25774 12860 25780 12912
rect 25832 12900 25838 12912
rect 26067 12909 26095 12940
rect 30101 12937 30113 12940
rect 30147 12937 30159 12971
rect 30101 12931 30159 12937
rect 30282 12928 30288 12980
rect 30340 12968 30346 12980
rect 32401 12971 32459 12977
rect 32401 12968 32413 12971
rect 30340 12940 32413 12968
rect 30340 12928 30346 12940
rect 32401 12937 32413 12940
rect 32447 12937 32459 12971
rect 32401 12931 32459 12937
rect 25961 12903 26019 12909
rect 25961 12900 25973 12903
rect 25832 12872 25973 12900
rect 25832 12860 25838 12872
rect 25961 12869 25973 12872
rect 26007 12869 26019 12903
rect 25961 12863 26019 12869
rect 26053 12903 26111 12909
rect 26053 12869 26065 12903
rect 26099 12869 26111 12903
rect 26053 12863 26111 12869
rect 26970 12860 26976 12912
rect 27028 12900 27034 12912
rect 27709 12903 27767 12909
rect 27709 12900 27721 12903
rect 27028 12872 27721 12900
rect 27028 12860 27034 12872
rect 27709 12869 27721 12872
rect 27755 12869 27767 12903
rect 27709 12863 27767 12869
rect 27801 12903 27859 12909
rect 27801 12869 27813 12903
rect 27847 12900 27859 12903
rect 29822 12900 29828 12912
rect 27847 12872 29828 12900
rect 27847 12869 27859 12872
rect 27801 12863 27859 12869
rect 29822 12860 29828 12872
rect 29880 12860 29886 12912
rect 32950 12900 32956 12912
rect 32911 12872 32956 12900
rect 32950 12860 32956 12872
rect 33008 12860 33014 12912
rect 24949 12835 25007 12841
rect 24949 12801 24961 12835
rect 24995 12801 25007 12835
rect 24949 12795 25007 12801
rect 28353 12835 28411 12841
rect 28353 12801 28365 12835
rect 28399 12832 28411 12835
rect 28902 12832 28908 12844
rect 28399 12804 28908 12832
rect 28399 12801 28411 12804
rect 28353 12795 28411 12801
rect 22097 12767 22155 12773
rect 22097 12733 22109 12767
rect 22143 12733 22155 12767
rect 23014 12764 23020 12776
rect 22975 12736 23020 12764
rect 22097 12727 22155 12733
rect 20312 12668 21588 12696
rect 20312 12656 20318 12668
rect 22112 12628 22140 12727
rect 23014 12724 23020 12736
rect 23072 12724 23078 12776
rect 23382 12724 23388 12776
rect 23440 12764 23446 12776
rect 23937 12767 23995 12773
rect 23937 12764 23949 12767
rect 23440 12736 23949 12764
rect 23440 12724 23446 12736
rect 23937 12733 23949 12736
rect 23983 12764 23995 12767
rect 24762 12764 24768 12776
rect 23983 12736 24768 12764
rect 23983 12733 23995 12736
rect 23937 12727 23995 12733
rect 24762 12724 24768 12736
rect 24820 12724 24826 12776
rect 24964 12696 24992 12795
rect 28902 12792 28908 12804
rect 28960 12792 28966 12844
rect 28994 12792 29000 12844
rect 29052 12832 29058 12844
rect 29052 12804 29097 12832
rect 29052 12792 29058 12804
rect 29638 12792 29644 12844
rect 29696 12830 29702 12844
rect 30929 12835 30987 12841
rect 29696 12802 29739 12830
rect 29696 12792 29702 12802
rect 30929 12801 30941 12835
rect 30975 12801 30987 12835
rect 31570 12832 31576 12844
rect 31531 12804 31576 12832
rect 30929 12795 30987 12801
rect 25777 12767 25835 12773
rect 25777 12733 25789 12767
rect 25823 12764 25835 12767
rect 25866 12764 25872 12776
rect 25823 12736 25872 12764
rect 25823 12733 25835 12736
rect 25777 12727 25835 12733
rect 25866 12724 25872 12736
rect 25924 12724 25930 12776
rect 26050 12724 26056 12776
rect 26108 12764 26114 12776
rect 29012 12764 29040 12792
rect 26108 12736 29040 12764
rect 26108 12724 26114 12736
rect 29178 12724 29184 12776
rect 29236 12764 29242 12776
rect 29549 12767 29607 12773
rect 29549 12764 29561 12767
rect 29236 12736 29561 12764
rect 29236 12724 29242 12736
rect 29549 12733 29561 12736
rect 29595 12733 29607 12767
rect 29549 12727 29607 12733
rect 30650 12724 30656 12776
rect 30708 12764 30714 12776
rect 30837 12767 30895 12773
rect 30837 12764 30849 12767
rect 30708 12736 30849 12764
rect 30708 12724 30714 12736
rect 30837 12733 30849 12736
rect 30883 12733 30895 12767
rect 30944 12764 30972 12795
rect 31570 12792 31576 12804
rect 31628 12792 31634 12844
rect 32493 12835 32551 12841
rect 32493 12801 32505 12835
rect 32539 12832 32551 12835
rect 33594 12832 33600 12844
rect 32539 12804 33600 12832
rect 32539 12801 32551 12804
rect 32493 12795 32551 12801
rect 33594 12792 33600 12804
rect 33652 12792 33658 12844
rect 31846 12764 31852 12776
rect 30944 12736 31852 12764
rect 30837 12727 30895 12733
rect 31846 12724 31852 12736
rect 31904 12724 31910 12776
rect 27890 12696 27896 12708
rect 24964 12668 27896 12696
rect 27890 12656 27896 12668
rect 27948 12656 27954 12708
rect 28442 12656 28448 12708
rect 28500 12696 28506 12708
rect 28500 12668 29592 12696
rect 28500 12656 28506 12668
rect 20180 12600 22140 12628
rect 25590 12588 25596 12640
rect 25648 12628 25654 12640
rect 26050 12628 26056 12640
rect 25648 12600 26056 12628
rect 25648 12588 25654 12600
rect 26050 12588 26056 12600
rect 26108 12588 26114 12640
rect 26326 12588 26332 12640
rect 26384 12628 26390 12640
rect 28905 12631 28963 12637
rect 28905 12628 28917 12631
rect 26384 12600 28917 12628
rect 26384 12588 26390 12600
rect 28905 12597 28917 12600
rect 28951 12597 28963 12631
rect 29564 12628 29592 12668
rect 31481 12631 31539 12637
rect 31481 12628 31493 12631
rect 29564 12600 31493 12628
rect 28905 12591 28963 12597
rect 31481 12597 31493 12600
rect 31527 12597 31539 12631
rect 31481 12591 31539 12597
rect 37642 12588 37648 12640
rect 37700 12628 37706 12640
rect 37921 12631 37979 12637
rect 37921 12628 37933 12631
rect 37700 12600 37933 12628
rect 37700 12588 37706 12600
rect 37921 12597 37933 12600
rect 37967 12597 37979 12631
rect 37921 12591 37979 12597
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 13722 12384 13728 12436
rect 13780 12424 13786 12436
rect 14274 12424 14280 12436
rect 13780 12396 14280 12424
rect 13780 12384 13786 12396
rect 14274 12384 14280 12396
rect 14332 12424 14338 12436
rect 14332 12396 18092 12424
rect 14332 12384 14338 12396
rect 14553 12359 14611 12365
rect 14553 12325 14565 12359
rect 14599 12356 14611 12359
rect 17862 12356 17868 12368
rect 14599 12328 17868 12356
rect 14599 12325 14611 12328
rect 14553 12319 14611 12325
rect 17862 12316 17868 12328
rect 17920 12356 17926 12368
rect 18064 12356 18092 12396
rect 18138 12384 18144 12436
rect 18196 12424 18202 12436
rect 19150 12424 19156 12436
rect 18196 12396 19156 12424
rect 18196 12384 18202 12396
rect 19150 12384 19156 12396
rect 19208 12384 19214 12436
rect 24118 12424 24124 12436
rect 20456 12396 24124 12424
rect 19334 12356 19340 12368
rect 17920 12328 18000 12356
rect 18064 12328 19340 12356
rect 17920 12316 17926 12328
rect 1854 12248 1860 12300
rect 1912 12288 1918 12300
rect 8294 12288 8300 12300
rect 1912 12260 8300 12288
rect 1912 12248 1918 12260
rect 8294 12248 8300 12260
rect 8352 12248 8358 12300
rect 12621 12291 12679 12297
rect 12621 12257 12633 12291
rect 12667 12288 12679 12291
rect 16850 12288 16856 12300
rect 12667 12260 15148 12288
rect 12667 12257 12679 12260
rect 12621 12251 12679 12257
rect 12069 12223 12127 12229
rect 12069 12189 12081 12223
rect 12115 12220 12127 12223
rect 14458 12220 14464 12232
rect 12115 12192 14464 12220
rect 12115 12189 12127 12192
rect 12069 12183 12127 12189
rect 14458 12180 14464 12192
rect 14516 12180 14522 12232
rect 15120 12229 15148 12260
rect 15948 12260 16856 12288
rect 15105 12223 15163 12229
rect 15105 12189 15117 12223
rect 15151 12220 15163 12223
rect 15838 12220 15844 12232
rect 15151 12192 15844 12220
rect 15151 12189 15163 12192
rect 15105 12183 15163 12189
rect 15838 12180 15844 12192
rect 15896 12180 15902 12232
rect 15948 12229 15976 12260
rect 16850 12248 16856 12260
rect 16908 12248 16914 12300
rect 17037 12291 17095 12297
rect 17037 12257 17049 12291
rect 17083 12288 17095 12291
rect 17586 12288 17592 12300
rect 17083 12260 17592 12288
rect 17083 12257 17095 12260
rect 17037 12251 17095 12257
rect 17586 12248 17592 12260
rect 17644 12248 17650 12300
rect 17972 12288 18000 12328
rect 19334 12316 19340 12328
rect 19392 12316 19398 12368
rect 18141 12291 18199 12297
rect 18141 12288 18153 12291
rect 17972 12260 18153 12288
rect 18141 12257 18153 12260
rect 18187 12257 18199 12291
rect 18141 12251 18199 12257
rect 18230 12248 18236 12300
rect 18288 12288 18294 12300
rect 20456 12297 20484 12396
rect 24118 12384 24124 12396
rect 24176 12384 24182 12436
rect 24486 12384 24492 12436
rect 24544 12424 24550 12436
rect 26326 12424 26332 12436
rect 24544 12396 26332 12424
rect 24544 12384 24550 12396
rect 26326 12384 26332 12396
rect 26384 12384 26390 12436
rect 26418 12384 26424 12436
rect 26476 12424 26482 12436
rect 28442 12424 28448 12436
rect 26476 12396 28448 12424
rect 26476 12384 26482 12396
rect 28442 12384 28448 12396
rect 28500 12384 28506 12436
rect 28534 12384 28540 12436
rect 28592 12424 28598 12436
rect 29825 12427 29883 12433
rect 29825 12424 29837 12427
rect 28592 12396 29837 12424
rect 28592 12384 28598 12396
rect 29825 12393 29837 12396
rect 29871 12393 29883 12427
rect 29825 12387 29883 12393
rect 31754 12384 31760 12436
rect 31812 12424 31818 12436
rect 31812 12396 31857 12424
rect 31812 12384 31818 12396
rect 21910 12316 21916 12368
rect 21968 12356 21974 12368
rect 21968 12328 22048 12356
rect 21968 12316 21974 12328
rect 20441 12291 20499 12297
rect 18288 12260 18828 12288
rect 18288 12248 18294 12260
rect 15933 12223 15991 12229
rect 15933 12189 15945 12223
rect 15979 12189 15991 12223
rect 15933 12183 15991 12189
rect 16022 12180 16028 12232
rect 16080 12220 16086 12232
rect 18800 12229 18828 12260
rect 20441 12257 20453 12291
rect 20487 12257 20499 12291
rect 20441 12251 20499 12257
rect 20714 12248 20720 12300
rect 20772 12288 20778 12300
rect 22020 12297 22048 12328
rect 22922 12316 22928 12368
rect 22980 12356 22986 12368
rect 27157 12359 27215 12365
rect 27157 12356 27169 12359
rect 22980 12328 27169 12356
rect 22980 12316 22986 12328
rect 27157 12325 27169 12328
rect 27203 12325 27215 12359
rect 27157 12319 27215 12325
rect 27430 12316 27436 12368
rect 27488 12356 27494 12368
rect 31113 12359 31171 12365
rect 31113 12356 31125 12359
rect 27488 12328 31125 12356
rect 27488 12316 27494 12328
rect 21177 12291 21235 12297
rect 21177 12288 21189 12291
rect 20772 12260 21189 12288
rect 20772 12248 20778 12260
rect 21177 12257 21189 12260
rect 21223 12257 21235 12291
rect 21177 12251 21235 12257
rect 22005 12291 22063 12297
rect 22005 12257 22017 12291
rect 22051 12257 22063 12291
rect 23106 12288 23112 12300
rect 23067 12260 23112 12288
rect 22005 12251 22063 12257
rect 23106 12248 23112 12260
rect 23164 12248 23170 12300
rect 23566 12248 23572 12300
rect 23624 12288 23630 12300
rect 23753 12291 23811 12297
rect 23753 12288 23765 12291
rect 23624 12260 23765 12288
rect 23624 12248 23630 12260
rect 23753 12257 23765 12260
rect 23799 12288 23811 12291
rect 24578 12288 24584 12300
rect 23799 12260 24584 12288
rect 23799 12257 23811 12260
rect 23753 12251 23811 12257
rect 24578 12248 24584 12260
rect 24636 12248 24642 12300
rect 25130 12248 25136 12300
rect 25188 12288 25194 12300
rect 25225 12291 25283 12297
rect 25225 12288 25237 12291
rect 25188 12260 25237 12288
rect 25188 12248 25194 12260
rect 25225 12257 25237 12260
rect 25271 12257 25283 12291
rect 25225 12251 25283 12257
rect 25866 12248 25872 12300
rect 25924 12288 25930 12300
rect 26142 12288 26148 12300
rect 25924 12260 26148 12288
rect 25924 12248 25930 12260
rect 26142 12248 26148 12260
rect 26200 12248 26206 12300
rect 27709 12291 27767 12297
rect 27709 12257 27721 12291
rect 27755 12288 27767 12291
rect 28994 12288 29000 12300
rect 27755 12260 29000 12288
rect 27755 12257 27767 12260
rect 27709 12251 27767 12257
rect 28994 12248 29000 12260
rect 29052 12248 29058 12300
rect 29104 12297 29132 12328
rect 31113 12325 31125 12328
rect 31159 12325 31171 12359
rect 31113 12319 31171 12325
rect 31570 12316 31576 12368
rect 31628 12356 31634 12368
rect 32953 12359 33011 12365
rect 32953 12356 32965 12359
rect 31628 12328 32965 12356
rect 31628 12316 31634 12328
rect 32953 12325 32965 12328
rect 32999 12325 33011 12359
rect 32953 12319 33011 12325
rect 29089 12291 29147 12297
rect 29089 12257 29101 12291
rect 29135 12257 29147 12291
rect 32398 12288 32404 12300
rect 32359 12260 32404 12288
rect 29089 12251 29147 12257
rect 32398 12248 32404 12260
rect 32456 12248 32462 12300
rect 16393 12223 16451 12229
rect 16393 12220 16405 12223
rect 16080 12192 16405 12220
rect 16080 12180 16086 12192
rect 16393 12189 16405 12192
rect 16439 12189 16451 12223
rect 16393 12183 16451 12189
rect 18785 12223 18843 12229
rect 18785 12189 18797 12223
rect 18831 12220 18843 12223
rect 19797 12223 19855 12229
rect 19797 12220 19809 12223
rect 18831 12192 19809 12220
rect 18831 12189 18843 12192
rect 18785 12183 18843 12189
rect 19797 12189 19809 12192
rect 19843 12189 19855 12223
rect 29914 12220 29920 12232
rect 29875 12192 29920 12220
rect 19797 12183 19855 12189
rect 29914 12180 29920 12192
rect 29972 12180 29978 12232
rect 30374 12220 30380 12232
rect 30335 12192 30380 12220
rect 30374 12180 30380 12192
rect 30432 12180 30438 12232
rect 31205 12223 31263 12229
rect 31205 12220 31217 12223
rect 30576 12192 31217 12220
rect 13725 12155 13783 12161
rect 13725 12121 13737 12155
rect 13771 12152 13783 12155
rect 16298 12152 16304 12164
rect 13771 12124 16304 12152
rect 13771 12121 13783 12124
rect 13725 12115 13783 12121
rect 16298 12112 16304 12124
rect 16356 12112 16362 12164
rect 16942 12152 16948 12164
rect 16903 12124 16948 12152
rect 16942 12112 16948 12124
rect 17000 12112 17006 12164
rect 18233 12155 18291 12161
rect 18233 12121 18245 12155
rect 18279 12152 18291 12155
rect 18506 12152 18512 12164
rect 18279 12124 18512 12152
rect 18279 12121 18291 12124
rect 18233 12115 18291 12121
rect 18506 12112 18512 12124
rect 18564 12112 18570 12164
rect 18874 12112 18880 12164
rect 18932 12152 18938 12164
rect 20349 12155 20407 12161
rect 20349 12152 20361 12155
rect 18932 12124 20361 12152
rect 18932 12112 18938 12124
rect 20349 12121 20361 12124
rect 20395 12121 20407 12155
rect 20349 12115 20407 12121
rect 21174 12112 21180 12164
rect 21232 12152 21238 12164
rect 21269 12155 21327 12161
rect 21269 12152 21281 12155
rect 21232 12124 21281 12152
rect 21232 12112 21238 12124
rect 21269 12121 21281 12124
rect 21315 12121 21327 12155
rect 21269 12115 21327 12121
rect 23661 12155 23719 12161
rect 23661 12121 23673 12155
rect 23707 12152 23719 12155
rect 23750 12152 23756 12164
rect 23707 12124 23756 12152
rect 23707 12121 23719 12124
rect 23661 12115 23719 12121
rect 23750 12112 23756 12124
rect 23808 12112 23814 12164
rect 24578 12152 24584 12164
rect 24539 12124 24584 12152
rect 24578 12112 24584 12124
rect 24636 12112 24642 12164
rect 25133 12155 25191 12161
rect 25133 12121 25145 12155
rect 25179 12121 25191 12155
rect 26418 12152 26424 12164
rect 26379 12124 26424 12152
rect 25133 12115 25191 12121
rect 13173 12087 13231 12093
rect 13173 12053 13185 12087
rect 13219 12084 13231 12087
rect 14918 12084 14924 12096
rect 13219 12056 14924 12084
rect 13219 12053 13231 12056
rect 13173 12047 13231 12053
rect 14918 12044 14924 12056
rect 14976 12044 14982 12096
rect 15194 12084 15200 12096
rect 15155 12056 15200 12084
rect 15194 12044 15200 12056
rect 15252 12044 15258 12096
rect 15841 12087 15899 12093
rect 15841 12053 15853 12087
rect 15887 12084 15899 12087
rect 19978 12084 19984 12096
rect 15887 12056 19984 12084
rect 15887 12053 15899 12056
rect 15841 12047 15899 12053
rect 19978 12044 19984 12056
rect 20036 12044 20042 12096
rect 20806 12044 20812 12096
rect 20864 12084 20870 12096
rect 23566 12084 23572 12096
rect 20864 12056 23572 12084
rect 20864 12044 20870 12056
rect 23566 12044 23572 12056
rect 23624 12044 23630 12096
rect 25148 12084 25176 12115
rect 26418 12112 26424 12124
rect 26476 12112 26482 12164
rect 26513 12155 26571 12161
rect 26513 12121 26525 12155
rect 26559 12152 26571 12155
rect 27522 12152 27528 12164
rect 26559 12124 27528 12152
rect 26559 12121 26571 12124
rect 26513 12115 26571 12121
rect 27522 12112 27528 12124
rect 27580 12112 27586 12164
rect 27617 12155 27675 12161
rect 27617 12121 27629 12155
rect 27663 12152 27675 12155
rect 28350 12152 28356 12164
rect 27663 12124 28356 12152
rect 27663 12121 27675 12124
rect 27617 12115 27675 12121
rect 28350 12112 28356 12124
rect 28408 12112 28414 12164
rect 28442 12112 28448 12164
rect 28500 12152 28506 12164
rect 28500 12124 28545 12152
rect 28500 12112 28506 12124
rect 28994 12112 29000 12164
rect 29052 12152 29058 12164
rect 30466 12152 30472 12164
rect 29052 12124 29097 12152
rect 30427 12124 30472 12152
rect 29052 12112 29058 12124
rect 30466 12112 30472 12124
rect 30524 12112 30530 12164
rect 29086 12084 29092 12096
rect 25148 12056 29092 12084
rect 29086 12044 29092 12056
rect 29144 12044 29150 12096
rect 30098 12044 30104 12096
rect 30156 12084 30162 12096
rect 30576 12084 30604 12192
rect 31205 12189 31217 12192
rect 31251 12189 31263 12223
rect 31662 12220 31668 12232
rect 31623 12192 31668 12220
rect 31205 12183 31263 12189
rect 31220 12152 31248 12183
rect 31662 12180 31668 12192
rect 31720 12180 31726 12232
rect 32493 12223 32551 12229
rect 32493 12189 32505 12223
rect 32539 12220 32551 12223
rect 34422 12220 34428 12232
rect 32539 12192 34428 12220
rect 32539 12189 32551 12192
rect 32493 12183 32551 12189
rect 34422 12180 34428 12192
rect 34480 12180 34486 12232
rect 37550 12152 37556 12164
rect 31220 12124 37556 12152
rect 37550 12112 37556 12124
rect 37608 12112 37614 12164
rect 30156 12056 30604 12084
rect 37461 12087 37519 12093
rect 30156 12044 30162 12056
rect 37461 12053 37473 12087
rect 37507 12084 37519 12087
rect 37826 12084 37832 12096
rect 37507 12056 37832 12084
rect 37507 12053 37519 12056
rect 37461 12047 37519 12053
rect 37826 12044 37832 12056
rect 37884 12044 37890 12096
rect 37918 12044 37924 12096
rect 37976 12084 37982 12096
rect 37976 12056 38021 12084
rect 37976 12044 37982 12056
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 6546 11880 6552 11892
rect 6507 11852 6552 11880
rect 6546 11840 6552 11852
rect 6604 11880 6610 11892
rect 6604 11852 6914 11880
rect 6604 11840 6610 11852
rect 5905 11747 5963 11753
rect 5905 11713 5917 11747
rect 5951 11744 5963 11747
rect 6886 11744 6914 11852
rect 15194 11840 15200 11892
rect 15252 11880 15258 11892
rect 19889 11883 19947 11889
rect 15252 11852 18644 11880
rect 15252 11840 15258 11852
rect 12897 11815 12955 11821
rect 12897 11781 12909 11815
rect 12943 11812 12955 11815
rect 15013 11815 15071 11821
rect 12943 11784 14320 11812
rect 12943 11781 12955 11784
rect 12897 11775 12955 11781
rect 14292 11756 14320 11784
rect 15013 11781 15025 11815
rect 15059 11812 15071 11815
rect 15746 11812 15752 11824
rect 15059 11784 15752 11812
rect 15059 11781 15071 11784
rect 15013 11775 15071 11781
rect 15746 11772 15752 11784
rect 15804 11772 15810 11824
rect 16117 11815 16175 11821
rect 16117 11781 16129 11815
rect 16163 11812 16175 11815
rect 17678 11812 17684 11824
rect 16163 11784 17172 11812
rect 17639 11784 17684 11812
rect 16163 11781 16175 11784
rect 16117 11775 16175 11781
rect 12345 11747 12403 11753
rect 12345 11744 12357 11747
rect 5951 11716 12357 11744
rect 5951 11713 5963 11716
rect 5905 11707 5963 11713
rect 12345 11713 12357 11716
rect 12391 11744 12403 11747
rect 13357 11747 13415 11753
rect 13357 11744 13369 11747
rect 12391 11716 13369 11744
rect 12391 11713 12403 11716
rect 12345 11707 12403 11713
rect 13357 11713 13369 11716
rect 13403 11713 13415 11747
rect 14274 11744 14280 11756
rect 14235 11716 14280 11744
rect 13357 11707 13415 11713
rect 14274 11704 14280 11716
rect 14332 11704 14338 11756
rect 15105 11747 15163 11753
rect 15105 11713 15117 11747
rect 15151 11744 15163 11747
rect 15562 11744 15568 11756
rect 15151 11716 15568 11744
rect 15151 11713 15163 11716
rect 15105 11707 15163 11713
rect 15562 11704 15568 11716
rect 15620 11704 15626 11756
rect 13449 11679 13507 11685
rect 13449 11645 13461 11679
rect 13495 11676 13507 11679
rect 16209 11679 16267 11685
rect 16209 11676 16221 11679
rect 13495 11648 16221 11676
rect 13495 11645 13507 11648
rect 13449 11639 13507 11645
rect 16209 11645 16221 11648
rect 16255 11676 16267 11679
rect 16390 11676 16396 11688
rect 16255 11648 16396 11676
rect 16255 11645 16267 11648
rect 16209 11639 16267 11645
rect 16390 11636 16396 11648
rect 16448 11636 16454 11688
rect 17144 11676 17172 11784
rect 17678 11772 17684 11784
rect 17736 11772 17742 11824
rect 17773 11815 17831 11821
rect 17773 11781 17785 11815
rect 17819 11812 17831 11815
rect 17954 11812 17960 11824
rect 17819 11784 17960 11812
rect 17819 11781 17831 11784
rect 17773 11775 17831 11781
rect 17954 11772 17960 11784
rect 18012 11772 18018 11824
rect 18616 11821 18644 11852
rect 19889 11849 19901 11883
rect 19935 11880 19947 11883
rect 20254 11880 20260 11892
rect 19935 11852 20260 11880
rect 19935 11849 19947 11852
rect 19889 11843 19947 11849
rect 20254 11840 20260 11852
rect 20312 11840 20318 11892
rect 22002 11840 22008 11892
rect 22060 11880 22066 11892
rect 22649 11883 22707 11889
rect 22060 11852 22232 11880
rect 22060 11840 22066 11852
rect 18601 11815 18659 11821
rect 18601 11781 18613 11815
rect 18647 11781 18659 11815
rect 18601 11775 18659 11781
rect 19153 11815 19211 11821
rect 19153 11781 19165 11815
rect 19199 11812 19211 11815
rect 20806 11812 20812 11824
rect 19199 11784 20812 11812
rect 19199 11781 19211 11784
rect 19153 11775 19211 11781
rect 20806 11772 20812 11784
rect 20864 11772 20870 11824
rect 20990 11812 20996 11824
rect 20951 11784 20996 11812
rect 20990 11772 20996 11784
rect 21048 11772 21054 11824
rect 21085 11815 21143 11821
rect 21085 11781 21097 11815
rect 21131 11812 21143 11815
rect 22094 11812 22100 11824
rect 21131 11784 22100 11812
rect 21131 11781 21143 11784
rect 21085 11775 21143 11781
rect 22094 11772 22100 11784
rect 22152 11772 22158 11824
rect 19794 11744 19800 11756
rect 19755 11716 19800 11744
rect 19794 11704 19800 11716
rect 19852 11704 19858 11756
rect 22204 11753 22232 11852
rect 22649 11849 22661 11883
rect 22695 11880 22707 11883
rect 23290 11880 23296 11892
rect 22695 11852 23296 11880
rect 22695 11849 22707 11852
rect 22649 11843 22707 11849
rect 23290 11840 23296 11852
rect 23348 11840 23354 11892
rect 24486 11880 24492 11892
rect 23676 11852 24492 11880
rect 23676 11821 23704 11852
rect 24486 11840 24492 11852
rect 24544 11840 24550 11892
rect 24596 11852 27200 11880
rect 23661 11815 23719 11821
rect 23661 11781 23673 11815
rect 23707 11781 23719 11815
rect 23661 11775 23719 11781
rect 23753 11815 23811 11821
rect 23753 11781 23765 11815
rect 23799 11812 23811 11815
rect 23934 11812 23940 11824
rect 23799 11784 23940 11812
rect 23799 11781 23811 11784
rect 23753 11775 23811 11781
rect 23934 11772 23940 11784
rect 23992 11772 23998 11824
rect 24302 11772 24308 11824
rect 24360 11812 24366 11824
rect 24596 11812 24624 11852
rect 24854 11812 24860 11824
rect 24360 11784 24624 11812
rect 24815 11784 24860 11812
rect 24360 11772 24366 11784
rect 24854 11772 24860 11784
rect 24912 11772 24918 11824
rect 24949 11815 25007 11821
rect 24949 11781 24961 11815
rect 24995 11812 25007 11815
rect 25130 11812 25136 11824
rect 24995 11784 25136 11812
rect 24995 11781 25007 11784
rect 24949 11775 25007 11781
rect 25130 11772 25136 11784
rect 25188 11772 25194 11824
rect 26234 11772 26240 11824
rect 26292 11812 26298 11824
rect 27172 11821 27200 11852
rect 28718 11840 28724 11892
rect 28776 11880 28782 11892
rect 29089 11883 29147 11889
rect 29089 11880 29101 11883
rect 28776 11852 29101 11880
rect 28776 11840 28782 11852
rect 29089 11849 29101 11852
rect 29135 11849 29147 11883
rect 30834 11880 30840 11892
rect 29089 11843 29147 11849
rect 29196 11852 30840 11880
rect 26329 11815 26387 11821
rect 26329 11812 26341 11815
rect 26292 11784 26341 11812
rect 26292 11772 26298 11784
rect 26329 11781 26341 11784
rect 26375 11781 26387 11815
rect 26329 11775 26387 11781
rect 27157 11815 27215 11821
rect 27157 11781 27169 11815
rect 27203 11781 27215 11815
rect 27157 11775 27215 11781
rect 27709 11815 27767 11821
rect 27709 11781 27721 11815
rect 27755 11812 27767 11815
rect 27755 11784 28994 11812
rect 27755 11781 27767 11784
rect 27709 11775 27767 11781
rect 22189 11747 22247 11753
rect 22189 11713 22201 11747
rect 22235 11713 22247 11747
rect 22189 11707 22247 11713
rect 28258 11704 28264 11756
rect 28316 11744 28322 11756
rect 28353 11747 28411 11753
rect 28353 11744 28365 11747
rect 28316 11716 28365 11744
rect 28316 11704 28322 11716
rect 28353 11713 28365 11716
rect 28399 11713 28411 11747
rect 28966 11744 28994 11784
rect 29086 11744 29092 11756
rect 28966 11716 29092 11744
rect 28353 11707 28411 11713
rect 29086 11704 29092 11716
rect 29144 11704 29150 11756
rect 29196 11753 29224 11852
rect 30834 11840 30840 11852
rect 30892 11880 30898 11892
rect 30892 11852 31156 11880
rect 30892 11840 30898 11852
rect 29730 11772 29736 11824
rect 29788 11812 29794 11824
rect 31021 11815 31079 11821
rect 31021 11812 31033 11815
rect 29788 11784 31033 11812
rect 29788 11772 29794 11784
rect 31021 11781 31033 11784
rect 31067 11781 31079 11815
rect 31021 11775 31079 11781
rect 29181 11747 29239 11753
rect 29181 11713 29193 11747
rect 29227 11713 29239 11747
rect 29822 11744 29828 11756
rect 29783 11716 29828 11744
rect 29181 11707 29239 11713
rect 29822 11704 29828 11716
rect 29880 11704 29886 11756
rect 30282 11704 30288 11756
rect 30340 11744 30346 11756
rect 31128 11753 31156 11852
rect 31202 11840 31208 11892
rect 31260 11880 31266 11892
rect 31665 11883 31723 11889
rect 31665 11880 31677 11883
rect 31260 11852 31677 11880
rect 31260 11840 31266 11852
rect 31665 11849 31677 11852
rect 31711 11849 31723 11883
rect 31665 11843 31723 11849
rect 30469 11747 30527 11753
rect 30469 11744 30481 11747
rect 30340 11716 30481 11744
rect 30340 11704 30346 11716
rect 30469 11713 30481 11716
rect 30515 11713 30527 11747
rect 30469 11707 30527 11713
rect 31113 11747 31171 11753
rect 31113 11713 31125 11747
rect 31159 11744 31171 11747
rect 31202 11744 31208 11756
rect 31159 11716 31208 11744
rect 31159 11713 31171 11716
rect 31113 11707 31171 11713
rect 17144 11648 17724 11676
rect 15654 11608 15660 11620
rect 15615 11580 15660 11608
rect 15654 11568 15660 11580
rect 15712 11568 15718 11620
rect 16022 11568 16028 11620
rect 16080 11608 16086 11620
rect 17221 11611 17279 11617
rect 17221 11608 17233 11611
rect 16080 11580 17233 11608
rect 16080 11568 16086 11580
rect 17221 11577 17233 11580
rect 17267 11577 17279 11611
rect 17696 11608 17724 11648
rect 17954 11636 17960 11688
rect 18012 11676 18018 11688
rect 18509 11679 18567 11685
rect 18509 11676 18521 11679
rect 18012 11648 18521 11676
rect 18012 11636 18018 11648
rect 18509 11645 18521 11648
rect 18555 11645 18567 11679
rect 18509 11639 18567 11645
rect 18598 11636 18604 11688
rect 18656 11676 18662 11688
rect 20441 11679 20499 11685
rect 20441 11676 20453 11679
rect 18656 11648 20453 11676
rect 18656 11636 18662 11648
rect 20441 11645 20453 11648
rect 20487 11645 20499 11679
rect 20441 11639 20499 11645
rect 21818 11636 21824 11688
rect 21876 11676 21882 11688
rect 22005 11679 22063 11685
rect 22005 11676 22017 11679
rect 21876 11648 22017 11676
rect 21876 11636 21882 11648
rect 22005 11645 22017 11648
rect 22051 11645 22063 11679
rect 22005 11639 22063 11645
rect 26421 11679 26479 11685
rect 26421 11645 26433 11679
rect 26467 11676 26479 11679
rect 27430 11676 27436 11688
rect 26467 11648 27436 11676
rect 26467 11645 26479 11648
rect 26421 11639 26479 11645
rect 27430 11636 27436 11648
rect 27488 11636 27494 11688
rect 27522 11636 27528 11688
rect 27580 11676 27586 11688
rect 27801 11679 27859 11685
rect 27801 11676 27813 11679
rect 27580 11648 27813 11676
rect 27580 11636 27586 11648
rect 27801 11645 27813 11648
rect 27847 11676 27859 11679
rect 30377 11679 30435 11685
rect 30377 11676 30389 11679
rect 27847 11648 30389 11676
rect 27847 11645 27859 11648
rect 27801 11639 27859 11645
rect 30377 11645 30389 11648
rect 30423 11645 30435 11679
rect 30484 11676 30512 11707
rect 31202 11704 31208 11716
rect 31260 11704 31266 11756
rect 31757 11747 31815 11753
rect 31757 11713 31769 11747
rect 31803 11744 31815 11747
rect 33410 11744 33416 11756
rect 31803 11716 33416 11744
rect 31803 11713 31815 11716
rect 31757 11707 31815 11713
rect 33410 11704 33416 11716
rect 33468 11704 33474 11756
rect 37553 11747 37611 11753
rect 37553 11713 37565 11747
rect 37599 11744 37611 11747
rect 38194 11744 38200 11756
rect 37599 11716 38200 11744
rect 37599 11713 37611 11716
rect 37553 11707 37611 11713
rect 38194 11704 38200 11716
rect 38252 11704 38258 11756
rect 31846 11676 31852 11688
rect 30484 11648 31852 11676
rect 30377 11639 30435 11645
rect 31846 11636 31852 11648
rect 31904 11676 31910 11688
rect 32953 11679 33011 11685
rect 32953 11676 32965 11679
rect 31904 11648 32965 11676
rect 31904 11636 31910 11648
rect 32953 11645 32965 11648
rect 32999 11676 33011 11679
rect 38378 11676 38384 11688
rect 32999 11648 38384 11676
rect 32999 11645 33011 11648
rect 32953 11639 33011 11645
rect 38378 11636 38384 11648
rect 38436 11636 38442 11688
rect 18782 11608 18788 11620
rect 17696 11580 18788 11608
rect 17221 11571 17279 11577
rect 18782 11568 18788 11580
rect 18840 11568 18846 11620
rect 21450 11608 21456 11620
rect 18892 11580 21456 11608
rect 5718 11540 5724 11552
rect 5679 11512 5724 11540
rect 5718 11500 5724 11512
rect 5776 11500 5782 11552
rect 14369 11543 14427 11549
rect 14369 11509 14381 11543
rect 14415 11540 14427 11543
rect 17034 11540 17040 11552
rect 14415 11512 17040 11540
rect 14415 11509 14427 11512
rect 14369 11503 14427 11509
rect 17034 11500 17040 11512
rect 17092 11500 17098 11552
rect 17402 11500 17408 11552
rect 17460 11540 17466 11552
rect 18892 11540 18920 11580
rect 21450 11568 21456 11580
rect 21508 11608 21514 11620
rect 23201 11611 23259 11617
rect 23201 11608 23213 11611
rect 21508 11580 23213 11608
rect 21508 11568 21514 11580
rect 23201 11577 23213 11580
rect 23247 11577 23259 11611
rect 23201 11571 23259 11577
rect 24397 11611 24455 11617
rect 24397 11577 24409 11611
rect 24443 11608 24455 11611
rect 25869 11611 25927 11617
rect 25869 11608 25881 11611
rect 24443 11580 25881 11608
rect 24443 11577 24455 11580
rect 24397 11571 24455 11577
rect 25869 11577 25881 11580
rect 25915 11577 25927 11611
rect 25869 11571 25927 11577
rect 17460 11512 18920 11540
rect 17460 11500 17466 11512
rect 20070 11500 20076 11552
rect 20128 11540 20134 11552
rect 21910 11540 21916 11552
rect 20128 11512 21916 11540
rect 20128 11500 20134 11512
rect 21910 11500 21916 11512
rect 21968 11500 21974 11552
rect 22002 11500 22008 11552
rect 22060 11540 22066 11552
rect 24412 11540 24440 11571
rect 28166 11568 28172 11620
rect 28224 11608 28230 11620
rect 28445 11611 28503 11617
rect 28445 11608 28457 11611
rect 28224 11580 28457 11608
rect 28224 11568 28230 11580
rect 28445 11577 28457 11580
rect 28491 11577 28503 11611
rect 28445 11571 28503 11577
rect 28534 11568 28540 11620
rect 28592 11608 28598 11620
rect 31110 11608 31116 11620
rect 28592 11580 31116 11608
rect 28592 11568 28598 11580
rect 31110 11568 31116 11580
rect 31168 11568 31174 11620
rect 38010 11608 38016 11620
rect 37971 11580 38016 11608
rect 38010 11568 38016 11580
rect 38068 11568 38074 11620
rect 22060 11512 24440 11540
rect 22060 11500 22066 11512
rect 29086 11500 29092 11552
rect 29144 11540 29150 11552
rect 29733 11543 29791 11549
rect 29733 11540 29745 11543
rect 29144 11512 29745 11540
rect 29144 11500 29150 11512
rect 29733 11509 29745 11512
rect 29779 11509 29791 11543
rect 29733 11503 29791 11509
rect 31202 11500 31208 11552
rect 31260 11540 31266 11552
rect 32401 11543 32459 11549
rect 32401 11540 32413 11543
rect 31260 11512 32413 11540
rect 31260 11500 31266 11512
rect 32401 11509 32413 11512
rect 32447 11540 32459 11543
rect 33413 11543 33471 11549
rect 33413 11540 33425 11543
rect 32447 11512 33425 11540
rect 32447 11509 32459 11512
rect 32401 11503 32459 11509
rect 33413 11509 33425 11512
rect 33459 11509 33471 11543
rect 33413 11503 33471 11509
rect 36909 11543 36967 11549
rect 36909 11509 36921 11543
rect 36955 11540 36967 11543
rect 37366 11540 37372 11552
rect 36955 11512 37372 11540
rect 36955 11509 36967 11512
rect 36909 11503 36967 11509
rect 37366 11500 37372 11512
rect 37424 11500 37430 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 12437 11339 12495 11345
rect 12437 11305 12449 11339
rect 12483 11336 12495 11339
rect 15470 11336 15476 11348
rect 12483 11308 15476 11336
rect 12483 11305 12495 11308
rect 12437 11299 12495 11305
rect 15470 11296 15476 11308
rect 15528 11296 15534 11348
rect 15654 11336 15660 11348
rect 15567 11308 15660 11336
rect 15580 11277 15608 11308
rect 15654 11296 15660 11308
rect 15712 11336 15718 11348
rect 15712 11308 20944 11336
rect 15712 11296 15718 11308
rect 15565 11271 15623 11277
rect 15565 11237 15577 11271
rect 15611 11237 15623 11271
rect 20806 11268 20812 11280
rect 15565 11231 15623 11237
rect 16224 11240 17540 11268
rect 14369 11203 14427 11209
rect 14369 11169 14381 11203
rect 14415 11200 14427 11203
rect 16224 11200 16252 11240
rect 16390 11200 16396 11212
rect 14415 11172 16252 11200
rect 16351 11172 16396 11200
rect 14415 11169 14427 11172
rect 14369 11163 14427 11169
rect 16390 11160 16396 11172
rect 16448 11160 16454 11212
rect 17037 11203 17095 11209
rect 17037 11169 17049 11203
rect 17083 11200 17095 11203
rect 17402 11200 17408 11212
rect 17083 11172 17408 11200
rect 17083 11169 17095 11172
rect 17037 11163 17095 11169
rect 17402 11160 17408 11172
rect 17460 11160 17466 11212
rect 5534 11092 5540 11144
rect 5592 11132 5598 11144
rect 6362 11132 6368 11144
rect 5592 11104 6368 11132
rect 5592 11092 5598 11104
rect 6362 11092 6368 11104
rect 6420 11132 6426 11144
rect 11793 11135 11851 11141
rect 11793 11132 11805 11135
rect 6420 11104 11805 11132
rect 6420 11092 6426 11104
rect 11793 11101 11805 11104
rect 11839 11132 11851 11135
rect 12345 11135 12403 11141
rect 12345 11132 12357 11135
rect 11839 11104 12357 11132
rect 11839 11101 11851 11104
rect 11793 11095 11851 11101
rect 12345 11101 12357 11104
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 13354 11092 13360 11144
rect 13412 11132 13418 11144
rect 13538 11132 13544 11144
rect 13412 11104 13544 11132
rect 13412 11092 13418 11104
rect 13538 11092 13544 11104
rect 13596 11092 13602 11144
rect 14274 11132 14280 11144
rect 14235 11104 14280 11132
rect 14274 11092 14280 11104
rect 14332 11092 14338 11144
rect 17512 11132 17540 11240
rect 17696 11240 20812 11268
rect 17696 11209 17724 11240
rect 20806 11228 20812 11240
rect 20864 11228 20870 11280
rect 20916 11268 20944 11308
rect 20990 11296 20996 11348
rect 21048 11336 21054 11348
rect 21048 11308 23612 11336
rect 21048 11296 21054 11308
rect 22830 11268 22836 11280
rect 20916 11240 22836 11268
rect 22830 11228 22836 11240
rect 22888 11228 22894 11280
rect 23474 11268 23480 11280
rect 22940 11240 23480 11268
rect 17681 11203 17739 11209
rect 17681 11169 17693 11203
rect 17727 11169 17739 11203
rect 17681 11163 17739 11169
rect 18233 11203 18291 11209
rect 18233 11169 18245 11203
rect 18279 11200 18291 11203
rect 18322 11200 18328 11212
rect 18279 11172 18328 11200
rect 18279 11169 18291 11172
rect 18233 11163 18291 11169
rect 18322 11160 18328 11172
rect 18380 11160 18386 11212
rect 18598 11200 18604 11212
rect 18559 11172 18604 11200
rect 18598 11160 18604 11172
rect 18656 11160 18662 11212
rect 20162 11160 20168 11212
rect 20220 11200 20226 11212
rect 20257 11203 20315 11209
rect 20257 11200 20269 11203
rect 20220 11172 20269 11200
rect 20220 11160 20226 11172
rect 20257 11169 20269 11172
rect 20303 11169 20315 11203
rect 22002 11200 22008 11212
rect 20257 11163 20315 11169
rect 20824 11172 22008 11200
rect 18046 11132 18052 11144
rect 17512 11104 18052 11132
rect 18046 11092 18052 11104
rect 18104 11092 18110 11144
rect 13633 11067 13691 11073
rect 13633 11033 13645 11067
rect 13679 11064 13691 11067
rect 15010 11064 15016 11076
rect 13679 11036 15016 11064
rect 13679 11033 13691 11036
rect 13633 11027 13691 11033
rect 15010 11024 15016 11036
rect 15068 11024 15074 11076
rect 15102 11024 15108 11076
rect 15160 11064 15166 11076
rect 15160 11036 15205 11064
rect 15160 11024 15166 11036
rect 16482 11024 16488 11076
rect 16540 11064 16546 11076
rect 17954 11064 17960 11076
rect 16540 11036 16585 11064
rect 16684 11036 17960 11064
rect 16540 11024 16546 11036
rect 13081 10999 13139 11005
rect 13081 10965 13093 10999
rect 13127 10996 13139 10999
rect 14274 10996 14280 11008
rect 13127 10968 14280 10996
rect 13127 10965 13139 10968
rect 13081 10959 13139 10965
rect 14274 10956 14280 10968
rect 14332 10996 14338 11008
rect 15194 10996 15200 11008
rect 14332 10968 15200 10996
rect 14332 10956 14338 10968
rect 15194 10956 15200 10968
rect 15252 10956 15258 11008
rect 15470 10956 15476 11008
rect 15528 10996 15534 11008
rect 16684 10996 16712 11036
rect 17954 11024 17960 11036
rect 18012 11024 18018 11076
rect 18322 11064 18328 11076
rect 18283 11036 18328 11064
rect 18322 11024 18328 11036
rect 18380 11024 18386 11076
rect 19058 11024 19064 11076
rect 19116 11064 19122 11076
rect 19981 11067 20039 11073
rect 19981 11064 19993 11067
rect 19116 11036 19993 11064
rect 19116 11024 19122 11036
rect 19981 11033 19993 11036
rect 20027 11033 20039 11067
rect 19981 11027 20039 11033
rect 15528 10968 16712 10996
rect 15528 10956 15534 10968
rect 16758 10956 16764 11008
rect 16816 10996 16822 11008
rect 17862 10996 17868 11008
rect 16816 10968 17868 10996
rect 16816 10956 16822 10968
rect 17862 10956 17868 10968
rect 17920 10956 17926 11008
rect 19996 10996 20024 11027
rect 20070 11024 20076 11076
rect 20128 11064 20134 11076
rect 20824 11064 20852 11172
rect 22002 11160 22008 11172
rect 22060 11160 22066 11212
rect 22097 11203 22155 11209
rect 22097 11169 22109 11203
rect 22143 11200 22155 11203
rect 22940 11200 22968 11240
rect 23474 11228 23480 11240
rect 23532 11228 23538 11280
rect 23584 11268 23612 11308
rect 23842 11296 23848 11348
rect 23900 11336 23906 11348
rect 23937 11339 23995 11345
rect 23937 11336 23949 11339
rect 23900 11308 23949 11336
rect 23900 11296 23906 11308
rect 23937 11305 23949 11308
rect 23983 11305 23995 11339
rect 27062 11336 27068 11348
rect 27023 11308 27068 11336
rect 23937 11299 23995 11305
rect 27062 11296 27068 11308
rect 27120 11296 27126 11348
rect 27246 11296 27252 11348
rect 27304 11336 27310 11348
rect 29086 11336 29092 11348
rect 27304 11308 29092 11336
rect 27304 11296 27310 11308
rect 29086 11296 29092 11308
rect 29144 11296 29150 11348
rect 30466 11336 30472 11348
rect 30427 11308 30472 11336
rect 30466 11296 30472 11308
rect 30524 11296 30530 11348
rect 31665 11339 31723 11345
rect 31665 11305 31677 11339
rect 31711 11336 31723 11339
rect 31846 11336 31852 11348
rect 31711 11308 31852 11336
rect 31711 11305 31723 11308
rect 31665 11299 31723 11305
rect 31846 11296 31852 11308
rect 31904 11296 31910 11348
rect 32217 11339 32275 11345
rect 32217 11305 32229 11339
rect 32263 11336 32275 11339
rect 34790 11336 34796 11348
rect 32263 11308 34796 11336
rect 32263 11305 32275 11308
rect 32217 11299 32275 11305
rect 24578 11268 24584 11280
rect 23584 11240 24584 11268
rect 24578 11228 24584 11240
rect 24636 11228 24642 11280
rect 27706 11268 27712 11280
rect 27667 11240 27712 11268
rect 27706 11228 27712 11240
rect 27764 11228 27770 11280
rect 29825 11271 29883 11277
rect 29825 11268 29837 11271
rect 27816 11240 29837 11268
rect 24946 11200 24952 11212
rect 22143 11172 22968 11200
rect 24504 11172 24952 11200
rect 22143 11169 22155 11172
rect 22097 11163 22155 11169
rect 21450 11132 21456 11144
rect 21411 11104 21456 11132
rect 21450 11092 21456 11104
rect 21508 11092 21514 11144
rect 23750 11092 23756 11144
rect 23808 11132 23814 11144
rect 24029 11135 24087 11141
rect 24029 11132 24041 11135
rect 23808 11104 24041 11132
rect 23808 11092 23814 11104
rect 24029 11101 24041 11104
rect 24075 11101 24087 11135
rect 24029 11095 24087 11101
rect 20128 11036 20173 11064
rect 20272 11036 20852 11064
rect 20128 11024 20134 11036
rect 20272 10996 20300 11036
rect 21634 11024 21640 11076
rect 21692 11064 21698 11076
rect 22005 11067 22063 11073
rect 22005 11064 22017 11067
rect 21692 11036 22017 11064
rect 21692 11024 21698 11036
rect 22005 11033 22017 11036
rect 22051 11033 22063 11067
rect 22646 11064 22652 11076
rect 22607 11036 22652 11064
rect 22005 11027 22063 11033
rect 22646 11024 22652 11036
rect 22704 11024 22710 11076
rect 23198 11064 23204 11076
rect 23159 11036 23204 11064
rect 23198 11024 23204 11036
rect 23256 11024 23262 11076
rect 23293 11067 23351 11073
rect 23293 11033 23305 11067
rect 23339 11064 23351 11067
rect 24504 11064 24532 11172
rect 24946 11160 24952 11172
rect 25004 11160 25010 11212
rect 25222 11200 25228 11212
rect 25183 11172 25228 11200
rect 25222 11160 25228 11172
rect 25280 11160 25286 11212
rect 26142 11200 26148 11212
rect 26103 11172 26148 11200
rect 26142 11160 26148 11172
rect 26200 11160 26206 11212
rect 26234 11160 26240 11212
rect 26292 11200 26298 11212
rect 27816 11200 27844 11240
rect 29825 11237 29837 11240
rect 29871 11237 29883 11271
rect 29825 11231 29883 11237
rect 29914 11228 29920 11280
rect 29972 11268 29978 11280
rect 32232 11268 32260 11299
rect 34790 11296 34796 11308
rect 34848 11296 34854 11348
rect 29972 11240 32260 11268
rect 29972 11228 29978 11240
rect 26292 11172 27844 11200
rect 26292 11160 26298 11172
rect 28350 11160 28356 11212
rect 28408 11200 28414 11212
rect 29730 11200 29736 11212
rect 28408 11172 29736 11200
rect 28408 11160 28414 11172
rect 29730 11160 29736 11172
rect 29788 11160 29794 11212
rect 30466 11160 30472 11212
rect 30524 11200 30530 11212
rect 31662 11200 31668 11212
rect 30524 11172 31668 11200
rect 30524 11160 30530 11172
rect 31662 11160 31668 11172
rect 31720 11160 31726 11212
rect 28537 11135 28595 11141
rect 28537 11132 28549 11135
rect 26620 11104 28549 11132
rect 23339 11036 24532 11064
rect 23339 11033 23351 11036
rect 23293 11027 23351 11033
rect 24578 11024 24584 11076
rect 24636 11064 24642 11076
rect 25130 11064 25136 11076
rect 24636 11036 24681 11064
rect 25091 11036 25136 11064
rect 24636 11024 24642 11036
rect 25130 11024 25136 11036
rect 25188 11024 25194 11076
rect 25222 11024 25228 11076
rect 25280 11064 25286 11076
rect 25869 11067 25927 11073
rect 25869 11064 25881 11067
rect 25280 11036 25881 11064
rect 25280 11024 25286 11036
rect 25869 11033 25881 11036
rect 25915 11033 25927 11067
rect 25869 11027 25927 11033
rect 25961 11067 26019 11073
rect 25961 11033 25973 11067
rect 26007 11064 26019 11067
rect 26007 11036 26464 11064
rect 26007 11033 26019 11036
rect 25961 11027 26019 11033
rect 19996 10968 20300 10996
rect 20714 10956 20720 11008
rect 20772 10996 20778 11008
rect 21726 10996 21732 11008
rect 20772 10968 21732 10996
rect 20772 10956 20778 10968
rect 21726 10956 21732 10968
rect 21784 10956 21790 11008
rect 26436 10996 26464 11036
rect 26620 10996 26648 11104
rect 28537 11101 28549 11104
rect 28583 11101 28595 11135
rect 28537 11095 28595 11101
rect 28629 11135 28687 11141
rect 28629 11101 28641 11135
rect 28675 11132 28687 11135
rect 28718 11132 28724 11144
rect 28675 11104 28724 11132
rect 28675 11101 28687 11104
rect 28629 11095 28687 11101
rect 28718 11092 28724 11104
rect 28776 11092 28782 11144
rect 29086 11132 29092 11144
rect 29047 11104 29092 11132
rect 29086 11092 29092 11104
rect 29144 11092 29150 11144
rect 29178 11092 29184 11144
rect 29236 11132 29242 11144
rect 29914 11132 29920 11144
rect 29236 11104 29920 11132
rect 29236 11092 29242 11104
rect 29914 11092 29920 11104
rect 29972 11092 29978 11144
rect 30558 11132 30564 11144
rect 30519 11104 30564 11132
rect 30558 11092 30564 11104
rect 30616 11132 30622 11144
rect 30616 11104 31754 11132
rect 30616 11092 30622 11104
rect 27157 11067 27215 11073
rect 27157 11033 27169 11067
rect 27203 11064 27215 11067
rect 27798 11064 27804 11076
rect 27203 11036 27804 11064
rect 27203 11033 27215 11036
rect 27157 11027 27215 11033
rect 27798 11024 27804 11036
rect 27856 11024 27862 11076
rect 27893 11067 27951 11073
rect 27893 11033 27905 11067
rect 27939 11064 27951 11067
rect 30282 11064 30288 11076
rect 27939 11036 30288 11064
rect 27939 11033 27951 11036
rect 27893 11027 27951 11033
rect 30282 11024 30288 11036
rect 30340 11024 30346 11076
rect 31021 11067 31079 11073
rect 31021 11064 31033 11067
rect 30392 11036 31033 11064
rect 26436 10968 26648 10996
rect 26786 10956 26792 11008
rect 26844 10996 26850 11008
rect 29178 10996 29184 11008
rect 26844 10968 29184 10996
rect 26844 10956 26850 10968
rect 29178 10956 29184 10968
rect 29236 10956 29242 11008
rect 29638 10956 29644 11008
rect 29696 10996 29702 11008
rect 30392 10996 30420 11036
rect 31021 11033 31033 11036
rect 31067 11033 31079 11067
rect 31726 11064 31754 11104
rect 32769 11067 32827 11073
rect 32769 11064 32781 11067
rect 31726 11036 32781 11064
rect 31021 11027 31079 11033
rect 32769 11033 32781 11036
rect 32815 11064 32827 11067
rect 33870 11064 33876 11076
rect 32815 11036 33876 11064
rect 32815 11033 32827 11036
rect 32769 11027 32827 11033
rect 33870 11024 33876 11036
rect 33928 11024 33934 11076
rect 34514 11024 34520 11076
rect 34572 11064 34578 11076
rect 35621 11067 35679 11073
rect 35621 11064 35633 11067
rect 34572 11036 35633 11064
rect 34572 11024 34578 11036
rect 35621 11033 35633 11036
rect 35667 11064 35679 11067
rect 35802 11064 35808 11076
rect 35667 11036 35808 11064
rect 35667 11033 35679 11036
rect 35621 11027 35679 11033
rect 35802 11024 35808 11036
rect 35860 11024 35866 11076
rect 36078 11064 36084 11076
rect 36039 11036 36084 11064
rect 36078 11024 36084 11036
rect 36136 11024 36142 11076
rect 36725 11067 36783 11073
rect 36725 11033 36737 11067
rect 36771 11064 36783 11067
rect 36814 11064 36820 11076
rect 36771 11036 36820 11064
rect 36771 11033 36783 11036
rect 36725 11027 36783 11033
rect 36814 11024 36820 11036
rect 36872 11024 36878 11076
rect 36906 11024 36912 11076
rect 36964 11064 36970 11076
rect 37277 11067 37335 11073
rect 37277 11064 37289 11067
rect 36964 11036 37289 11064
rect 36964 11024 36970 11036
rect 37277 11033 37289 11036
rect 37323 11033 37335 11067
rect 37277 11027 37335 11033
rect 38102 11024 38108 11076
rect 38160 11064 38166 11076
rect 38197 11067 38255 11073
rect 38197 11064 38209 11067
rect 38160 11036 38209 11064
rect 38160 11024 38166 11036
rect 38197 11033 38209 11036
rect 38243 11033 38255 11067
rect 38197 11027 38255 11033
rect 29696 10968 30420 10996
rect 29696 10956 29702 10968
rect 30926 10956 30932 11008
rect 30984 10996 30990 11008
rect 32858 10996 32864 11008
rect 30984 10968 32864 10996
rect 30984 10956 30990 10968
rect 32858 10956 32864 10968
rect 32916 10956 32922 11008
rect 35069 10999 35127 11005
rect 35069 10965 35081 10999
rect 35115 10996 35127 10999
rect 35710 10996 35716 11008
rect 35115 10968 35716 10996
rect 35115 10965 35127 10968
rect 35069 10959 35127 10965
rect 35710 10956 35716 10968
rect 35768 10956 35774 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 21542 10792 21548 10804
rect 14476 10764 21548 10792
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10656 1915 10659
rect 5718 10656 5724 10668
rect 1903 10628 5724 10656
rect 1903 10625 1915 10628
rect 1857 10619 1915 10625
rect 5718 10616 5724 10628
rect 5776 10616 5782 10668
rect 14476 10665 14504 10764
rect 21542 10752 21548 10764
rect 21600 10752 21606 10804
rect 23753 10795 23811 10801
rect 23753 10761 23765 10795
rect 23799 10792 23811 10795
rect 28166 10792 28172 10804
rect 23799 10764 28172 10792
rect 23799 10761 23811 10764
rect 23753 10755 23811 10761
rect 28166 10752 28172 10764
rect 28224 10752 28230 10804
rect 29273 10795 29331 10801
rect 29273 10761 29285 10795
rect 29319 10792 29331 10795
rect 29822 10792 29828 10804
rect 29319 10764 29828 10792
rect 29319 10761 29331 10764
rect 29273 10755 29331 10761
rect 29822 10752 29828 10764
rect 29880 10752 29886 10804
rect 30098 10752 30104 10804
rect 30156 10792 30162 10804
rect 33321 10795 33379 10801
rect 33321 10792 33333 10795
rect 30156 10764 33333 10792
rect 30156 10752 30162 10764
rect 33321 10761 33333 10764
rect 33367 10761 33379 10795
rect 33321 10755 33379 10761
rect 14642 10684 14648 10736
rect 14700 10724 14706 10736
rect 15105 10727 15163 10733
rect 15105 10724 15117 10727
rect 14700 10696 15117 10724
rect 14700 10684 14706 10696
rect 15105 10693 15117 10696
rect 15151 10693 15163 10727
rect 17313 10727 17371 10733
rect 17313 10724 17325 10727
rect 15105 10687 15163 10693
rect 17052 10696 17325 10724
rect 17052 10668 17080 10696
rect 17313 10693 17325 10696
rect 17359 10693 17371 10727
rect 18506 10724 18512 10736
rect 18467 10696 18512 10724
rect 17313 10687 17371 10693
rect 18506 10684 18512 10696
rect 18564 10684 18570 10736
rect 19058 10724 19064 10736
rect 19019 10696 19064 10724
rect 19058 10684 19064 10696
rect 19116 10684 19122 10736
rect 19334 10684 19340 10736
rect 19392 10724 19398 10736
rect 19705 10727 19763 10733
rect 19705 10724 19717 10727
rect 19392 10696 19717 10724
rect 19392 10684 19398 10696
rect 19705 10693 19717 10696
rect 19751 10693 19763 10727
rect 19705 10687 19763 10693
rect 20070 10684 20076 10736
rect 20128 10724 20134 10736
rect 20901 10727 20959 10733
rect 20901 10724 20913 10727
rect 20128 10696 20913 10724
rect 20128 10684 20134 10696
rect 20901 10693 20913 10696
rect 20947 10693 20959 10727
rect 20901 10687 20959 10693
rect 21453 10727 21511 10733
rect 21453 10693 21465 10727
rect 21499 10724 21511 10727
rect 22554 10724 22560 10736
rect 21499 10696 22560 10724
rect 21499 10693 21511 10696
rect 21453 10687 21511 10693
rect 14461 10659 14519 10665
rect 14461 10625 14473 10659
rect 14507 10625 14519 10659
rect 16114 10656 16120 10668
rect 16075 10628 16120 10656
rect 14461 10619 14519 10625
rect 16114 10616 16120 10628
rect 16172 10616 16178 10668
rect 17034 10616 17040 10668
rect 17092 10616 17098 10668
rect 20254 10616 20260 10668
rect 20312 10656 20318 10668
rect 20312 10628 20357 10656
rect 20312 10616 20318 10628
rect 15010 10588 15016 10600
rect 14971 10560 15016 10588
rect 15010 10548 15016 10560
rect 15068 10548 15074 10600
rect 17218 10588 17224 10600
rect 17179 10560 17224 10588
rect 17218 10548 17224 10560
rect 17276 10548 17282 10600
rect 18230 10588 18236 10600
rect 17512 10560 18236 10588
rect 14369 10523 14427 10529
rect 14369 10489 14381 10523
rect 14415 10520 14427 10523
rect 15102 10520 15108 10532
rect 14415 10492 15108 10520
rect 14415 10489 14427 10492
rect 14369 10483 14427 10489
rect 15102 10480 15108 10492
rect 15160 10480 15166 10532
rect 15565 10523 15623 10529
rect 15565 10489 15577 10523
rect 15611 10520 15623 10523
rect 15838 10520 15844 10532
rect 15611 10492 15844 10520
rect 15611 10489 15623 10492
rect 15565 10483 15623 10489
rect 15838 10480 15844 10492
rect 15896 10520 15902 10532
rect 17512 10520 17540 10560
rect 18230 10548 18236 10560
rect 18288 10548 18294 10600
rect 18414 10588 18420 10600
rect 18375 10560 18420 10588
rect 18414 10548 18420 10560
rect 18472 10588 18478 10600
rect 19610 10588 19616 10600
rect 18472 10560 19616 10588
rect 18472 10548 18478 10560
rect 19610 10548 19616 10560
rect 19668 10548 19674 10600
rect 20806 10588 20812 10600
rect 20767 10560 20812 10588
rect 20806 10548 20812 10560
rect 20864 10548 20870 10600
rect 17770 10520 17776 10532
rect 15896 10492 17540 10520
rect 17731 10492 17776 10520
rect 15896 10480 15902 10492
rect 17770 10480 17776 10492
rect 17828 10480 17834 10532
rect 18138 10480 18144 10532
rect 18196 10520 18202 10532
rect 21468 10520 21496 10687
rect 22554 10684 22560 10696
rect 22612 10684 22618 10736
rect 22830 10684 22836 10736
rect 22888 10684 22894 10736
rect 23658 10684 23664 10736
rect 23716 10724 23722 10736
rect 24765 10727 24823 10733
rect 24765 10724 24777 10727
rect 23716 10696 24777 10724
rect 23716 10684 23722 10696
rect 24765 10693 24777 10696
rect 24811 10693 24823 10727
rect 24765 10687 24823 10693
rect 24857 10727 24915 10733
rect 24857 10693 24869 10727
rect 24903 10724 24915 10727
rect 25038 10724 25044 10736
rect 24903 10696 25044 10724
rect 24903 10693 24915 10696
rect 24857 10687 24915 10693
rect 25038 10684 25044 10696
rect 25096 10684 25102 10736
rect 25406 10724 25412 10736
rect 25367 10696 25412 10724
rect 25406 10684 25412 10696
rect 25464 10684 25470 10736
rect 25961 10727 26019 10733
rect 25961 10693 25973 10727
rect 26007 10724 26019 10727
rect 27798 10724 27804 10736
rect 26007 10696 27804 10724
rect 26007 10693 26019 10696
rect 25961 10687 26019 10693
rect 27798 10684 27804 10696
rect 27856 10684 27862 10736
rect 29730 10684 29736 10736
rect 29788 10724 29794 10736
rect 29917 10727 29975 10733
rect 29917 10724 29929 10727
rect 29788 10696 29929 10724
rect 29788 10684 29794 10696
rect 29917 10693 29929 10696
rect 29963 10693 29975 10727
rect 29917 10687 29975 10693
rect 22002 10656 22008 10668
rect 21963 10628 22008 10656
rect 22002 10616 22008 10628
rect 22060 10616 22066 10668
rect 30009 10659 30067 10665
rect 21542 10548 21548 10600
rect 21600 10588 21606 10600
rect 22646 10588 22652 10600
rect 21600 10560 22652 10588
rect 21600 10548 21606 10560
rect 22646 10548 22652 10560
rect 22704 10588 22710 10600
rect 24213 10591 24271 10597
rect 24213 10588 24225 10591
rect 22704 10560 24225 10588
rect 22704 10548 22710 10560
rect 24213 10557 24225 10560
rect 24259 10557 24271 10591
rect 24213 10551 24271 10557
rect 26053 10591 26111 10597
rect 26053 10557 26065 10591
rect 26099 10588 26111 10591
rect 26099 10560 26372 10588
rect 26099 10557 26111 10560
rect 26053 10551 26111 10557
rect 18196 10492 21496 10520
rect 18196 10480 18202 10492
rect 24118 10480 24124 10532
rect 24176 10520 24182 10532
rect 26068 10520 26096 10551
rect 24176 10492 26096 10520
rect 24176 10480 24182 10492
rect 1670 10452 1676 10464
rect 1631 10424 1676 10452
rect 1670 10412 1676 10424
rect 1728 10412 1734 10464
rect 13265 10455 13323 10461
rect 13265 10421 13277 10455
rect 13311 10452 13323 10455
rect 13354 10452 13360 10464
rect 13311 10424 13360 10452
rect 13311 10421 13323 10424
rect 13265 10415 13323 10421
rect 13354 10412 13360 10424
rect 13412 10412 13418 10464
rect 13814 10452 13820 10464
rect 13727 10424 13820 10452
rect 13814 10412 13820 10424
rect 13872 10452 13878 10464
rect 16114 10452 16120 10464
rect 13872 10424 16120 10452
rect 13872 10412 13878 10424
rect 16114 10412 16120 10424
rect 16172 10412 16178 10464
rect 16209 10455 16267 10461
rect 16209 10421 16221 10455
rect 16255 10452 16267 10455
rect 20070 10452 20076 10464
rect 16255 10424 20076 10452
rect 16255 10421 16267 10424
rect 16209 10415 16267 10421
rect 20070 10412 20076 10424
rect 20128 10412 20134 10464
rect 20254 10412 20260 10464
rect 20312 10452 20318 10464
rect 22094 10452 22100 10464
rect 20312 10424 22100 10452
rect 20312 10412 20318 10424
rect 22094 10412 22100 10424
rect 22152 10412 22158 10464
rect 22278 10461 22284 10464
rect 22268 10455 22284 10461
rect 22268 10452 22280 10455
rect 22191 10424 22280 10452
rect 22268 10421 22280 10424
rect 22336 10452 22342 10464
rect 22646 10452 22652 10464
rect 22336 10424 22652 10452
rect 22268 10415 22284 10421
rect 22278 10412 22284 10415
rect 22336 10412 22342 10424
rect 22646 10412 22652 10424
rect 22704 10412 22710 10464
rect 26344 10452 26372 10560
rect 27154 10548 27160 10600
rect 27212 10588 27218 10600
rect 27525 10591 27583 10597
rect 27525 10588 27537 10591
rect 27212 10560 27537 10588
rect 27212 10548 27218 10560
rect 27525 10557 27537 10560
rect 27571 10557 27583 10591
rect 27801 10591 27859 10597
rect 27801 10588 27813 10591
rect 27525 10551 27583 10557
rect 27632 10560 27813 10588
rect 26418 10480 26424 10532
rect 26476 10520 26482 10532
rect 27632 10520 27660 10560
rect 27801 10557 27813 10560
rect 27847 10557 27859 10591
rect 28920 10588 28948 10642
rect 30009 10625 30021 10659
rect 30055 10656 30067 10659
rect 30650 10656 30656 10668
rect 30055 10628 30656 10656
rect 30055 10625 30067 10628
rect 30009 10619 30067 10625
rect 30650 10616 30656 10628
rect 30708 10616 30714 10668
rect 33413 10659 33471 10665
rect 33413 10625 33425 10659
rect 33459 10656 33471 10659
rect 33686 10656 33692 10668
rect 33459 10628 33692 10656
rect 33459 10625 33471 10628
rect 33413 10619 33471 10625
rect 33686 10616 33692 10628
rect 33744 10616 33750 10668
rect 34422 10616 34428 10668
rect 34480 10656 34486 10668
rect 38013 10659 38071 10665
rect 38013 10656 38025 10659
rect 34480 10628 38025 10656
rect 34480 10616 34486 10628
rect 38013 10625 38025 10628
rect 38059 10625 38071 10659
rect 38013 10619 38071 10625
rect 34698 10588 34704 10600
rect 28920 10560 34704 10588
rect 27801 10551 27859 10557
rect 34698 10548 34704 10560
rect 34756 10548 34762 10600
rect 38286 10588 38292 10600
rect 38247 10560 38292 10588
rect 38286 10548 38292 10560
rect 38344 10548 38350 10600
rect 26476 10492 27660 10520
rect 26476 10480 26482 10492
rect 29914 10480 29920 10532
rect 29972 10520 29978 10532
rect 31573 10523 31631 10529
rect 31573 10520 31585 10523
rect 29972 10492 31585 10520
rect 29972 10480 29978 10492
rect 31573 10489 31585 10492
rect 31619 10489 31631 10523
rect 31573 10483 31631 10489
rect 34793 10523 34851 10529
rect 34793 10489 34805 10523
rect 34839 10520 34851 10523
rect 35437 10523 35495 10529
rect 35437 10520 35449 10523
rect 34839 10492 35449 10520
rect 34839 10489 34851 10492
rect 34793 10483 34851 10489
rect 35437 10489 35449 10492
rect 35483 10520 35495 10523
rect 35618 10520 35624 10532
rect 35483 10492 35624 10520
rect 35483 10489 35495 10492
rect 35437 10483 35495 10489
rect 35618 10480 35624 10492
rect 35676 10520 35682 10532
rect 36817 10523 36875 10529
rect 36817 10520 36829 10523
rect 35676 10492 36829 10520
rect 35676 10480 35682 10492
rect 36817 10489 36829 10492
rect 36863 10489 36875 10523
rect 36817 10483 36875 10489
rect 30098 10452 30104 10464
rect 26344 10424 30104 10452
rect 30098 10412 30104 10424
rect 30156 10412 30162 10464
rect 30282 10412 30288 10464
rect 30340 10452 30346 10464
rect 30469 10455 30527 10461
rect 30469 10452 30481 10455
rect 30340 10424 30481 10452
rect 30340 10412 30346 10424
rect 30469 10421 30481 10424
rect 30515 10421 30527 10455
rect 30469 10415 30527 10421
rect 30558 10412 30564 10464
rect 30616 10452 30622 10464
rect 31021 10455 31079 10461
rect 31021 10452 31033 10455
rect 30616 10424 31033 10452
rect 30616 10412 30622 10424
rect 31021 10421 31033 10424
rect 31067 10421 31079 10455
rect 32398 10452 32404 10464
rect 32359 10424 32404 10452
rect 31021 10415 31079 10421
rect 32398 10412 32404 10424
rect 32456 10412 32462 10464
rect 33870 10452 33876 10464
rect 33831 10424 33876 10452
rect 33870 10412 33876 10424
rect 33928 10412 33934 10464
rect 35710 10412 35716 10464
rect 35768 10452 35774 10464
rect 36265 10455 36323 10461
rect 36265 10452 36277 10455
rect 35768 10424 36277 10452
rect 35768 10412 35774 10424
rect 36265 10421 36277 10424
rect 36311 10421 36323 10455
rect 36265 10415 36323 10421
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 14642 10248 14648 10260
rect 14603 10220 14648 10248
rect 14642 10208 14648 10220
rect 14700 10208 14706 10260
rect 14734 10208 14740 10260
rect 14792 10248 14798 10260
rect 18414 10248 18420 10260
rect 14792 10220 18420 10248
rect 14792 10208 14798 10220
rect 18414 10208 18420 10220
rect 18472 10208 18478 10260
rect 18782 10248 18788 10260
rect 18743 10220 18788 10248
rect 18782 10208 18788 10220
rect 18840 10208 18846 10260
rect 19610 10208 19616 10260
rect 19668 10248 19674 10260
rect 21818 10248 21824 10260
rect 19668 10220 21824 10248
rect 19668 10208 19674 10220
rect 21818 10208 21824 10220
rect 21876 10208 21882 10260
rect 22186 10208 22192 10260
rect 22244 10248 22250 10260
rect 22738 10248 22744 10260
rect 22244 10220 22744 10248
rect 22244 10208 22250 10220
rect 22738 10208 22744 10220
rect 22796 10248 22802 10260
rect 23106 10248 23112 10260
rect 22796 10220 23112 10248
rect 22796 10208 22802 10220
rect 23106 10208 23112 10220
rect 23164 10248 23170 10260
rect 24673 10251 24731 10257
rect 23164 10220 24624 10248
rect 23164 10208 23170 10220
rect 14090 10140 14096 10192
rect 14148 10180 14154 10192
rect 16669 10183 16727 10189
rect 14148 10152 15976 10180
rect 14148 10140 14154 10152
rect 15654 10112 15660 10124
rect 14752 10084 15660 10112
rect 14752 10053 14780 10084
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 15838 10112 15844 10124
rect 15799 10084 15844 10112
rect 15838 10072 15844 10084
rect 15896 10072 15902 10124
rect 15948 10112 15976 10152
rect 16669 10149 16681 10183
rect 16715 10180 16727 10183
rect 18874 10180 18880 10192
rect 16715 10152 18880 10180
rect 16715 10149 16727 10152
rect 16669 10143 16727 10149
rect 18874 10140 18880 10152
rect 18932 10140 18938 10192
rect 20530 10140 20536 10192
rect 20588 10140 20594 10192
rect 21910 10140 21916 10192
rect 21968 10180 21974 10192
rect 22281 10183 22339 10189
rect 22281 10180 22293 10183
rect 21968 10152 22293 10180
rect 21968 10140 21974 10152
rect 22281 10149 22293 10152
rect 22327 10149 22339 10183
rect 22281 10143 22339 10149
rect 22554 10140 22560 10192
rect 22612 10180 22618 10192
rect 22925 10183 22983 10189
rect 22925 10180 22937 10183
rect 22612 10152 22937 10180
rect 22612 10140 22618 10152
rect 22925 10149 22937 10152
rect 22971 10180 22983 10183
rect 24302 10180 24308 10192
rect 22971 10152 24308 10180
rect 22971 10149 22983 10152
rect 22925 10143 22983 10149
rect 24302 10140 24308 10152
rect 24360 10140 24366 10192
rect 24596 10180 24624 10220
rect 24673 10217 24685 10251
rect 24719 10248 24731 10251
rect 24854 10248 24860 10260
rect 24719 10220 24860 10248
rect 24719 10217 24731 10220
rect 24673 10211 24731 10217
rect 24854 10208 24860 10220
rect 24912 10208 24918 10260
rect 26142 10208 26148 10260
rect 26200 10248 26206 10260
rect 29638 10248 29644 10260
rect 26200 10220 29644 10248
rect 26200 10208 26206 10220
rect 29638 10208 29644 10220
rect 29696 10248 29702 10260
rect 29733 10251 29791 10257
rect 29733 10248 29745 10251
rect 29696 10220 29745 10248
rect 29696 10208 29702 10220
rect 29733 10217 29745 10220
rect 29779 10217 29791 10251
rect 29733 10211 29791 10217
rect 30190 10208 30196 10260
rect 30248 10248 30254 10260
rect 32033 10251 32091 10257
rect 32033 10248 32045 10251
rect 30248 10220 32045 10248
rect 30248 10208 30254 10220
rect 32033 10217 32045 10220
rect 32079 10217 32091 10251
rect 32033 10211 32091 10217
rect 36633 10251 36691 10257
rect 36633 10217 36645 10251
rect 36679 10248 36691 10251
rect 36906 10248 36912 10260
rect 36679 10220 36912 10248
rect 36679 10217 36691 10220
rect 36633 10211 36691 10217
rect 36906 10208 36912 10220
rect 36964 10208 36970 10260
rect 37642 10248 37648 10260
rect 37603 10220 37648 10248
rect 37642 10208 37648 10220
rect 37700 10208 37706 10260
rect 38286 10248 38292 10260
rect 38247 10220 38292 10248
rect 38286 10208 38292 10220
rect 38344 10208 38350 10260
rect 24596 10152 25360 10180
rect 17221 10115 17279 10121
rect 17221 10112 17233 10115
rect 15948 10084 17233 10112
rect 17221 10081 17233 10084
rect 17267 10081 17279 10115
rect 17221 10075 17279 10081
rect 17402 10072 17408 10124
rect 17460 10112 17466 10124
rect 17865 10115 17923 10121
rect 17865 10112 17877 10115
rect 17460 10084 17877 10112
rect 17460 10072 17466 10084
rect 17865 10081 17877 10084
rect 17911 10081 17923 10115
rect 20548 10112 20576 10140
rect 20806 10112 20812 10124
rect 17865 10075 17923 10081
rect 18892 10084 20576 10112
rect 20719 10084 20812 10112
rect 13541 10047 13599 10053
rect 13541 10044 13553 10047
rect 13004 10016 13553 10044
rect 12894 9868 12900 9920
rect 12952 9908 12958 9920
rect 13004 9917 13032 10016
rect 13541 10013 13553 10016
rect 13587 10013 13599 10047
rect 13541 10007 13599 10013
rect 14737 10047 14795 10053
rect 14737 10013 14749 10047
rect 14783 10013 14795 10047
rect 16574 10044 16580 10056
rect 16535 10016 16580 10044
rect 14737 10007 14795 10013
rect 16574 10004 16580 10016
rect 16632 10004 16638 10056
rect 18892 10053 18920 10084
rect 20806 10072 20812 10084
rect 20864 10112 20870 10124
rect 21818 10112 21824 10124
rect 20864 10084 21824 10112
rect 20864 10072 20870 10084
rect 21818 10072 21824 10084
rect 21876 10072 21882 10124
rect 22186 10072 22192 10124
rect 22244 10112 22250 10124
rect 23477 10115 23535 10121
rect 23477 10112 23489 10115
rect 22244 10084 23489 10112
rect 22244 10072 22250 10084
rect 23477 10081 23489 10084
rect 23523 10112 23535 10115
rect 25222 10112 25228 10124
rect 23523 10084 25228 10112
rect 23523 10081 23535 10084
rect 23477 10075 23535 10081
rect 25222 10072 25228 10084
rect 25280 10072 25286 10124
rect 25332 10112 25360 10152
rect 26878 10140 26884 10192
rect 26936 10180 26942 10192
rect 28445 10183 28503 10189
rect 28445 10180 28457 10183
rect 26936 10152 28457 10180
rect 26936 10140 26942 10152
rect 28445 10149 28457 10152
rect 28491 10149 28503 10183
rect 28445 10143 28503 10149
rect 28994 10140 29000 10192
rect 29052 10180 29058 10192
rect 29454 10180 29460 10192
rect 29052 10152 29460 10180
rect 29052 10140 29058 10152
rect 29454 10140 29460 10152
rect 29512 10140 29518 10192
rect 30650 10140 30656 10192
rect 30708 10180 30714 10192
rect 31389 10183 31447 10189
rect 31389 10180 31401 10183
rect 30708 10152 31401 10180
rect 30708 10140 30714 10152
rect 31389 10149 31401 10152
rect 31435 10149 31447 10183
rect 31389 10143 31447 10149
rect 25685 10115 25743 10121
rect 25685 10112 25697 10115
rect 25332 10084 25697 10112
rect 25685 10081 25697 10084
rect 25731 10081 25743 10115
rect 25685 10075 25743 10081
rect 27080 10112 27292 10124
rect 34054 10112 34060 10124
rect 27080 10096 34060 10112
rect 18877 10047 18935 10053
rect 18877 10013 18889 10047
rect 18923 10013 18935 10047
rect 18877 10007 18935 10013
rect 19889 10047 19947 10053
rect 19889 10013 19901 10047
rect 19935 10044 19947 10047
rect 20070 10044 20076 10056
rect 19935 10016 20076 10044
rect 19935 10013 19947 10016
rect 19889 10007 19947 10013
rect 20070 10004 20076 10016
rect 20128 10004 20134 10056
rect 20533 10047 20591 10053
rect 20533 10013 20545 10047
rect 20579 10013 20591 10047
rect 20533 10007 20591 10013
rect 15197 9979 15255 9985
rect 15197 9945 15209 9979
rect 15243 9976 15255 9979
rect 15654 9976 15660 9988
rect 15243 9948 15660 9976
rect 15243 9945 15255 9948
rect 15197 9939 15255 9945
rect 15654 9936 15660 9948
rect 15712 9936 15718 9988
rect 15749 9979 15807 9985
rect 15749 9945 15761 9979
rect 15795 9945 15807 9979
rect 17770 9976 17776 9988
rect 17731 9948 17776 9976
rect 15749 9939 15807 9945
rect 12989 9911 13047 9917
rect 12989 9908 13001 9911
rect 12952 9880 13001 9908
rect 12952 9868 12958 9880
rect 12989 9877 13001 9880
rect 13035 9877 13047 9911
rect 12989 9871 13047 9877
rect 13633 9911 13691 9917
rect 13633 9877 13645 9911
rect 13679 9908 13691 9911
rect 15102 9908 15108 9920
rect 13679 9880 15108 9908
rect 13679 9877 13691 9880
rect 13633 9871 13691 9877
rect 15102 9868 15108 9880
rect 15160 9868 15166 9920
rect 15771 9908 15799 9939
rect 17770 9936 17776 9948
rect 17828 9936 17834 9988
rect 20548 9976 20576 10007
rect 21910 10004 21916 10056
rect 21968 10004 21974 10056
rect 24026 10004 24032 10056
rect 24084 10044 24090 10056
rect 24581 10047 24639 10053
rect 24581 10044 24593 10047
rect 24084 10016 24593 10044
rect 24084 10004 24090 10016
rect 24581 10013 24593 10016
rect 24627 10013 24639 10047
rect 24581 10007 24639 10013
rect 25038 10004 25044 10056
rect 25096 10044 25102 10056
rect 25409 10047 25467 10053
rect 25409 10044 25421 10047
rect 25096 10016 25421 10044
rect 25096 10004 25102 10016
rect 25409 10013 25421 10016
rect 25455 10013 25467 10047
rect 27080 10044 27108 10096
rect 27264 10084 34060 10096
rect 34054 10072 34060 10084
rect 34112 10072 34118 10124
rect 27798 10044 27804 10056
rect 26818 10016 27108 10044
rect 27172 10016 27660 10044
rect 27759 10016 27804 10044
rect 25409 10007 25467 10013
rect 20714 9976 20720 9988
rect 20548 9948 20720 9976
rect 20714 9936 20720 9948
rect 20772 9936 20778 9988
rect 23392 9979 23450 9985
rect 23392 9945 23404 9979
rect 23438 9945 23450 9979
rect 23392 9939 23450 9945
rect 16482 9908 16488 9920
rect 15771 9880 16488 9908
rect 16482 9868 16488 9880
rect 16540 9868 16546 9920
rect 16574 9868 16580 9920
rect 16632 9908 16638 9920
rect 17310 9908 17316 9920
rect 16632 9880 17316 9908
rect 16632 9868 16638 9880
rect 17310 9868 17316 9880
rect 17368 9868 17374 9920
rect 19981 9911 20039 9917
rect 19981 9877 19993 9911
rect 20027 9908 20039 9911
rect 22186 9908 22192 9920
rect 20027 9880 22192 9908
rect 20027 9877 20039 9880
rect 19981 9871 20039 9877
rect 22186 9868 22192 9880
rect 22244 9868 22250 9920
rect 23400 9908 23428 9939
rect 24670 9908 24676 9920
rect 23400 9880 24676 9908
rect 24670 9868 24676 9880
rect 24728 9868 24734 9920
rect 27172 9917 27200 10016
rect 27632 9976 27660 10016
rect 27798 10004 27804 10016
rect 27856 10004 27862 10056
rect 27893 10047 27951 10053
rect 27893 10013 27905 10047
rect 27939 10013 27951 10047
rect 27893 10007 27951 10013
rect 28537 10047 28595 10053
rect 28537 10013 28549 10047
rect 28583 10044 28595 10047
rect 29638 10044 29644 10056
rect 28583 10016 29644 10044
rect 28583 10013 28595 10016
rect 28537 10007 28595 10013
rect 27908 9976 27936 10007
rect 29638 10004 29644 10016
rect 29696 10004 29702 10056
rect 32125 10047 32183 10053
rect 32125 10013 32137 10047
rect 32171 10044 32183 10047
rect 32306 10044 32312 10056
rect 32171 10016 32312 10044
rect 32171 10013 32183 10016
rect 32125 10007 32183 10013
rect 32306 10004 32312 10016
rect 32364 10004 32370 10056
rect 32398 10004 32404 10056
rect 32456 10044 32462 10056
rect 32677 10047 32735 10053
rect 32677 10044 32689 10047
rect 32456 10016 32689 10044
rect 32456 10004 32462 10016
rect 32677 10013 32689 10016
rect 32723 10044 32735 10047
rect 33229 10047 33287 10053
rect 33229 10044 33241 10047
rect 32723 10016 33241 10044
rect 32723 10013 32735 10016
rect 32677 10007 32735 10013
rect 33229 10013 33241 10016
rect 33275 10044 33287 10047
rect 33781 10047 33839 10053
rect 33781 10044 33793 10047
rect 33275 10016 33793 10044
rect 33275 10013 33287 10016
rect 33229 10007 33287 10013
rect 33781 10013 33793 10016
rect 33827 10044 33839 10047
rect 34241 10047 34299 10053
rect 34241 10044 34253 10047
rect 33827 10016 34253 10044
rect 33827 10013 33839 10016
rect 33781 10007 33839 10013
rect 34241 10013 34253 10016
rect 34287 10013 34299 10047
rect 34241 10007 34299 10013
rect 28902 9976 28908 9988
rect 27632 9948 28908 9976
rect 28902 9936 28908 9948
rect 28960 9936 28966 9988
rect 29086 9976 29092 9988
rect 29047 9948 29092 9976
rect 29086 9936 29092 9948
rect 29144 9976 29150 9988
rect 30282 9976 30288 9988
rect 29144 9948 30288 9976
rect 29144 9936 29150 9948
rect 30282 9936 30288 9948
rect 30340 9976 30346 9988
rect 30837 9979 30895 9985
rect 30837 9976 30849 9979
rect 30340 9948 30849 9976
rect 30340 9936 30346 9948
rect 30837 9945 30849 9948
rect 30883 9976 30895 9979
rect 32416 9976 32444 10004
rect 35710 9976 35716 9988
rect 30883 9948 32444 9976
rect 34992 9948 35716 9976
rect 30883 9945 30895 9948
rect 30837 9939 30895 9945
rect 34992 9920 35020 9948
rect 35710 9936 35716 9948
rect 35768 9976 35774 9988
rect 35989 9979 36047 9985
rect 35989 9976 36001 9979
rect 35768 9948 36001 9976
rect 35768 9936 35774 9948
rect 35989 9945 36001 9948
rect 36035 9976 36047 9979
rect 37093 9979 37151 9985
rect 37093 9976 37105 9979
rect 36035 9948 37105 9976
rect 36035 9945 36047 9948
rect 35989 9939 36047 9945
rect 37093 9945 37105 9948
rect 37139 9945 37151 9979
rect 37093 9939 37151 9945
rect 27157 9911 27215 9917
rect 27157 9877 27169 9911
rect 27203 9877 27215 9911
rect 27157 9871 27215 9877
rect 27246 9868 27252 9920
rect 27304 9908 27310 9920
rect 30650 9908 30656 9920
rect 27304 9880 30656 9908
rect 27304 9868 27310 9880
rect 30650 9868 30656 9880
rect 30708 9868 30714 9920
rect 34974 9908 34980 9920
rect 34935 9880 34980 9908
rect 34974 9868 34980 9880
rect 35032 9868 35038 9920
rect 35434 9908 35440 9920
rect 35395 9880 35440 9908
rect 35434 9868 35440 9880
rect 35492 9868 35498 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 13817 9707 13875 9713
rect 13817 9673 13829 9707
rect 13863 9704 13875 9707
rect 13863 9676 15884 9704
rect 13863 9673 13875 9676
rect 13817 9667 13875 9673
rect 4062 9596 4068 9648
rect 4120 9636 4126 9648
rect 4709 9639 4767 9645
rect 4709 9636 4721 9639
rect 4120 9608 4721 9636
rect 4120 9596 4126 9608
rect 4709 9605 4721 9608
rect 4755 9605 4767 9639
rect 4709 9599 4767 9605
rect 10962 9596 10968 9648
rect 11020 9636 11026 9648
rect 13078 9636 13084 9648
rect 11020 9608 13084 9636
rect 11020 9596 11026 9608
rect 13078 9596 13084 9608
rect 13136 9596 13142 9648
rect 13265 9639 13323 9645
rect 13265 9605 13277 9639
rect 13311 9636 13323 9639
rect 13446 9636 13452 9648
rect 13311 9608 13452 9636
rect 13311 9605 13323 9608
rect 13265 9599 13323 9605
rect 13446 9596 13452 9608
rect 13504 9636 13510 9648
rect 14369 9639 14427 9645
rect 13504 9608 14320 9636
rect 13504 9596 13510 9608
rect 4801 9571 4859 9577
rect 4801 9537 4813 9571
rect 4847 9568 4859 9571
rect 5353 9571 5411 9577
rect 5353 9568 5365 9571
rect 4847 9540 5365 9568
rect 4847 9537 4859 9540
rect 4801 9531 4859 9537
rect 5353 9537 5365 9540
rect 5399 9568 5411 9571
rect 14182 9568 14188 9580
rect 5399 9540 14188 9568
rect 5399 9537 5411 9540
rect 5353 9531 5411 9537
rect 14182 9528 14188 9540
rect 14240 9528 14246 9580
rect 14292 9577 14320 9608
rect 14369 9605 14381 9639
rect 14415 9636 14427 9639
rect 15749 9639 15807 9645
rect 15749 9636 15761 9639
rect 14415 9608 15761 9636
rect 14415 9605 14427 9608
rect 14369 9599 14427 9605
rect 15749 9605 15761 9608
rect 15795 9605 15807 9639
rect 15856 9636 15884 9676
rect 16114 9664 16120 9716
rect 16172 9704 16178 9716
rect 16172 9676 17540 9704
rect 16172 9664 16178 9676
rect 16574 9636 16580 9648
rect 15856 9608 16580 9636
rect 15749 9599 15807 9605
rect 16574 9596 16580 9608
rect 16632 9596 16638 9648
rect 17034 9636 17040 9648
rect 16995 9608 17040 9636
rect 17034 9596 17040 9608
rect 17092 9596 17098 9648
rect 17512 9636 17540 9676
rect 17586 9664 17592 9716
rect 17644 9704 17650 9716
rect 21542 9704 21548 9716
rect 17644 9676 21548 9704
rect 17644 9664 17650 9676
rect 21542 9664 21548 9676
rect 21600 9664 21606 9716
rect 24946 9704 24952 9716
rect 22066 9676 24952 9704
rect 22066 9674 22094 9676
rect 21928 9648 22094 9674
rect 24946 9664 24952 9676
rect 25004 9664 25010 9716
rect 28718 9704 28724 9716
rect 27632 9676 28724 9704
rect 17954 9636 17960 9648
rect 17512 9608 17960 9636
rect 17954 9596 17960 9608
rect 18012 9596 18018 9648
rect 18046 9596 18052 9648
rect 18104 9636 18110 9648
rect 19061 9639 19119 9645
rect 19061 9636 19073 9639
rect 18104 9608 19073 9636
rect 18104 9596 18110 9608
rect 19061 9605 19073 9608
rect 19107 9605 19119 9639
rect 19978 9636 19984 9648
rect 19939 9608 19984 9636
rect 19061 9599 19119 9605
rect 19978 9596 19984 9608
rect 20036 9596 20042 9648
rect 20438 9596 20444 9648
rect 20496 9596 20502 9648
rect 21910 9596 21916 9648
rect 21968 9646 22094 9648
rect 21968 9596 21974 9646
rect 23842 9596 23848 9648
rect 23900 9636 23906 9648
rect 24029 9639 24087 9645
rect 24029 9636 24041 9639
rect 23900 9608 24041 9636
rect 23900 9596 23906 9608
rect 24029 9605 24041 9608
rect 24075 9636 24087 9639
rect 24210 9636 24216 9648
rect 24075 9608 24216 9636
rect 24075 9605 24087 9608
rect 24029 9599 24087 9605
rect 24210 9596 24216 9608
rect 24268 9596 24274 9648
rect 25038 9636 25044 9648
rect 24504 9608 25044 9636
rect 14277 9571 14335 9577
rect 14277 9537 14289 9571
rect 14323 9568 14335 9571
rect 14918 9568 14924 9580
rect 14323 9540 14780 9568
rect 14879 9540 14924 9568
rect 14323 9537 14335 9540
rect 14277 9531 14335 9537
rect 14752 9432 14780 9540
rect 14918 9528 14924 9540
rect 14976 9528 14982 9580
rect 16298 9528 16304 9580
rect 16356 9568 16362 9580
rect 24118 9568 24124 9580
rect 16356 9540 16401 9568
rect 23414 9540 24124 9568
rect 16356 9528 16362 9540
rect 24118 9528 24124 9540
rect 24176 9528 24182 9580
rect 24504 9577 24532 9608
rect 25038 9596 25044 9608
rect 25096 9596 25102 9648
rect 27430 9636 27436 9648
rect 25990 9608 27436 9636
rect 27430 9596 27436 9608
rect 27488 9596 27494 9648
rect 24489 9571 24547 9577
rect 24489 9568 24501 9571
rect 24228 9540 24501 9568
rect 15470 9460 15476 9512
rect 15528 9500 15534 9512
rect 15657 9503 15715 9509
rect 15657 9500 15669 9503
rect 15528 9472 15669 9500
rect 15528 9460 15534 9472
rect 15657 9469 15669 9472
rect 15703 9500 15715 9503
rect 16945 9503 17003 9509
rect 16945 9500 16957 9503
rect 15703 9472 16957 9500
rect 15703 9469 15715 9472
rect 15657 9463 15715 9469
rect 16945 9469 16957 9472
rect 16991 9469 17003 9503
rect 16945 9463 17003 9469
rect 17126 9460 17132 9512
rect 17184 9500 17190 9512
rect 17402 9500 17408 9512
rect 17184 9472 17408 9500
rect 17184 9460 17190 9472
rect 17402 9460 17408 9472
rect 17460 9460 17466 9512
rect 17586 9500 17592 9512
rect 17547 9472 17592 9500
rect 17586 9460 17592 9472
rect 17644 9460 17650 9512
rect 18877 9503 18935 9509
rect 18877 9469 18889 9503
rect 18923 9469 18935 9503
rect 19150 9500 19156 9512
rect 19111 9472 19156 9500
rect 18877 9463 18935 9469
rect 16666 9432 16672 9444
rect 14752 9404 16672 9432
rect 16666 9392 16672 9404
rect 16724 9392 16730 9444
rect 16758 9392 16764 9444
rect 16816 9432 16822 9444
rect 17604 9432 17632 9460
rect 18046 9432 18052 9444
rect 16816 9404 17632 9432
rect 17696 9404 18052 9432
rect 16816 9392 16822 9404
rect 15013 9367 15071 9373
rect 15013 9333 15025 9367
rect 15059 9364 15071 9367
rect 17696 9364 17724 9404
rect 18046 9392 18052 9404
rect 18104 9392 18110 9444
rect 18892 9432 18920 9463
rect 19150 9460 19156 9472
rect 19208 9460 19214 9512
rect 19705 9503 19763 9509
rect 19705 9469 19717 9503
rect 19751 9500 19763 9503
rect 20714 9500 20720 9512
rect 19751 9472 20720 9500
rect 19751 9469 19763 9472
rect 19705 9463 19763 9469
rect 20714 9460 20720 9472
rect 20772 9500 20778 9512
rect 20990 9500 20996 9512
rect 20772 9472 20996 9500
rect 20772 9460 20778 9472
rect 20990 9460 20996 9472
rect 21048 9460 21054 9512
rect 22002 9460 22008 9512
rect 22060 9500 22066 9512
rect 22060 9472 22105 9500
rect 22060 9460 22066 9472
rect 22278 9460 22284 9512
rect 22336 9500 22342 9512
rect 24228 9500 24256 9540
rect 24489 9537 24501 9540
rect 24535 9537 24547 9571
rect 27632 9568 27660 9676
rect 28718 9664 28724 9676
rect 28776 9704 28782 9716
rect 30558 9704 30564 9716
rect 28776 9676 30564 9704
rect 28776 9664 28782 9676
rect 30558 9664 30564 9676
rect 30616 9664 30622 9716
rect 32490 9664 32496 9716
rect 32548 9704 32554 9716
rect 37274 9704 37280 9716
rect 32548 9676 37280 9704
rect 32548 9664 32554 9676
rect 37274 9664 37280 9676
rect 37332 9664 37338 9716
rect 32950 9636 32956 9648
rect 28474 9608 32956 9636
rect 32950 9596 32956 9608
rect 33008 9596 33014 9648
rect 36262 9636 36268 9648
rect 36175 9608 36268 9636
rect 36262 9596 36268 9608
rect 36320 9636 36326 9648
rect 36817 9639 36875 9645
rect 36817 9636 36829 9639
rect 36320 9608 36829 9636
rect 36320 9596 36326 9608
rect 36817 9605 36829 9608
rect 36863 9636 36875 9639
rect 36906 9636 36912 9648
rect 36863 9608 36912 9636
rect 36863 9605 36875 9608
rect 36817 9599 36875 9605
rect 36906 9596 36912 9608
rect 36964 9596 36970 9648
rect 24489 9531 24547 9537
rect 26344 9540 27660 9568
rect 22336 9472 24256 9500
rect 22336 9460 22342 9472
rect 24302 9460 24308 9512
rect 24360 9500 24366 9512
rect 24765 9503 24823 9509
rect 24765 9500 24777 9503
rect 24360 9472 24777 9500
rect 24360 9460 24366 9472
rect 24765 9469 24777 9472
rect 24811 9469 24823 9503
rect 24765 9463 24823 9469
rect 25314 9460 25320 9512
rect 25372 9500 25378 9512
rect 26344 9500 26372 9540
rect 26510 9500 26516 9512
rect 25372 9472 26372 9500
rect 26471 9472 26516 9500
rect 25372 9460 25378 9472
rect 26510 9460 26516 9472
rect 26568 9460 26574 9512
rect 27157 9503 27215 9509
rect 27157 9469 27169 9503
rect 27203 9469 27215 9503
rect 27157 9463 27215 9469
rect 28905 9503 28963 9509
rect 28905 9469 28917 9503
rect 28951 9500 28963 9503
rect 29181 9503 29239 9509
rect 28951 9472 29132 9500
rect 28951 9469 28963 9472
rect 28905 9463 28963 9469
rect 19242 9432 19248 9444
rect 18892 9404 19248 9432
rect 19242 9392 19248 9404
rect 19300 9392 19306 9444
rect 15059 9336 17724 9364
rect 15059 9333 15071 9336
rect 15013 9327 15071 9333
rect 17862 9324 17868 9376
rect 17920 9364 17926 9376
rect 19702 9364 19708 9376
rect 17920 9336 19708 9364
rect 17920 9324 17926 9336
rect 19702 9324 19708 9336
rect 19760 9324 19766 9376
rect 21453 9367 21511 9373
rect 21453 9333 21465 9367
rect 21499 9364 21511 9367
rect 22094 9364 22100 9376
rect 21499 9336 22100 9364
rect 21499 9333 21511 9336
rect 21453 9327 21511 9333
rect 22094 9324 22100 9336
rect 22152 9324 22158 9376
rect 22268 9367 22326 9373
rect 22268 9333 22280 9367
rect 22314 9364 22326 9367
rect 24026 9364 24032 9376
rect 22314 9336 24032 9364
rect 22314 9333 22326 9336
rect 22268 9327 22326 9333
rect 24026 9324 24032 9336
rect 24084 9324 24090 9376
rect 25222 9324 25228 9376
rect 25280 9364 25286 9376
rect 27172 9364 27200 9463
rect 29104 9432 29132 9472
rect 29181 9469 29193 9503
rect 29227 9500 29239 9503
rect 29733 9503 29791 9509
rect 29733 9500 29745 9503
rect 29227 9472 29745 9500
rect 29227 9469 29239 9472
rect 29181 9463 29239 9469
rect 29733 9469 29745 9472
rect 29779 9500 29791 9503
rect 31389 9503 31447 9509
rect 31389 9500 31401 9503
rect 29779 9472 31401 9500
rect 29779 9469 29791 9472
rect 29733 9463 29791 9469
rect 31389 9469 31401 9472
rect 31435 9500 31447 9503
rect 33505 9503 33563 9509
rect 31435 9472 32904 9500
rect 31435 9469 31447 9472
rect 31389 9463 31447 9469
rect 32766 9432 32772 9444
rect 29104 9404 32772 9432
rect 32766 9392 32772 9404
rect 32824 9392 32830 9444
rect 32876 9376 32904 9472
rect 33505 9469 33517 9503
rect 33551 9500 33563 9503
rect 34057 9503 34115 9509
rect 34057 9500 34069 9503
rect 33551 9472 34069 9500
rect 33551 9469 33563 9472
rect 33505 9463 33563 9469
rect 34057 9469 34069 9472
rect 34103 9500 34115 9503
rect 35161 9503 35219 9509
rect 35161 9500 35173 9503
rect 34103 9472 35173 9500
rect 34103 9469 34115 9472
rect 34057 9463 34115 9469
rect 35161 9469 35173 9472
rect 35207 9500 35219 9503
rect 37274 9500 37280 9512
rect 35207 9472 37280 9500
rect 35207 9469 35219 9472
rect 35161 9463 35219 9469
rect 37274 9460 37280 9472
rect 37332 9500 37338 9512
rect 37461 9503 37519 9509
rect 37461 9500 37473 9503
rect 37332 9472 37473 9500
rect 37332 9460 37338 9472
rect 37461 9469 37473 9472
rect 37507 9500 37519 9503
rect 37918 9500 37924 9512
rect 37507 9472 37924 9500
rect 37507 9469 37519 9472
rect 37461 9463 37519 9469
rect 37918 9460 37924 9472
rect 37976 9460 37982 9512
rect 34609 9435 34667 9441
rect 34609 9401 34621 9435
rect 34655 9432 34667 9435
rect 34974 9432 34980 9444
rect 34655 9404 34980 9432
rect 34655 9401 34667 9404
rect 34609 9395 34667 9401
rect 34974 9392 34980 9404
rect 35032 9432 35038 9444
rect 35342 9432 35348 9444
rect 35032 9404 35348 9432
rect 35032 9392 35038 9404
rect 35342 9392 35348 9404
rect 35400 9392 35406 9444
rect 29730 9364 29736 9376
rect 25280 9336 29736 9364
rect 25280 9324 25286 9336
rect 29730 9324 29736 9336
rect 29788 9324 29794 9376
rect 30190 9364 30196 9376
rect 30151 9336 30196 9364
rect 30190 9324 30196 9336
rect 30248 9324 30254 9376
rect 30282 9324 30288 9376
rect 30340 9364 30346 9376
rect 30745 9367 30803 9373
rect 30745 9364 30757 9367
rect 30340 9336 30757 9364
rect 30340 9324 30346 9336
rect 30745 9333 30757 9336
rect 30791 9364 30803 9367
rect 30834 9364 30840 9376
rect 30791 9336 30840 9364
rect 30791 9333 30803 9336
rect 30745 9327 30803 9333
rect 30834 9324 30840 9336
rect 30892 9324 30898 9376
rect 31110 9324 31116 9376
rect 31168 9364 31174 9376
rect 32309 9367 32367 9373
rect 32309 9364 32321 9367
rect 31168 9336 32321 9364
rect 31168 9324 31174 9336
rect 32309 9333 32321 9336
rect 32355 9333 32367 9367
rect 32858 9364 32864 9376
rect 32819 9336 32864 9364
rect 32309 9327 32367 9333
rect 32858 9324 32864 9336
rect 32916 9324 32922 9376
rect 35710 9364 35716 9376
rect 35671 9336 35716 9364
rect 35710 9324 35716 9336
rect 35768 9364 35774 9376
rect 37642 9364 37648 9376
rect 35768 9336 37648 9364
rect 35768 9324 35774 9336
rect 37642 9324 37648 9336
rect 37700 9324 37706 9376
rect 38194 9364 38200 9376
rect 38155 9336 38200 9364
rect 38194 9324 38200 9336
rect 38252 9324 38258 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 15013 9163 15071 9169
rect 15013 9129 15025 9163
rect 15059 9160 15071 9163
rect 17034 9160 17040 9172
rect 15059 9132 17040 9160
rect 15059 9129 15071 9132
rect 15013 9123 15071 9129
rect 17034 9120 17040 9132
rect 17092 9120 17098 9172
rect 17126 9120 17132 9172
rect 17184 9160 17190 9172
rect 23477 9163 23535 9169
rect 17184 9132 23428 9160
rect 17184 9120 17190 9132
rect 1854 9092 1860 9104
rect 1815 9064 1860 9092
rect 1854 9052 1860 9064
rect 1912 9052 1918 9104
rect 16850 9092 16856 9104
rect 15488 9064 16856 9092
rect 13538 8916 13544 8968
rect 13596 8956 13602 8968
rect 13725 8959 13783 8965
rect 13725 8956 13737 8959
rect 13596 8928 13737 8956
rect 13596 8916 13602 8928
rect 13725 8925 13737 8928
rect 13771 8956 13783 8959
rect 14274 8956 14280 8968
rect 13771 8928 14280 8956
rect 13771 8925 13783 8928
rect 13725 8919 13783 8925
rect 14274 8916 14280 8928
rect 14332 8916 14338 8968
rect 14918 8956 14924 8968
rect 14831 8928 14924 8956
rect 14918 8916 14924 8928
rect 14976 8956 14982 8968
rect 15488 8956 15516 9064
rect 16850 9052 16856 9064
rect 16908 9052 16914 9104
rect 16945 9095 17003 9101
rect 16945 9061 16957 9095
rect 16991 9092 17003 9095
rect 18506 9092 18512 9104
rect 16991 9064 18512 9092
rect 16991 9061 17003 9064
rect 16945 9055 17003 9061
rect 18506 9052 18512 9064
rect 18564 9052 18570 9104
rect 18598 9052 18604 9104
rect 18656 9092 18662 9104
rect 20530 9092 20536 9104
rect 18656 9064 20536 9092
rect 18656 9052 18662 9064
rect 20530 9052 20536 9064
rect 20588 9052 20594 9104
rect 23400 9092 23428 9132
rect 23477 9129 23489 9163
rect 23523 9160 23535 9163
rect 23658 9160 23664 9172
rect 23523 9132 23664 9160
rect 23523 9129 23535 9132
rect 23477 9123 23535 9129
rect 23658 9120 23664 9132
rect 23716 9120 23722 9172
rect 24670 9160 24676 9172
rect 24631 9132 24676 9160
rect 24670 9120 24676 9132
rect 24728 9120 24734 9172
rect 24762 9120 24768 9172
rect 24820 9160 24826 9172
rect 26142 9169 26148 9172
rect 25317 9163 25375 9169
rect 25317 9160 25329 9163
rect 24820 9132 25329 9160
rect 24820 9120 24826 9132
rect 25317 9129 25329 9132
rect 25363 9129 25375 9163
rect 25317 9123 25375 9129
rect 26126 9163 26148 9169
rect 26126 9129 26138 9163
rect 26126 9123 26148 9129
rect 26142 9120 26148 9123
rect 26200 9120 26206 9172
rect 26786 9120 26792 9172
rect 26844 9160 26850 9172
rect 35529 9163 35587 9169
rect 26844 9132 30512 9160
rect 26844 9120 26850 9132
rect 24210 9092 24216 9104
rect 23400 9064 24216 9092
rect 24210 9052 24216 9064
rect 24268 9052 24274 9104
rect 27246 9052 27252 9104
rect 27304 9092 27310 9104
rect 30282 9092 30288 9104
rect 27304 9064 30288 9092
rect 27304 9052 27310 9064
rect 30282 9052 30288 9064
rect 30340 9052 30346 9104
rect 15657 9027 15715 9033
rect 15657 8993 15669 9027
rect 15703 9024 15715 9027
rect 15930 9024 15936 9036
rect 15703 8996 15936 9024
rect 15703 8993 15715 8996
rect 15657 8987 15715 8993
rect 15930 8984 15936 8996
rect 15988 8984 15994 9036
rect 16301 9027 16359 9033
rect 16301 8993 16313 9027
rect 16347 9024 16359 9027
rect 17494 9024 17500 9036
rect 16347 8996 17500 9024
rect 16347 8993 16359 8996
rect 16301 8987 16359 8993
rect 17494 8984 17500 8996
rect 17552 9024 17558 9036
rect 19797 9027 19855 9033
rect 19797 9024 19809 9027
rect 17552 8996 19809 9024
rect 17552 8984 17558 8996
rect 19797 8993 19809 8996
rect 19843 8993 19855 9027
rect 19797 8987 19855 8993
rect 21177 9027 21235 9033
rect 21177 8993 21189 9027
rect 21223 9024 21235 9027
rect 21726 9024 21732 9036
rect 21223 8996 21732 9024
rect 21223 8993 21235 8996
rect 21177 8987 21235 8993
rect 21726 8984 21732 8996
rect 21784 8984 21790 9036
rect 22186 8984 22192 9036
rect 22244 9024 22250 9036
rect 22925 9027 22983 9033
rect 22244 8996 22416 9024
rect 22244 8984 22250 8996
rect 14976 8928 15516 8956
rect 14976 8916 14982 8928
rect 16666 8916 16672 8968
rect 16724 8956 16730 8968
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 16724 8928 16865 8956
rect 16724 8916 16730 8928
rect 16853 8925 16865 8928
rect 16899 8925 16911 8959
rect 16853 8919 16911 8925
rect 17681 8959 17739 8965
rect 17681 8925 17693 8959
rect 17727 8956 17739 8959
rect 17770 8956 17776 8968
rect 17727 8928 17776 8956
rect 17727 8925 17739 8928
rect 17681 8919 17739 8925
rect 17770 8916 17776 8928
rect 17828 8916 17834 8968
rect 20898 8956 20904 8968
rect 20859 8928 20904 8956
rect 20898 8916 20904 8928
rect 20956 8916 20962 8968
rect 22388 8956 22416 8996
rect 22925 8993 22937 9027
rect 22971 9024 22983 9027
rect 23106 9024 23112 9036
rect 22971 8996 23112 9024
rect 22971 8993 22983 8996
rect 22925 8987 22983 8993
rect 23106 8984 23112 8996
rect 23164 8984 23170 9036
rect 23658 8984 23664 9036
rect 23716 9024 23722 9036
rect 23716 8996 24992 9024
rect 23716 8984 23722 8996
rect 23382 8956 23388 8968
rect 22388 8928 23388 8956
rect 23382 8916 23388 8928
rect 23440 8916 23446 8968
rect 24762 8956 24768 8968
rect 24723 8928 24768 8956
rect 24762 8916 24768 8928
rect 24820 8916 24826 8968
rect 24964 8956 24992 8996
rect 25038 8984 25044 9036
rect 25096 9024 25102 9036
rect 26234 9024 26240 9036
rect 25096 8996 26240 9024
rect 25096 8984 25102 8996
rect 25314 8956 25320 8968
rect 24964 8928 25320 8956
rect 25314 8916 25320 8928
rect 25372 8916 25378 8968
rect 25409 8959 25467 8965
rect 25409 8925 25421 8959
rect 25455 8956 25467 8959
rect 25682 8956 25688 8968
rect 25455 8928 25688 8956
rect 25455 8925 25467 8928
rect 25409 8919 25467 8925
rect 25682 8916 25688 8928
rect 25740 8916 25746 8968
rect 25884 8965 25912 8996
rect 26234 8984 26240 8996
rect 26292 8984 26298 9036
rect 29454 9024 29460 9036
rect 27264 8996 29460 9024
rect 25869 8959 25927 8965
rect 25869 8925 25881 8959
rect 25915 8925 25927 8959
rect 27264 8942 27292 8996
rect 29454 8984 29460 8996
rect 29512 8984 29518 9036
rect 30484 9024 30512 9132
rect 35529 9129 35541 9163
rect 35575 9160 35587 9163
rect 36262 9160 36268 9172
rect 35575 9132 36268 9160
rect 35575 9129 35587 9132
rect 35529 9123 35587 9129
rect 36262 9120 36268 9132
rect 36320 9120 36326 9172
rect 31018 9024 31024 9036
rect 30484 8996 31024 9024
rect 31018 8984 31024 8996
rect 31076 8984 31082 9036
rect 27893 8959 27951 8965
rect 25869 8919 25927 8925
rect 27893 8925 27905 8959
rect 27939 8956 27951 8959
rect 27982 8956 27988 8968
rect 27939 8928 27988 8956
rect 27939 8925 27951 8928
rect 27893 8919 27951 8925
rect 27982 8916 27988 8928
rect 28040 8916 28046 8968
rect 31757 8959 31815 8965
rect 31757 8925 31769 8959
rect 31803 8956 31815 8959
rect 32858 8956 32864 8968
rect 31803 8928 32864 8956
rect 31803 8925 31815 8928
rect 31757 8919 31815 8925
rect 32858 8916 32864 8928
rect 32916 8916 32922 8968
rect 1670 8888 1676 8900
rect 1631 8860 1676 8888
rect 1670 8848 1676 8860
rect 1728 8848 1734 8900
rect 15742 8891 15800 8897
rect 15742 8857 15754 8891
rect 15788 8857 15800 8891
rect 15742 8851 15800 8857
rect 14366 8820 14372 8832
rect 14327 8792 14372 8820
rect 14366 8780 14372 8792
rect 14424 8780 14430 8832
rect 15102 8780 15108 8832
rect 15160 8820 15166 8832
rect 15764 8820 15792 8851
rect 15930 8848 15936 8900
rect 15988 8888 15994 8900
rect 17218 8888 17224 8900
rect 15988 8860 17224 8888
rect 15988 8848 15994 8860
rect 17218 8848 17224 8860
rect 17276 8848 17282 8900
rect 18141 8891 18199 8897
rect 18141 8888 18153 8891
rect 17328 8860 18153 8888
rect 15160 8792 15792 8820
rect 15160 8780 15166 8792
rect 15838 8780 15844 8832
rect 15896 8820 15902 8832
rect 17328 8820 17356 8860
rect 18141 8857 18153 8860
rect 18187 8888 18199 8891
rect 18506 8888 18512 8900
rect 18187 8860 18512 8888
rect 18187 8857 18199 8860
rect 18141 8851 18199 8857
rect 18506 8848 18512 8860
rect 18564 8848 18570 8900
rect 18690 8888 18696 8900
rect 18651 8860 18696 8888
rect 18690 8848 18696 8860
rect 18748 8848 18754 8900
rect 18782 8848 18788 8900
rect 18840 8888 18846 8900
rect 18840 8860 18885 8888
rect 18840 8848 18846 8860
rect 19150 8848 19156 8900
rect 19208 8888 19214 8900
rect 19521 8891 19579 8897
rect 19521 8888 19533 8891
rect 19208 8860 19533 8888
rect 19208 8848 19214 8860
rect 19521 8857 19533 8860
rect 19567 8857 19579 8891
rect 19521 8851 19579 8857
rect 19613 8891 19671 8897
rect 19613 8857 19625 8891
rect 19659 8857 19671 8891
rect 19613 8851 19671 8857
rect 15896 8792 17356 8820
rect 17589 8823 17647 8829
rect 15896 8780 15902 8792
rect 17589 8789 17601 8823
rect 17635 8820 17647 8823
rect 19628 8820 19656 8851
rect 19702 8848 19708 8900
rect 19760 8888 19766 8900
rect 23934 8888 23940 8900
rect 19760 8860 21036 8888
rect 22402 8860 23940 8888
rect 19760 8848 19766 8860
rect 17635 8792 19656 8820
rect 21008 8820 21036 8860
rect 23934 8848 23940 8860
rect 23992 8848 23998 8900
rect 24394 8848 24400 8900
rect 24452 8888 24458 8900
rect 26418 8888 26424 8900
rect 24452 8860 26424 8888
rect 24452 8848 24458 8860
rect 26418 8848 26424 8860
rect 26476 8848 26482 8900
rect 27522 8848 27528 8900
rect 27580 8888 27586 8900
rect 29733 8891 29791 8897
rect 29733 8888 29745 8891
rect 27580 8860 29745 8888
rect 27580 8848 27586 8860
rect 29733 8857 29745 8860
rect 29779 8857 29791 8891
rect 29733 8851 29791 8857
rect 31018 8848 31024 8900
rect 31076 8848 31082 8900
rect 31481 8891 31539 8897
rect 31481 8857 31493 8891
rect 31527 8888 31539 8891
rect 31938 8888 31944 8900
rect 31527 8860 31944 8888
rect 31527 8857 31539 8860
rect 31481 8851 31539 8857
rect 31938 8848 31944 8860
rect 31996 8848 32002 8900
rect 34790 8888 34796 8900
rect 32232 8860 34796 8888
rect 23658 8820 23664 8832
rect 21008 8792 23664 8820
rect 17635 8789 17647 8792
rect 17589 8783 17647 8789
rect 23658 8780 23664 8792
rect 23716 8780 23722 8832
rect 23750 8780 23756 8832
rect 23808 8820 23814 8832
rect 26510 8820 26516 8832
rect 23808 8792 26516 8820
rect 23808 8780 23814 8792
rect 26510 8780 26516 8792
rect 26568 8780 26574 8832
rect 27154 8780 27160 8832
rect 27212 8820 27218 8832
rect 28353 8823 28411 8829
rect 28353 8820 28365 8823
rect 27212 8792 28365 8820
rect 27212 8780 27218 8792
rect 28353 8789 28365 8792
rect 28399 8820 28411 8823
rect 28905 8823 28963 8829
rect 28905 8820 28917 8823
rect 28399 8792 28917 8820
rect 28399 8789 28411 8792
rect 28353 8783 28411 8789
rect 28905 8789 28917 8792
rect 28951 8820 28963 8823
rect 29086 8820 29092 8832
rect 28951 8792 29092 8820
rect 28951 8789 28963 8792
rect 28905 8783 28963 8789
rect 29086 8780 29092 8792
rect 29144 8780 29150 8832
rect 29822 8780 29828 8832
rect 29880 8820 29886 8832
rect 32232 8820 32260 8860
rect 34790 8848 34796 8860
rect 34848 8848 34854 8900
rect 35342 8848 35348 8900
rect 35400 8888 35406 8900
rect 35989 8891 36047 8897
rect 35989 8888 36001 8891
rect 35400 8860 36001 8888
rect 35400 8848 35406 8860
rect 35989 8857 36001 8860
rect 36035 8888 36047 8891
rect 38197 8891 38255 8897
rect 38197 8888 38209 8891
rect 36035 8860 38209 8888
rect 36035 8857 36047 8860
rect 35989 8851 36047 8857
rect 38197 8857 38209 8860
rect 38243 8857 38255 8891
rect 38197 8851 38255 8857
rect 29880 8792 32260 8820
rect 32309 8823 32367 8829
rect 29880 8780 29886 8792
rect 32309 8789 32321 8823
rect 32355 8820 32367 8823
rect 32858 8820 32864 8832
rect 32355 8792 32864 8820
rect 32355 8789 32367 8792
rect 32309 8783 32367 8789
rect 32858 8780 32864 8792
rect 32916 8820 32922 8832
rect 33321 8823 33379 8829
rect 33321 8820 33333 8823
rect 32916 8792 33333 8820
rect 32916 8780 32922 8792
rect 33321 8789 33333 8792
rect 33367 8820 33379 8823
rect 33873 8823 33931 8829
rect 33873 8820 33885 8823
rect 33367 8792 33885 8820
rect 33367 8789 33379 8792
rect 33321 8783 33379 8789
rect 33873 8789 33885 8792
rect 33919 8789 33931 8823
rect 33873 8783 33931 8789
rect 34422 8780 34428 8832
rect 34480 8820 34486 8832
rect 34885 8823 34943 8829
rect 34885 8820 34897 8823
rect 34480 8792 34897 8820
rect 34480 8780 34486 8792
rect 34885 8789 34897 8792
rect 34931 8820 34943 8823
rect 35710 8820 35716 8832
rect 34931 8792 35716 8820
rect 34931 8789 34943 8792
rect 34885 8783 34943 8789
rect 35710 8780 35716 8792
rect 35768 8820 35774 8832
rect 36541 8823 36599 8829
rect 36541 8820 36553 8823
rect 35768 8792 36553 8820
rect 35768 8780 35774 8792
rect 36541 8789 36553 8792
rect 36587 8789 36599 8823
rect 36541 8783 36599 8789
rect 37185 8823 37243 8829
rect 37185 8789 37197 8823
rect 37231 8820 37243 8823
rect 37274 8820 37280 8832
rect 37231 8792 37280 8820
rect 37231 8789 37243 8792
rect 37185 8783 37243 8789
rect 37274 8780 37280 8792
rect 37332 8820 37338 8832
rect 37645 8823 37703 8829
rect 37645 8820 37657 8823
rect 37332 8792 37657 8820
rect 37332 8780 37338 8792
rect 37645 8789 37657 8792
rect 37691 8789 37703 8823
rect 37645 8783 37703 8789
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1670 8616 1676 8628
rect 1631 8588 1676 8616
rect 1670 8576 1676 8588
rect 1728 8576 1734 8628
rect 10873 8619 10931 8625
rect 10873 8585 10885 8619
rect 10919 8616 10931 8619
rect 10919 8588 14320 8616
rect 10919 8585 10931 8588
rect 10873 8579 10931 8585
rect 14090 8548 14096 8560
rect 14051 8520 14096 8548
rect 14090 8508 14096 8520
rect 14148 8508 14154 8560
rect 14292 8548 14320 8588
rect 14366 8576 14372 8628
rect 14424 8616 14430 8628
rect 14424 8588 16712 8616
rect 14424 8576 14430 8588
rect 14550 8548 14556 8560
rect 14292 8520 14556 8548
rect 14550 8508 14556 8520
rect 14608 8508 14614 8560
rect 14645 8551 14703 8557
rect 14645 8517 14657 8551
rect 14691 8548 14703 8551
rect 15746 8548 15752 8560
rect 14691 8520 15752 8548
rect 14691 8517 14703 8520
rect 14645 8511 14703 8517
rect 15746 8508 15752 8520
rect 15804 8508 15810 8560
rect 15841 8551 15899 8557
rect 15841 8517 15853 8551
rect 15887 8548 15899 8551
rect 16574 8548 16580 8560
rect 15887 8520 16580 8548
rect 15887 8517 15899 8520
rect 15841 8511 15899 8517
rect 16574 8508 16580 8520
rect 16632 8508 16638 8560
rect 2498 8440 2504 8492
rect 2556 8480 2562 8492
rect 10781 8483 10839 8489
rect 10781 8480 10793 8483
rect 2556 8452 10793 8480
rect 2556 8440 2562 8452
rect 10781 8449 10793 8452
rect 10827 8449 10839 8483
rect 10781 8443 10839 8449
rect 13633 8415 13691 8421
rect 13633 8381 13645 8415
rect 13679 8412 13691 8415
rect 14550 8412 14556 8424
rect 13679 8384 14556 8412
rect 13679 8381 13691 8384
rect 13633 8375 13691 8381
rect 14550 8372 14556 8384
rect 14608 8412 14614 8424
rect 14737 8415 14795 8421
rect 14737 8412 14749 8415
rect 14608 8384 14749 8412
rect 14608 8372 14614 8384
rect 14737 8381 14749 8384
rect 14783 8412 14795 8415
rect 15838 8412 15844 8424
rect 14783 8384 15844 8412
rect 14783 8381 14795 8384
rect 14737 8375 14795 8381
rect 15838 8372 15844 8384
rect 15896 8372 15902 8424
rect 15933 8415 15991 8421
rect 15933 8381 15945 8415
rect 15979 8381 15991 8415
rect 16684 8412 16712 8588
rect 17402 8576 17408 8628
rect 17460 8616 17466 8628
rect 18598 8616 18604 8628
rect 17460 8588 18604 8616
rect 17460 8576 17466 8588
rect 18598 8576 18604 8588
rect 18656 8576 18662 8628
rect 18690 8576 18696 8628
rect 18748 8616 18754 8628
rect 19426 8616 19432 8628
rect 18748 8588 19432 8616
rect 18748 8576 18754 8588
rect 19426 8576 19432 8588
rect 19484 8576 19490 8628
rect 19705 8619 19763 8625
rect 19705 8585 19717 8619
rect 19751 8616 19763 8619
rect 19886 8616 19892 8628
rect 19751 8588 19892 8616
rect 19751 8585 19763 8588
rect 19705 8579 19763 8585
rect 19886 8576 19892 8588
rect 19944 8576 19950 8628
rect 22002 8576 22008 8628
rect 22060 8576 22066 8628
rect 31202 8616 31208 8628
rect 24688 8588 31208 8616
rect 17034 8548 17040 8560
rect 16995 8520 17040 8548
rect 17034 8508 17040 8520
rect 17092 8508 17098 8560
rect 17586 8508 17592 8560
rect 17644 8548 17650 8560
rect 18233 8551 18291 8557
rect 18233 8548 18245 8551
rect 17644 8520 18245 8548
rect 17644 8508 17650 8520
rect 18233 8517 18245 8520
rect 18279 8517 18291 8551
rect 18233 8511 18291 8517
rect 18506 8508 18512 8560
rect 18564 8548 18570 8560
rect 18564 8520 20010 8548
rect 18564 8508 18570 8520
rect 20898 8508 20904 8560
rect 20956 8548 20962 8560
rect 20956 8520 21496 8548
rect 20956 8508 20962 8520
rect 18785 8483 18843 8489
rect 18785 8449 18797 8483
rect 18831 8480 18843 8483
rect 19242 8480 19248 8492
rect 18831 8452 19248 8480
rect 18831 8449 18843 8452
rect 18785 8443 18843 8449
rect 19242 8440 19248 8452
rect 19300 8440 19306 8492
rect 21468 8480 21496 8520
rect 22020 8480 22048 8576
rect 24688 8548 24716 8588
rect 31202 8576 31208 8588
rect 31260 8576 31266 8628
rect 32766 8576 32772 8628
rect 32824 8616 32830 8628
rect 38105 8619 38163 8625
rect 38105 8616 38117 8619
rect 32824 8588 38117 8616
rect 32824 8576 32830 8588
rect 38105 8585 38117 8588
rect 38151 8585 38163 8619
rect 38105 8579 38163 8585
rect 23598 8520 24716 8548
rect 25682 8508 25688 8560
rect 25740 8548 25746 8560
rect 27522 8548 27528 8560
rect 25740 8520 27528 8548
rect 25740 8508 25746 8520
rect 27522 8508 27528 8520
rect 27580 8508 27586 8560
rect 29822 8548 29828 8560
rect 28658 8520 29828 8548
rect 29822 8508 29828 8520
rect 29880 8508 29886 8560
rect 30098 8508 30104 8560
rect 30156 8508 30162 8560
rect 30834 8508 30840 8560
rect 30892 8548 30898 8560
rect 31113 8551 31171 8557
rect 31113 8548 31125 8551
rect 30892 8520 31125 8548
rect 30892 8508 30898 8520
rect 31113 8517 31125 8520
rect 31159 8517 31171 8551
rect 31113 8511 31171 8517
rect 31938 8508 31944 8560
rect 31996 8548 32002 8560
rect 32214 8548 32220 8560
rect 31996 8520 32220 8548
rect 31996 8508 32002 8520
rect 32214 8508 32220 8520
rect 32272 8508 32278 8560
rect 22097 8483 22155 8489
rect 22097 8480 22109 8483
rect 21468 8452 22109 8480
rect 21468 8424 21496 8452
rect 22097 8449 22109 8452
rect 22143 8449 22155 8483
rect 22097 8443 22155 8449
rect 24854 8440 24860 8492
rect 24912 8440 24918 8492
rect 31389 8483 31447 8489
rect 28736 8452 29684 8480
rect 16945 8415 17003 8421
rect 16945 8412 16957 8415
rect 16684 8384 16957 8412
rect 15933 8375 15991 8381
rect 16945 8381 16957 8384
rect 16991 8412 17003 8415
rect 18141 8415 18199 8421
rect 18141 8412 18153 8415
rect 16991 8384 18153 8412
rect 16991 8381 17003 8384
rect 16945 8375 17003 8381
rect 18141 8381 18153 8384
rect 18187 8381 18199 8415
rect 20714 8412 20720 8424
rect 18141 8375 18199 8381
rect 18248 8384 20720 8412
rect 14090 8304 14096 8356
rect 14148 8344 14154 8356
rect 15381 8347 15439 8353
rect 15381 8344 15393 8347
rect 14148 8316 15393 8344
rect 14148 8304 14154 8316
rect 15381 8313 15393 8316
rect 15427 8313 15439 8347
rect 15948 8344 15976 8375
rect 17494 8344 17500 8356
rect 15948 8316 17500 8344
rect 15381 8307 15439 8313
rect 17494 8304 17500 8316
rect 17552 8304 17558 8356
rect 18248 8344 18276 8384
rect 20714 8372 20720 8384
rect 20772 8372 20778 8424
rect 21174 8412 21180 8424
rect 21135 8384 21180 8412
rect 21174 8372 21180 8384
rect 21232 8372 21238 8424
rect 21450 8412 21456 8424
rect 21411 8384 21456 8412
rect 21450 8372 21456 8384
rect 21508 8372 21514 8424
rect 22002 8372 22008 8424
rect 22060 8412 22066 8424
rect 22373 8415 22431 8421
rect 22373 8412 22385 8415
rect 22060 8384 22385 8412
rect 22060 8372 22066 8384
rect 22373 8381 22385 8384
rect 22419 8381 22431 8415
rect 22373 8375 22431 8381
rect 23845 8415 23903 8421
rect 23845 8381 23857 8415
rect 23891 8412 23903 8415
rect 24026 8412 24032 8424
rect 23891 8384 24032 8412
rect 23891 8381 23903 8384
rect 23845 8375 23903 8381
rect 24026 8372 24032 8384
rect 24084 8372 24090 8424
rect 24489 8415 24547 8421
rect 24489 8381 24501 8415
rect 24535 8412 24547 8415
rect 25222 8412 25228 8424
rect 24535 8384 25228 8412
rect 24535 8381 24547 8384
rect 24489 8375 24547 8381
rect 25222 8372 25228 8384
rect 25280 8372 25286 8424
rect 25314 8372 25320 8424
rect 25372 8412 25378 8424
rect 25961 8415 26019 8421
rect 25961 8412 25973 8415
rect 25372 8384 25973 8412
rect 25372 8372 25378 8384
rect 25961 8381 25973 8384
rect 26007 8381 26019 8415
rect 26234 8412 26240 8424
rect 26195 8384 26240 8412
rect 25961 8375 26019 8381
rect 26234 8372 26240 8384
rect 26292 8372 26298 8424
rect 27154 8412 27160 8424
rect 27115 8384 27160 8412
rect 27154 8372 27160 8384
rect 27212 8372 27218 8424
rect 27433 8415 27491 8421
rect 27433 8412 27445 8415
rect 27264 8384 27445 8412
rect 17880 8316 18276 8344
rect 15194 8236 15200 8288
rect 15252 8276 15258 8288
rect 16390 8276 16396 8288
rect 15252 8248 16396 8276
rect 15252 8236 15258 8248
rect 16390 8236 16396 8248
rect 16448 8236 16454 8288
rect 16666 8236 16672 8288
rect 16724 8276 16730 8288
rect 17880 8276 17908 8316
rect 18598 8304 18604 8356
rect 18656 8344 18662 8356
rect 20162 8344 20168 8356
rect 18656 8316 20168 8344
rect 18656 8304 18662 8316
rect 20162 8304 20168 8316
rect 20220 8304 20226 8356
rect 21818 8304 21824 8356
rect 21876 8344 21882 8356
rect 22094 8344 22100 8356
rect 21876 8316 22100 8344
rect 21876 8304 21882 8316
rect 22094 8304 22100 8316
rect 22152 8304 22158 8356
rect 26418 8304 26424 8356
rect 26476 8344 26482 8356
rect 27062 8344 27068 8356
rect 26476 8316 27068 8344
rect 26476 8304 26482 8316
rect 27062 8304 27068 8316
rect 27120 8344 27126 8356
rect 27264 8344 27292 8384
rect 27433 8381 27445 8384
rect 27479 8381 27491 8415
rect 27433 8375 27491 8381
rect 27522 8372 27528 8424
rect 27580 8412 27586 8424
rect 28736 8412 28764 8452
rect 27580 8384 28764 8412
rect 29181 8415 29239 8421
rect 27580 8372 27586 8384
rect 29181 8381 29193 8415
rect 29227 8412 29239 8415
rect 29270 8412 29276 8424
rect 29227 8384 29276 8412
rect 29227 8381 29239 8384
rect 29181 8375 29239 8381
rect 29270 8372 29276 8384
rect 29328 8372 29334 8424
rect 29656 8421 29684 8452
rect 31389 8449 31401 8483
rect 31435 8480 31447 8483
rect 32858 8480 32864 8492
rect 31435 8452 32864 8480
rect 31435 8449 31447 8452
rect 31389 8443 31447 8449
rect 32858 8440 32864 8452
rect 32916 8440 32922 8492
rect 35710 8480 35716 8492
rect 35623 8452 35716 8480
rect 35710 8440 35716 8452
rect 35768 8480 35774 8492
rect 36173 8483 36231 8489
rect 36173 8480 36185 8483
rect 35768 8452 36185 8480
rect 35768 8440 35774 8452
rect 36173 8449 36185 8452
rect 36219 8449 36231 8483
rect 36173 8443 36231 8449
rect 37645 8483 37703 8489
rect 37645 8449 37657 8483
rect 37691 8480 37703 8483
rect 38286 8480 38292 8492
rect 37691 8452 38292 8480
rect 37691 8449 37703 8452
rect 37645 8443 37703 8449
rect 38286 8440 38292 8452
rect 38344 8440 38350 8492
rect 29641 8415 29699 8421
rect 29641 8381 29653 8415
rect 29687 8412 29699 8415
rect 30650 8412 30656 8424
rect 29687 8384 30656 8412
rect 29687 8381 29699 8384
rect 29641 8375 29699 8381
rect 30650 8372 30656 8384
rect 30708 8372 30714 8424
rect 31018 8372 31024 8424
rect 31076 8412 31082 8424
rect 32309 8415 32367 8421
rect 32309 8412 32321 8415
rect 31076 8384 32321 8412
rect 31076 8372 31082 8384
rect 32309 8381 32321 8384
rect 32355 8381 32367 8415
rect 32309 8375 32367 8381
rect 30098 8344 30104 8356
rect 27120 8316 27292 8344
rect 28460 8316 30104 8344
rect 27120 8304 27126 8316
rect 16724 8248 17908 8276
rect 16724 8236 16730 8248
rect 18874 8236 18880 8288
rect 18932 8276 18938 8288
rect 28460 8276 28488 8316
rect 30098 8304 30104 8316
rect 30156 8304 30162 8356
rect 34517 8347 34575 8353
rect 34517 8344 34529 8347
rect 31312 8316 34529 8344
rect 18932 8248 28488 8276
rect 18932 8236 18938 8248
rect 29914 8236 29920 8288
rect 29972 8276 29978 8288
rect 31312 8276 31340 8316
rect 34517 8313 34529 8316
rect 34563 8313 34575 8347
rect 34517 8307 34575 8313
rect 35161 8347 35219 8353
rect 35161 8313 35173 8347
rect 35207 8344 35219 8347
rect 35342 8344 35348 8356
rect 35207 8316 35348 8344
rect 35207 8313 35219 8316
rect 35161 8307 35219 8313
rect 35342 8304 35348 8316
rect 35400 8304 35406 8356
rect 29972 8248 31340 8276
rect 29972 8236 29978 8248
rect 32858 8236 32864 8288
rect 32916 8276 32922 8288
rect 32953 8279 33011 8285
rect 32953 8276 32965 8279
rect 32916 8248 32965 8276
rect 32916 8236 32922 8248
rect 32953 8245 32965 8248
rect 32999 8276 33011 8279
rect 33505 8279 33563 8285
rect 33505 8276 33517 8279
rect 32999 8248 33517 8276
rect 32999 8245 33011 8248
rect 32953 8239 33011 8245
rect 33505 8245 33517 8248
rect 33551 8276 33563 8279
rect 34057 8279 34115 8285
rect 34057 8276 34069 8279
rect 33551 8248 34069 8276
rect 33551 8245 33563 8248
rect 33505 8239 33563 8245
rect 34057 8245 34069 8248
rect 34103 8276 34115 8279
rect 34606 8276 34612 8288
rect 34103 8248 34612 8276
rect 34103 8245 34115 8248
rect 34057 8239 34115 8245
rect 34606 8236 34612 8248
rect 34664 8236 34670 8288
rect 36817 8279 36875 8285
rect 36817 8245 36829 8279
rect 36863 8276 36875 8279
rect 37274 8276 37280 8288
rect 36863 8248 37280 8276
rect 36863 8245 36875 8248
rect 36817 8239 36875 8245
rect 37274 8236 37280 8248
rect 37332 8236 37338 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 16209 8075 16267 8081
rect 16209 8041 16221 8075
rect 16255 8072 16267 8075
rect 17034 8072 17040 8084
rect 16255 8044 17040 8072
rect 16255 8041 16267 8044
rect 16209 8035 16267 8041
rect 17034 8032 17040 8044
rect 17092 8032 17098 8084
rect 17497 8075 17555 8081
rect 17497 8041 17509 8075
rect 17543 8072 17555 8075
rect 17586 8072 17592 8084
rect 17543 8044 17592 8072
rect 17543 8041 17555 8044
rect 17497 8035 17555 8041
rect 17586 8032 17592 8044
rect 17644 8032 17650 8084
rect 18141 8075 18199 8081
rect 18141 8041 18153 8075
rect 18187 8072 18199 8075
rect 18322 8072 18328 8084
rect 18187 8044 18328 8072
rect 18187 8041 18199 8044
rect 18141 8035 18199 8041
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 18785 8075 18843 8081
rect 18785 8041 18797 8075
rect 18831 8072 18843 8075
rect 19334 8072 19340 8084
rect 18831 8044 19340 8072
rect 18831 8041 18843 8044
rect 18785 8035 18843 8041
rect 19334 8032 19340 8044
rect 19392 8032 19398 8084
rect 19797 8075 19855 8081
rect 19797 8041 19809 8075
rect 19843 8072 19855 8075
rect 21634 8072 21640 8084
rect 19843 8044 21640 8072
rect 19843 8041 19855 8044
rect 19797 8035 19855 8041
rect 21634 8032 21640 8044
rect 21692 8032 21698 8084
rect 27414 8075 27472 8081
rect 27414 8072 27426 8075
rect 22940 8044 27426 8072
rect 15657 8007 15715 8013
rect 15657 7973 15669 8007
rect 15703 8004 15715 8007
rect 16666 8004 16672 8016
rect 15703 7976 16672 8004
rect 15703 7973 15715 7976
rect 15657 7967 15715 7973
rect 16666 7964 16672 7976
rect 16724 7964 16730 8016
rect 16853 8007 16911 8013
rect 16853 7973 16865 8007
rect 16899 8004 16911 8007
rect 17218 8004 17224 8016
rect 16899 7976 17224 8004
rect 16899 7973 16911 7976
rect 16853 7967 16911 7973
rect 17218 7964 17224 7976
rect 17276 7964 17282 8016
rect 17954 8004 17960 8016
rect 17328 7976 17960 8004
rect 14642 7936 14648 7948
rect 14603 7908 14648 7936
rect 14642 7896 14648 7908
rect 14700 7896 14706 7948
rect 15010 7896 15016 7948
rect 15068 7936 15074 7948
rect 17328 7936 17356 7976
rect 17954 7964 17960 7976
rect 18012 7964 18018 8016
rect 18690 7964 18696 8016
rect 18748 8004 18754 8016
rect 20806 8004 20812 8016
rect 18748 7976 20812 8004
rect 18748 7964 18754 7976
rect 20806 7964 20812 7976
rect 20864 7964 20870 8016
rect 15068 7908 17356 7936
rect 17604 7908 20024 7936
rect 15068 7896 15074 7908
rect 16132 7877 16160 7908
rect 16117 7871 16175 7877
rect 16117 7837 16129 7871
rect 16163 7837 16175 7871
rect 16942 7868 16948 7880
rect 16903 7840 16948 7868
rect 16117 7831 16175 7837
rect 16942 7828 16948 7840
rect 17000 7828 17006 7880
rect 17604 7877 17632 7908
rect 19996 7880 20024 7908
rect 21358 7896 21364 7948
rect 21416 7936 21422 7948
rect 22940 7936 22968 8044
rect 27414 8041 27426 8044
rect 27460 8072 27472 8075
rect 27460 8044 31340 8072
rect 27460 8041 27472 8044
rect 27414 8035 27472 8041
rect 28626 7964 28632 8016
rect 28684 8004 28690 8016
rect 28905 8007 28963 8013
rect 28905 8004 28917 8007
rect 28684 7976 28917 8004
rect 28684 7964 28690 7976
rect 28905 7973 28917 7976
rect 28951 7973 28963 8007
rect 29730 8004 29736 8016
rect 29691 7976 29736 8004
rect 28905 7967 28963 7973
rect 29730 7964 29736 7976
rect 29788 7964 29794 8016
rect 30285 8007 30343 8013
rect 30285 7973 30297 8007
rect 30331 8004 30343 8007
rect 30558 8004 30564 8016
rect 30331 7976 30564 8004
rect 30331 7973 30343 7976
rect 30285 7967 30343 7973
rect 30558 7964 30564 7976
rect 30616 7964 30622 8016
rect 30374 7936 30380 7948
rect 21416 7908 22968 7936
rect 25976 7908 30380 7936
rect 21416 7896 21422 7908
rect 17589 7871 17647 7877
rect 17589 7837 17601 7871
rect 17635 7837 17647 7871
rect 17589 7831 17647 7837
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7837 18291 7871
rect 18690 7868 18696 7880
rect 18651 7840 18696 7868
rect 18233 7831 18291 7837
rect 14921 7803 14979 7809
rect 14921 7769 14933 7803
rect 14967 7769 14979 7803
rect 14921 7763 14979 7769
rect 15013 7803 15071 7809
rect 15013 7769 15025 7803
rect 15059 7800 15071 7803
rect 18138 7800 18144 7812
rect 15059 7772 18144 7800
rect 15059 7769 15071 7772
rect 15013 7763 15071 7769
rect 14936 7732 14964 7763
rect 18138 7760 18144 7772
rect 18196 7760 18202 7812
rect 18248 7800 18276 7831
rect 18690 7828 18696 7840
rect 18748 7828 18754 7880
rect 19334 7828 19340 7880
rect 19392 7868 19398 7880
rect 19705 7871 19763 7877
rect 19705 7868 19717 7871
rect 19392 7840 19717 7868
rect 19392 7828 19398 7840
rect 19705 7837 19717 7840
rect 19751 7837 19763 7871
rect 19705 7831 19763 7837
rect 19978 7828 19984 7880
rect 20036 7868 20042 7880
rect 20349 7871 20407 7877
rect 20349 7868 20361 7871
rect 20036 7862 20208 7868
rect 20272 7862 20361 7868
rect 20036 7840 20361 7862
rect 20036 7828 20042 7840
rect 20180 7834 20300 7840
rect 20349 7837 20361 7840
rect 20395 7837 20407 7871
rect 20349 7831 20407 7837
rect 20622 7828 20628 7880
rect 20680 7868 20686 7880
rect 20993 7871 21051 7877
rect 20993 7868 21005 7871
rect 20680 7840 21005 7868
rect 20680 7828 20686 7840
rect 20993 7837 21005 7840
rect 21039 7837 21051 7871
rect 20993 7831 21051 7837
rect 23017 7871 23075 7877
rect 23017 7837 23029 7871
rect 23063 7868 23075 7871
rect 24578 7868 24584 7880
rect 23063 7840 24584 7868
rect 23063 7837 23075 7840
rect 23017 7831 23075 7837
rect 24578 7828 24584 7840
rect 24636 7828 24642 7880
rect 25976 7854 26004 7908
rect 30374 7896 30380 7908
rect 30432 7896 30438 7948
rect 31312 7936 31340 8044
rect 31662 8032 31668 8084
rect 31720 8072 31726 8084
rect 32585 8075 32643 8081
rect 32585 8072 32597 8075
rect 31720 8044 32597 8072
rect 31720 8032 31726 8044
rect 32585 8041 32597 8044
rect 32631 8072 32643 8075
rect 33137 8075 33195 8081
rect 33137 8072 33149 8075
rect 32631 8044 33149 8072
rect 32631 8041 32643 8044
rect 32585 8035 32643 8041
rect 33137 8041 33149 8044
rect 33183 8072 33195 8075
rect 33689 8075 33747 8081
rect 33689 8072 33701 8075
rect 33183 8044 33701 8072
rect 33183 8041 33195 8044
rect 33137 8035 33195 8041
rect 33689 8041 33701 8044
rect 33735 8072 33747 8075
rect 34241 8075 34299 8081
rect 34241 8072 34253 8075
rect 33735 8044 34253 8072
rect 33735 8041 33747 8044
rect 33689 8035 33747 8041
rect 34241 8041 34253 8044
rect 34287 8072 34299 8075
rect 34606 8072 34612 8084
rect 34287 8044 34612 8072
rect 34287 8041 34299 8044
rect 34241 8035 34299 8041
rect 34606 8032 34612 8044
rect 34664 8072 34670 8084
rect 34885 8075 34943 8081
rect 34885 8072 34897 8075
rect 34664 8044 34897 8072
rect 34664 8032 34670 8044
rect 34885 8041 34897 8044
rect 34931 8041 34943 8075
rect 34885 8035 34943 8041
rect 35529 8075 35587 8081
rect 35529 8041 35541 8075
rect 35575 8072 35587 8075
rect 36262 8072 36268 8084
rect 35575 8044 36268 8072
rect 35575 8041 35587 8044
rect 35529 8035 35587 8041
rect 36262 8032 36268 8044
rect 36320 8072 36326 8084
rect 36541 8075 36599 8081
rect 36541 8072 36553 8075
rect 36320 8044 36553 8072
rect 36320 8032 36326 8044
rect 36541 8041 36553 8044
rect 36587 8072 36599 8075
rect 37182 8072 37188 8084
rect 36587 8044 37188 8072
rect 36587 8041 36599 8044
rect 36541 8035 36599 8041
rect 37182 8032 37188 8044
rect 37240 8072 37246 8084
rect 37645 8075 37703 8081
rect 37645 8072 37657 8075
rect 37240 8044 37657 8072
rect 37240 8032 37246 8044
rect 37645 8041 37657 8044
rect 37691 8072 37703 8075
rect 38197 8075 38255 8081
rect 38197 8072 38209 8075
rect 37691 8044 38209 8072
rect 37691 8041 37703 8044
rect 37645 8035 37703 8041
rect 38197 8041 38209 8044
rect 38243 8041 38255 8075
rect 38197 8035 38255 8041
rect 31941 7939 31999 7945
rect 31941 7936 31953 7939
rect 31312 7908 31953 7936
rect 31941 7905 31953 7908
rect 31987 7905 31999 7939
rect 31941 7899 31999 7905
rect 27154 7868 27160 7880
rect 27115 7840 27160 7868
rect 27154 7828 27160 7840
rect 27212 7828 27218 7880
rect 30282 7828 30288 7880
rect 30340 7868 30346 7880
rect 30837 7871 30895 7877
rect 30837 7868 30849 7871
rect 30340 7840 30849 7868
rect 30340 7828 30346 7840
rect 30837 7837 30849 7840
rect 30883 7868 30895 7871
rect 31389 7871 31447 7877
rect 31389 7868 31401 7871
rect 30883 7840 31401 7868
rect 30883 7837 30895 7840
rect 30837 7831 30895 7837
rect 31389 7837 31401 7840
rect 31435 7837 31447 7871
rect 35618 7868 35624 7880
rect 31389 7831 31447 7837
rect 31496 7840 35624 7868
rect 20806 7800 20812 7812
rect 18248 7772 20812 7800
rect 20806 7760 20812 7772
rect 20864 7760 20870 7812
rect 20898 7760 20904 7812
rect 20956 7800 20962 7812
rect 20956 7772 21574 7800
rect 20956 7760 20962 7772
rect 22462 7760 22468 7812
rect 22520 7800 22526 7812
rect 22741 7803 22799 7809
rect 22741 7800 22753 7803
rect 22520 7772 22753 7800
rect 22520 7760 22526 7772
rect 22741 7769 22753 7772
rect 22787 7800 22799 7803
rect 23106 7800 23112 7812
rect 22787 7772 23112 7800
rect 22787 7769 22799 7772
rect 22741 7763 22799 7769
rect 23106 7760 23112 7772
rect 23164 7760 23170 7812
rect 23566 7760 23572 7812
rect 23624 7800 23630 7812
rect 24762 7800 24768 7812
rect 23624 7772 24768 7800
rect 23624 7760 23630 7772
rect 24762 7760 24768 7772
rect 24820 7800 24826 7812
rect 24857 7803 24915 7809
rect 24857 7800 24869 7803
rect 24820 7772 24869 7800
rect 24820 7760 24826 7772
rect 24857 7769 24869 7772
rect 24903 7769 24915 7803
rect 31496 7800 31524 7840
rect 35618 7828 35624 7840
rect 35676 7828 35682 7880
rect 33042 7800 33048 7812
rect 28658 7772 31524 7800
rect 31726 7772 33048 7800
rect 24857 7763 24915 7769
rect 15470 7732 15476 7744
rect 14936 7704 15476 7732
rect 15470 7692 15476 7704
rect 15528 7692 15534 7744
rect 18046 7692 18052 7744
rect 18104 7732 18110 7744
rect 20254 7732 20260 7744
rect 18104 7704 20260 7732
rect 18104 7692 18110 7704
rect 20254 7692 20260 7704
rect 20312 7692 20318 7744
rect 20441 7735 20499 7741
rect 20441 7701 20453 7735
rect 20487 7732 20499 7735
rect 23198 7732 23204 7744
rect 20487 7704 23204 7732
rect 20487 7701 20499 7704
rect 20441 7695 20499 7701
rect 23198 7692 23204 7704
rect 23256 7692 23262 7744
rect 23382 7692 23388 7744
rect 23440 7732 23446 7744
rect 23477 7735 23535 7741
rect 23477 7732 23489 7735
rect 23440 7704 23489 7732
rect 23440 7692 23446 7704
rect 23477 7701 23489 7704
rect 23523 7701 23535 7735
rect 23477 7695 23535 7701
rect 24302 7692 24308 7744
rect 24360 7732 24366 7744
rect 26329 7735 26387 7741
rect 26329 7732 26341 7735
rect 24360 7704 26341 7732
rect 24360 7692 24366 7704
rect 26329 7701 26341 7704
rect 26375 7732 26387 7735
rect 27246 7732 27252 7744
rect 26375 7704 27252 7732
rect 26375 7701 26387 7704
rect 26329 7695 26387 7701
rect 27246 7692 27252 7704
rect 27304 7692 27310 7744
rect 27614 7692 27620 7744
rect 27672 7732 27678 7744
rect 28994 7732 29000 7744
rect 27672 7704 29000 7732
rect 27672 7692 27678 7704
rect 28994 7692 29000 7704
rect 29052 7692 29058 7744
rect 30374 7692 30380 7744
rect 30432 7732 30438 7744
rect 31726 7732 31754 7772
rect 33042 7760 33048 7772
rect 33100 7760 33106 7812
rect 30432 7704 31754 7732
rect 30432 7692 30438 7704
rect 33778 7692 33784 7744
rect 33836 7732 33842 7744
rect 35989 7735 36047 7741
rect 35989 7732 36001 7735
rect 33836 7704 36001 7732
rect 33836 7692 33842 7704
rect 35989 7701 36001 7704
rect 36035 7701 36047 7735
rect 35989 7695 36047 7701
rect 37185 7735 37243 7741
rect 37185 7701 37197 7735
rect 37231 7732 37243 7735
rect 37274 7732 37280 7744
rect 37231 7704 37280 7732
rect 37231 7701 37243 7704
rect 37185 7695 37243 7701
rect 37274 7692 37280 7704
rect 37332 7692 37338 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 13630 7488 13636 7540
rect 13688 7528 13694 7540
rect 13725 7531 13783 7537
rect 13725 7528 13737 7531
rect 13688 7500 13737 7528
rect 13688 7488 13694 7500
rect 13725 7497 13737 7500
rect 13771 7497 13783 7531
rect 15010 7528 15016 7540
rect 14971 7500 15016 7528
rect 13725 7491 13783 7497
rect 15010 7488 15016 7500
rect 15068 7488 15074 7540
rect 17696 7500 17908 7528
rect 14182 7420 14188 7472
rect 14240 7460 14246 7472
rect 15565 7463 15623 7469
rect 15565 7460 15577 7463
rect 14240 7432 15577 7460
rect 14240 7420 14246 7432
rect 15565 7429 15577 7432
rect 15611 7429 15623 7463
rect 15565 7423 15623 7429
rect 16117 7463 16175 7469
rect 16117 7429 16129 7463
rect 16163 7460 16175 7463
rect 17218 7460 17224 7472
rect 16163 7432 17224 7460
rect 16163 7429 16175 7432
rect 16117 7423 16175 7429
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7392 1915 7395
rect 2498 7392 2504 7404
rect 1903 7364 2360 7392
rect 2459 7364 2504 7392
rect 1903 7361 1915 7364
rect 1857 7355 1915 7361
rect 2332 7265 2360 7364
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 10042 7352 10048 7404
rect 10100 7392 10106 7404
rect 13633 7395 13691 7401
rect 13633 7392 13645 7395
rect 10100 7364 13645 7392
rect 10100 7352 10106 7364
rect 13633 7361 13645 7364
rect 13679 7361 13691 7395
rect 13633 7355 13691 7361
rect 2317 7259 2375 7265
rect 2317 7225 2329 7259
rect 2363 7225 2375 7259
rect 15580 7256 15608 7423
rect 17218 7420 17224 7432
rect 17276 7420 17282 7472
rect 17402 7460 17408 7472
rect 17363 7432 17408 7460
rect 17402 7420 17408 7432
rect 17460 7420 17466 7472
rect 17497 7463 17555 7469
rect 17497 7429 17509 7463
rect 17543 7460 17555 7463
rect 17696 7460 17724 7500
rect 17543 7432 17724 7460
rect 17880 7460 17908 7500
rect 17954 7488 17960 7540
rect 18012 7528 18018 7540
rect 18322 7528 18328 7540
rect 18012 7500 18328 7528
rect 18012 7488 18018 7500
rect 18322 7488 18328 7500
rect 18380 7488 18386 7540
rect 18601 7531 18659 7537
rect 18601 7497 18613 7531
rect 18647 7528 18659 7531
rect 18782 7528 18788 7540
rect 18647 7500 18788 7528
rect 18647 7497 18659 7500
rect 18601 7491 18659 7497
rect 18782 7488 18788 7500
rect 18840 7488 18846 7540
rect 19150 7528 19156 7540
rect 19111 7500 19156 7528
rect 19150 7488 19156 7500
rect 19208 7488 19214 7540
rect 19352 7500 22692 7528
rect 19242 7460 19248 7472
rect 17880 7432 19248 7460
rect 17543 7429 17555 7432
rect 17497 7423 17555 7429
rect 19242 7420 19248 7432
rect 19300 7420 19306 7472
rect 16758 7392 16764 7404
rect 16592 7364 16764 7392
rect 16209 7327 16267 7333
rect 16209 7293 16221 7327
rect 16255 7324 16267 7327
rect 16592 7324 16620 7364
rect 16758 7352 16764 7364
rect 16816 7352 16822 7404
rect 19058 7392 19064 7404
rect 19019 7364 19064 7392
rect 19058 7352 19064 7364
rect 19116 7352 19122 7404
rect 16255 7296 16620 7324
rect 16255 7293 16267 7296
rect 16209 7287 16267 7293
rect 16666 7284 16672 7336
rect 16724 7324 16730 7336
rect 19352 7324 19380 7500
rect 21177 7463 21235 7469
rect 21177 7429 21189 7463
rect 21223 7460 21235 7463
rect 22186 7460 22192 7472
rect 21223 7432 22192 7460
rect 21223 7429 21235 7432
rect 21177 7423 21235 7429
rect 22186 7420 22192 7432
rect 22244 7420 22250 7472
rect 22664 7460 22692 7500
rect 22922 7488 22928 7540
rect 22980 7528 22986 7540
rect 24489 7531 24547 7537
rect 24489 7528 24501 7531
rect 22980 7500 24501 7528
rect 22980 7488 22986 7500
rect 24489 7497 24501 7500
rect 24535 7528 24547 7531
rect 24535 7500 26096 7528
rect 24535 7497 24547 7500
rect 24489 7491 24547 7497
rect 22664 7432 22770 7460
rect 24946 7420 24952 7472
rect 25004 7420 25010 7472
rect 25958 7460 25964 7472
rect 25919 7432 25964 7460
rect 25958 7420 25964 7432
rect 26016 7420 26022 7472
rect 26068 7460 26096 7500
rect 27062 7488 27068 7540
rect 27120 7528 27126 7540
rect 28905 7531 28963 7537
rect 27120 7500 28764 7528
rect 27120 7488 27126 7500
rect 27338 7460 27344 7472
rect 26068 7432 27344 7460
rect 27338 7420 27344 7432
rect 27396 7420 27402 7472
rect 28736 7460 28764 7500
rect 28905 7497 28917 7531
rect 28951 7528 28963 7531
rect 29546 7528 29552 7540
rect 28951 7500 29552 7528
rect 28951 7497 28963 7500
rect 28905 7491 28963 7497
rect 29546 7488 29552 7500
rect 29604 7488 29610 7540
rect 29822 7488 29828 7540
rect 29880 7528 29886 7540
rect 31110 7528 31116 7540
rect 29880 7500 31116 7528
rect 29880 7488 29886 7500
rect 31110 7488 31116 7500
rect 31168 7488 31174 7540
rect 31662 7488 31668 7540
rect 31720 7528 31726 7540
rect 32401 7531 32459 7537
rect 32401 7528 32413 7531
rect 31720 7500 32413 7528
rect 31720 7488 31726 7500
rect 32401 7497 32413 7500
rect 32447 7528 32459 7531
rect 33505 7531 33563 7537
rect 33505 7528 33517 7531
rect 32447 7500 33517 7528
rect 32447 7497 32459 7500
rect 32401 7491 32459 7497
rect 33505 7497 33517 7500
rect 33551 7528 33563 7531
rect 34057 7531 34115 7537
rect 34057 7528 34069 7531
rect 33551 7500 34069 7528
rect 33551 7497 33563 7500
rect 33505 7491 33563 7497
rect 34057 7497 34069 7500
rect 34103 7528 34115 7531
rect 34609 7531 34667 7537
rect 34609 7528 34621 7531
rect 34103 7500 34621 7528
rect 34103 7497 34115 7500
rect 34057 7491 34115 7497
rect 34609 7497 34621 7500
rect 34655 7528 34667 7531
rect 35161 7531 35219 7537
rect 35161 7528 35173 7531
rect 34655 7500 35173 7528
rect 34655 7497 34667 7500
rect 34609 7491 34667 7497
rect 35161 7497 35173 7500
rect 35207 7528 35219 7531
rect 35710 7528 35716 7540
rect 35207 7500 35716 7528
rect 35207 7497 35219 7500
rect 35161 7491 35219 7497
rect 35710 7488 35716 7500
rect 35768 7488 35774 7540
rect 37182 7488 37188 7540
rect 37240 7528 37246 7540
rect 37461 7531 37519 7537
rect 37461 7528 37473 7531
rect 37240 7500 37473 7528
rect 37240 7488 37246 7500
rect 37461 7497 37473 7500
rect 37507 7497 37519 7531
rect 37461 7491 37519 7497
rect 30561 7463 30619 7469
rect 30561 7460 30573 7463
rect 28736 7432 30573 7460
rect 30561 7429 30573 7432
rect 30607 7429 30619 7463
rect 30561 7423 30619 7429
rect 32950 7420 32956 7472
rect 33008 7460 33014 7472
rect 36725 7463 36783 7469
rect 36725 7460 36737 7463
rect 33008 7432 36737 7460
rect 33008 7420 33014 7432
rect 36725 7429 36737 7432
rect 36771 7429 36783 7463
rect 36725 7423 36783 7429
rect 20070 7352 20076 7404
rect 20128 7352 20134 7404
rect 21450 7352 21456 7404
rect 21508 7392 21514 7404
rect 21634 7392 21640 7404
rect 21508 7364 21640 7392
rect 21508 7352 21514 7364
rect 21634 7352 21640 7364
rect 21692 7392 21698 7404
rect 22005 7395 22063 7401
rect 22005 7392 22017 7395
rect 21692 7364 22017 7392
rect 21692 7352 21698 7364
rect 22005 7361 22017 7364
rect 22051 7361 22063 7395
rect 22005 7355 22063 7361
rect 26234 7352 26240 7404
rect 26292 7392 26298 7404
rect 26292 7364 27200 7392
rect 26292 7352 26298 7364
rect 27172 7336 27200 7364
rect 16724 7296 19380 7324
rect 16724 7284 16730 7296
rect 20622 7284 20628 7336
rect 20680 7324 20686 7336
rect 22281 7327 22339 7333
rect 22281 7324 22293 7327
rect 20680 7296 22293 7324
rect 20680 7284 20686 7296
rect 22281 7293 22293 7296
rect 22327 7293 22339 7327
rect 22281 7287 22339 7293
rect 22370 7284 22376 7336
rect 22428 7324 22434 7336
rect 23753 7327 23811 7333
rect 23753 7324 23765 7327
rect 22428 7296 23765 7324
rect 22428 7284 22434 7296
rect 23753 7293 23765 7296
rect 23799 7324 23811 7327
rect 25866 7324 25872 7336
rect 23799 7296 25872 7324
rect 23799 7293 23811 7296
rect 23753 7287 23811 7293
rect 25866 7284 25872 7296
rect 25924 7284 25930 7336
rect 26326 7284 26332 7336
rect 26384 7324 26390 7336
rect 26694 7324 26700 7336
rect 26384 7296 26700 7324
rect 26384 7284 26390 7296
rect 26694 7284 26700 7296
rect 26752 7284 26758 7336
rect 27154 7324 27160 7336
rect 27115 7296 27160 7324
rect 27154 7284 27160 7296
rect 27212 7284 27218 7336
rect 27433 7327 27491 7333
rect 27433 7293 27445 7327
rect 27479 7324 27491 7327
rect 28552 7324 28580 7378
rect 28994 7352 29000 7404
rect 29052 7392 29058 7404
rect 30006 7392 30012 7404
rect 29052 7364 30012 7392
rect 29052 7352 29058 7364
rect 30006 7352 30012 7364
rect 30064 7352 30070 7404
rect 36817 7395 36875 7401
rect 36817 7361 36829 7395
rect 36863 7392 36875 7395
rect 37274 7392 37280 7404
rect 36863 7364 37280 7392
rect 36863 7361 36875 7364
rect 36817 7355 36875 7361
rect 37274 7352 37280 7364
rect 37332 7352 37338 7404
rect 31018 7324 31024 7336
rect 27479 7296 28488 7324
rect 28552 7296 31024 7324
rect 27479 7293 27491 7296
rect 27433 7287 27491 7293
rect 16945 7259 17003 7265
rect 16945 7256 16957 7259
rect 15580 7228 16957 7256
rect 2317 7219 2375 7225
rect 16945 7225 16957 7228
rect 16991 7256 17003 7259
rect 17126 7256 17132 7268
rect 16991 7228 17132 7256
rect 16991 7225 17003 7228
rect 16945 7219 17003 7225
rect 17126 7216 17132 7228
rect 17184 7216 17190 7268
rect 17310 7216 17316 7268
rect 17368 7256 17374 7268
rect 28460 7256 28488 7296
rect 31018 7284 31024 7296
rect 31076 7284 31082 7336
rect 28626 7256 28632 7268
rect 17368 7228 20116 7256
rect 28460 7228 28632 7256
rect 17368 7216 17374 7228
rect 1670 7188 1676 7200
rect 1631 7160 1676 7188
rect 1670 7148 1676 7160
rect 1728 7148 1734 7200
rect 15562 7148 15568 7200
rect 15620 7188 15626 7200
rect 18782 7188 18788 7200
rect 15620 7160 18788 7188
rect 15620 7148 15626 7160
rect 18782 7148 18788 7160
rect 18840 7148 18846 7200
rect 19705 7191 19763 7197
rect 19705 7157 19717 7191
rect 19751 7188 19763 7191
rect 19978 7188 19984 7200
rect 19751 7160 19984 7188
rect 19751 7157 19763 7160
rect 19705 7151 19763 7157
rect 19978 7148 19984 7160
rect 20036 7148 20042 7200
rect 20088 7188 20116 7228
rect 28626 7216 28632 7228
rect 28684 7216 28690 7268
rect 28902 7216 28908 7268
rect 28960 7256 28966 7268
rect 29457 7259 29515 7265
rect 29457 7256 29469 7259
rect 28960 7228 29469 7256
rect 28960 7216 28966 7228
rect 29457 7225 29469 7228
rect 29503 7256 29515 7259
rect 30190 7256 30196 7268
rect 29503 7228 30196 7256
rect 29503 7225 29515 7228
rect 29457 7219 29515 7225
rect 30190 7216 30196 7228
rect 30248 7216 30254 7268
rect 31113 7259 31171 7265
rect 31113 7225 31125 7259
rect 31159 7225 31171 7259
rect 31113 7219 31171 7225
rect 21910 7188 21916 7200
rect 20088 7160 21916 7188
rect 21910 7148 21916 7160
rect 21968 7148 21974 7200
rect 22094 7148 22100 7200
rect 22152 7188 22158 7200
rect 22646 7188 22652 7200
rect 22152 7160 22652 7188
rect 22152 7148 22158 7160
rect 22646 7148 22652 7160
rect 22704 7188 22710 7200
rect 23382 7188 23388 7200
rect 22704 7160 23388 7188
rect 22704 7148 22710 7160
rect 23382 7148 23388 7160
rect 23440 7148 23446 7200
rect 25222 7148 25228 7200
rect 25280 7188 25286 7200
rect 29270 7188 29276 7200
rect 25280 7160 29276 7188
rect 25280 7148 25286 7160
rect 29270 7148 29276 7160
rect 29328 7148 29334 7200
rect 29730 7148 29736 7200
rect 29788 7188 29794 7200
rect 30009 7191 30067 7197
rect 30009 7188 30021 7191
rect 29788 7160 30021 7188
rect 29788 7148 29794 7160
rect 30009 7157 30021 7160
rect 30055 7188 30067 7191
rect 30282 7188 30288 7200
rect 30055 7160 30288 7188
rect 30055 7157 30067 7160
rect 30009 7151 30067 7157
rect 30282 7148 30288 7160
rect 30340 7188 30346 7200
rect 31128 7188 31156 7219
rect 31662 7188 31668 7200
rect 30340 7160 31668 7188
rect 30340 7148 30346 7160
rect 31662 7148 31668 7160
rect 31720 7148 31726 7200
rect 32858 7188 32864 7200
rect 32819 7160 32864 7188
rect 32858 7148 32864 7160
rect 32916 7148 32922 7200
rect 38010 7188 38016 7200
rect 37971 7160 38016 7188
rect 38010 7148 38016 7160
rect 38068 7148 38074 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 16040 6956 18644 6984
rect 15286 6848 15292 6860
rect 15247 6820 15292 6848
rect 15286 6808 15292 6820
rect 15344 6808 15350 6860
rect 15746 6808 15752 6860
rect 15804 6848 15810 6860
rect 15933 6851 15991 6857
rect 15933 6848 15945 6851
rect 15804 6820 15945 6848
rect 15804 6808 15810 6820
rect 15933 6817 15945 6820
rect 15979 6817 15991 6851
rect 15933 6811 15991 6817
rect 6362 6780 6368 6792
rect 6323 6752 6368 6780
rect 6362 6740 6368 6752
rect 6420 6780 6426 6792
rect 16040 6789 16068 6956
rect 17310 6876 17316 6928
rect 17368 6916 17374 6928
rect 18230 6916 18236 6928
rect 17368 6888 18236 6916
rect 17368 6876 17374 6888
rect 18230 6876 18236 6888
rect 18288 6876 18294 6928
rect 16574 6848 16580 6860
rect 16535 6820 16580 6848
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 18414 6848 18420 6860
rect 16684 6820 18276 6848
rect 18375 6820 18420 6848
rect 16684 6789 16712 6820
rect 7009 6783 7067 6789
rect 7009 6780 7021 6783
rect 6420 6752 7021 6780
rect 6420 6740 6426 6752
rect 7009 6749 7021 6752
rect 7055 6749 7067 6783
rect 7009 6743 7067 6749
rect 16025 6783 16083 6789
rect 16025 6749 16037 6783
rect 16071 6749 16083 6783
rect 16025 6743 16083 6749
rect 16669 6783 16727 6789
rect 16669 6749 16681 6783
rect 16715 6749 16727 6783
rect 16669 6743 16727 6749
rect 17313 6783 17371 6789
rect 17313 6749 17325 6783
rect 17359 6780 17371 6783
rect 18138 6780 18144 6792
rect 17359 6752 18144 6780
rect 17359 6749 17371 6752
rect 17313 6743 17371 6749
rect 18138 6740 18144 6752
rect 18196 6740 18202 6792
rect 18248 6780 18276 6820
rect 18414 6808 18420 6820
rect 18472 6808 18478 6860
rect 18616 6848 18644 6956
rect 18782 6944 18788 6996
rect 18840 6984 18846 6996
rect 23290 6984 23296 6996
rect 18840 6956 23296 6984
rect 18840 6944 18846 6956
rect 23290 6944 23296 6956
rect 23348 6944 23354 6996
rect 26050 6944 26056 6996
rect 26108 6984 26114 6996
rect 27249 6987 27307 6993
rect 27249 6984 27261 6987
rect 26108 6956 27261 6984
rect 26108 6944 26114 6956
rect 27249 6953 27261 6956
rect 27295 6953 27307 6987
rect 27249 6947 27307 6953
rect 28739 6987 28797 6993
rect 28739 6953 28751 6987
rect 28785 6984 28797 6987
rect 28994 6984 29000 6996
rect 28785 6956 29000 6984
rect 28785 6953 28797 6956
rect 28739 6947 28797 6953
rect 28994 6944 29000 6956
rect 29052 6944 29058 6996
rect 29546 6944 29552 6996
rect 29604 6984 29610 6996
rect 29990 6987 30048 6993
rect 29990 6984 30002 6987
rect 29604 6956 30002 6984
rect 29604 6944 29610 6956
rect 29990 6953 30002 6956
rect 30036 6953 30048 6987
rect 29990 6947 30048 6953
rect 30742 6944 30748 6996
rect 30800 6984 30806 6996
rect 31481 6987 31539 6993
rect 31481 6984 31493 6987
rect 30800 6956 31493 6984
rect 30800 6944 30806 6956
rect 31481 6953 31493 6956
rect 31527 6953 31539 6987
rect 31481 6947 31539 6953
rect 31754 6944 31760 6996
rect 31812 6984 31818 6996
rect 33686 6984 33692 6996
rect 31812 6956 33692 6984
rect 31812 6944 31818 6956
rect 33686 6944 33692 6956
rect 33744 6944 33750 6996
rect 19150 6876 19156 6928
rect 19208 6916 19214 6928
rect 20070 6916 20076 6928
rect 19208 6888 20076 6916
rect 19208 6876 19214 6888
rect 20070 6876 20076 6888
rect 20128 6876 20134 6928
rect 22370 6876 22376 6928
rect 22428 6916 22434 6928
rect 25130 6916 25136 6928
rect 22428 6888 25136 6916
rect 22428 6876 22434 6888
rect 25130 6876 25136 6888
rect 25188 6876 25194 6928
rect 31202 6876 31208 6928
rect 31260 6916 31266 6928
rect 33318 6916 33324 6928
rect 31260 6888 33324 6916
rect 31260 6876 31266 6888
rect 33318 6876 33324 6888
rect 33376 6876 33382 6928
rect 18616 6820 18920 6848
rect 18509 6783 18567 6789
rect 18248 6752 18368 6780
rect 14642 6712 14648 6724
rect 14603 6684 14648 6712
rect 14642 6672 14648 6684
rect 14700 6672 14706 6724
rect 15197 6715 15255 6721
rect 15197 6681 15209 6715
rect 15243 6712 15255 6715
rect 15838 6712 15844 6724
rect 15243 6684 15844 6712
rect 15243 6681 15255 6684
rect 15197 6675 15255 6681
rect 15838 6672 15844 6684
rect 15896 6672 15902 6724
rect 16482 6672 16488 6724
rect 16540 6712 16546 6724
rect 17221 6715 17279 6721
rect 17221 6712 17233 6715
rect 16540 6684 17233 6712
rect 16540 6672 16546 6684
rect 17221 6681 17233 6684
rect 17267 6681 17279 6715
rect 17770 6712 17776 6724
rect 17731 6684 17776 6712
rect 17221 6675 17279 6681
rect 17770 6672 17776 6684
rect 17828 6672 17834 6724
rect 6546 6644 6552 6656
rect 6507 6616 6552 6644
rect 6546 6604 6552 6616
rect 6604 6604 6610 6656
rect 18340 6644 18368 6752
rect 18509 6749 18521 6783
rect 18555 6780 18567 6783
rect 18782 6780 18788 6792
rect 18555 6752 18788 6780
rect 18555 6749 18567 6752
rect 18509 6743 18567 6749
rect 18782 6740 18788 6752
rect 18840 6740 18846 6792
rect 18892 6712 18920 6820
rect 19426 6808 19432 6860
rect 19484 6848 19490 6860
rect 19521 6851 19579 6857
rect 19521 6848 19533 6851
rect 19484 6820 19533 6848
rect 19484 6808 19490 6820
rect 19521 6817 19533 6820
rect 19567 6817 19579 6851
rect 20254 6848 20260 6860
rect 19521 6811 19579 6817
rect 19628 6820 20260 6848
rect 19242 6740 19248 6792
rect 19300 6780 19306 6792
rect 19628 6789 19656 6820
rect 20254 6808 20260 6820
rect 20312 6808 20318 6860
rect 20349 6851 20407 6857
rect 20349 6817 20361 6851
rect 20395 6848 20407 6851
rect 21726 6848 21732 6860
rect 20395 6820 21732 6848
rect 20395 6817 20407 6820
rect 20349 6811 20407 6817
rect 21726 6808 21732 6820
rect 21784 6808 21790 6860
rect 22554 6808 22560 6860
rect 22612 6848 22618 6860
rect 22833 6851 22891 6857
rect 22833 6848 22845 6851
rect 22612 6820 22845 6848
rect 22612 6808 22618 6820
rect 22833 6817 22845 6820
rect 22879 6817 22891 6851
rect 22833 6811 22891 6817
rect 24394 6808 24400 6860
rect 24452 6848 24458 6860
rect 24765 6851 24823 6857
rect 24765 6848 24777 6851
rect 24452 6820 24777 6848
rect 24452 6808 24458 6820
rect 24765 6817 24777 6820
rect 24811 6817 24823 6851
rect 25148 6848 25176 6876
rect 26142 6848 26148 6860
rect 25148 6820 26148 6848
rect 24765 6811 24823 6817
rect 26142 6808 26148 6820
rect 26200 6808 26206 6860
rect 27338 6808 27344 6860
rect 27396 6848 27402 6860
rect 30558 6848 30564 6860
rect 27396 6820 30564 6848
rect 27396 6808 27402 6820
rect 30558 6808 30564 6820
rect 30616 6808 30622 6860
rect 36541 6851 36599 6857
rect 36541 6848 36553 6851
rect 31128 6820 36553 6848
rect 19613 6783 19671 6789
rect 19613 6780 19625 6783
rect 19300 6752 19625 6780
rect 19300 6740 19306 6752
rect 19613 6749 19625 6752
rect 19659 6749 19671 6783
rect 19613 6743 19671 6749
rect 19702 6740 19708 6792
rect 19760 6780 19766 6792
rect 22373 6783 22431 6789
rect 19760 6752 21022 6780
rect 19760 6740 19766 6752
rect 22373 6749 22385 6783
rect 22419 6780 22431 6783
rect 22462 6780 22468 6792
rect 22419 6752 22468 6780
rect 22419 6749 22431 6752
rect 22373 6743 22431 6749
rect 22462 6740 22468 6752
rect 22520 6780 22526 6792
rect 23385 6783 23443 6789
rect 23385 6780 23397 6783
rect 22520 6752 23397 6780
rect 22520 6740 22526 6752
rect 23385 6749 23397 6752
rect 23431 6749 23443 6783
rect 23385 6743 23443 6749
rect 26513 6783 26571 6789
rect 26513 6749 26525 6783
rect 26559 6780 26571 6783
rect 27154 6780 27160 6792
rect 26559 6752 27160 6780
rect 26559 6749 26571 6752
rect 26513 6743 26571 6749
rect 27154 6740 27160 6752
rect 27212 6740 27218 6792
rect 28994 6740 29000 6792
rect 29052 6780 29058 6792
rect 29730 6780 29736 6792
rect 29052 6752 29736 6780
rect 29052 6740 29058 6752
rect 29730 6740 29736 6752
rect 29788 6740 29794 6792
rect 31128 6766 31156 6820
rect 36541 6817 36553 6820
rect 36587 6817 36599 6851
rect 36541 6811 36599 6817
rect 33042 6740 33048 6792
rect 33100 6780 33106 6792
rect 33413 6783 33471 6789
rect 33413 6780 33425 6783
rect 33100 6752 33425 6780
rect 33100 6740 33106 6752
rect 33413 6749 33425 6752
rect 33459 6749 33471 6783
rect 33413 6743 33471 6749
rect 33502 6740 33508 6792
rect 33560 6780 33566 6792
rect 34054 6780 34060 6792
rect 33560 6752 33605 6780
rect 34015 6752 34060 6780
rect 33560 6740 33566 6752
rect 34054 6740 34060 6752
rect 34112 6740 34118 6792
rect 34149 6783 34207 6789
rect 34149 6749 34161 6783
rect 34195 6780 34207 6783
rect 34882 6780 34888 6792
rect 34195 6752 34888 6780
rect 34195 6749 34207 6752
rect 34149 6743 34207 6749
rect 34882 6740 34888 6752
rect 34940 6740 34946 6792
rect 35526 6740 35532 6792
rect 35584 6780 35590 6792
rect 36633 6783 36691 6789
rect 36633 6780 36645 6783
rect 35584 6752 36645 6780
rect 35584 6740 35590 6752
rect 36633 6749 36645 6752
rect 36679 6780 36691 6783
rect 37274 6780 37280 6792
rect 36679 6752 37280 6780
rect 36679 6749 36691 6752
rect 36633 6743 36691 6749
rect 37274 6740 37280 6752
rect 37332 6780 37338 6792
rect 38197 6783 38255 6789
rect 38197 6780 38209 6783
rect 37332 6752 38209 6780
rect 37332 6740 37338 6752
rect 38197 6749 38209 6752
rect 38243 6749 38255 6783
rect 38197 6743 38255 6749
rect 22097 6715 22155 6721
rect 18892 6684 20852 6712
rect 20714 6644 20720 6656
rect 18340 6616 20720 6644
rect 20714 6604 20720 6616
rect 20772 6604 20778 6656
rect 20824 6644 20852 6684
rect 22097 6681 22109 6715
rect 22143 6681 22155 6715
rect 22097 6675 22155 6681
rect 21910 6644 21916 6656
rect 20824 6616 21916 6644
rect 21910 6604 21916 6616
rect 21968 6604 21974 6656
rect 22112 6644 22140 6675
rect 22186 6672 22192 6724
rect 22244 6712 22250 6724
rect 26234 6712 26240 6724
rect 22244 6684 25070 6712
rect 26195 6684 26240 6712
rect 22244 6672 22250 6684
rect 26234 6672 26240 6684
rect 26292 6672 26298 6724
rect 30282 6712 30288 6724
rect 26344 6684 27554 6712
rect 28920 6684 30288 6712
rect 22370 6644 22376 6656
rect 22112 6616 22376 6644
rect 22370 6604 22376 6616
rect 22428 6604 22434 6656
rect 22738 6604 22744 6656
rect 22796 6644 22802 6656
rect 24029 6647 24087 6653
rect 24029 6644 24041 6647
rect 22796 6616 24041 6644
rect 22796 6604 22802 6616
rect 24029 6613 24041 6616
rect 24075 6644 24087 6647
rect 24302 6644 24308 6656
rect 24075 6616 24308 6644
rect 24075 6613 24087 6616
rect 24029 6607 24087 6613
rect 24302 6604 24308 6616
rect 24360 6604 24366 6656
rect 24854 6604 24860 6656
rect 24912 6644 24918 6656
rect 26344 6644 26372 6684
rect 28920 6656 28948 6684
rect 30282 6672 30288 6684
rect 30340 6672 30346 6724
rect 31662 6672 31668 6724
rect 31720 6712 31726 6724
rect 32585 6715 32643 6721
rect 32585 6712 32597 6715
rect 31720 6684 32597 6712
rect 31720 6672 31726 6684
rect 32585 6681 32597 6684
rect 32631 6681 32643 6715
rect 34900 6712 34928 6740
rect 35342 6712 35348 6724
rect 34900 6684 35348 6712
rect 32585 6675 32643 6681
rect 35342 6672 35348 6684
rect 35400 6712 35406 6724
rect 37645 6715 37703 6721
rect 37645 6712 37657 6715
rect 35400 6684 37657 6712
rect 35400 6672 35406 6684
rect 37645 6681 37657 6684
rect 37691 6681 37703 6715
rect 37645 6675 37703 6681
rect 24912 6616 26372 6644
rect 24912 6604 24918 6616
rect 26418 6604 26424 6656
rect 26476 6644 26482 6656
rect 27982 6644 27988 6656
rect 26476 6616 27988 6644
rect 26476 6604 26482 6616
rect 27982 6604 27988 6616
rect 28040 6644 28046 6656
rect 28810 6644 28816 6656
rect 28040 6616 28816 6644
rect 28040 6604 28046 6616
rect 28810 6604 28816 6616
rect 28868 6604 28874 6656
rect 28902 6604 28908 6656
rect 28960 6604 28966 6656
rect 29546 6604 29552 6656
rect 29604 6644 29610 6656
rect 30926 6644 30932 6656
rect 29604 6616 30932 6644
rect 29604 6604 29610 6616
rect 30926 6604 30932 6616
rect 30984 6604 30990 6656
rect 31018 6604 31024 6656
rect 31076 6644 31082 6656
rect 32033 6647 32091 6653
rect 32033 6644 32045 6647
rect 31076 6616 32045 6644
rect 31076 6604 31082 6616
rect 32033 6613 32045 6616
rect 32079 6613 32091 6647
rect 32033 6607 32091 6613
rect 34514 6604 34520 6656
rect 34572 6644 34578 6656
rect 34885 6647 34943 6653
rect 34885 6644 34897 6647
rect 34572 6616 34897 6644
rect 34572 6604 34578 6616
rect 34885 6613 34897 6616
rect 34931 6644 34943 6647
rect 35437 6647 35495 6653
rect 35437 6644 35449 6647
rect 34931 6616 35449 6644
rect 34931 6613 34943 6616
rect 34885 6607 34943 6613
rect 35437 6613 35449 6616
rect 35483 6613 35495 6647
rect 35437 6607 35495 6613
rect 36630 6604 36636 6656
rect 36688 6644 36694 6656
rect 37093 6647 37151 6653
rect 37093 6644 37105 6647
rect 36688 6616 37105 6644
rect 36688 6604 36694 6616
rect 37093 6613 37105 6616
rect 37139 6644 37151 6647
rect 38010 6644 38016 6656
rect 37139 6616 38016 6644
rect 37139 6613 37151 6616
rect 37093 6607 37151 6613
rect 38010 6604 38016 6616
rect 38068 6604 38074 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 15470 6400 15476 6452
rect 15528 6440 15534 6452
rect 17221 6443 17279 6449
rect 17221 6440 17233 6443
rect 15528 6412 17233 6440
rect 15528 6400 15534 6412
rect 17221 6409 17233 6412
rect 17267 6409 17279 6443
rect 17221 6403 17279 6409
rect 18509 6443 18567 6449
rect 18509 6409 18521 6443
rect 18555 6440 18567 6443
rect 18690 6440 18696 6452
rect 18555 6412 18696 6440
rect 18555 6409 18567 6412
rect 18509 6403 18567 6409
rect 18690 6400 18696 6412
rect 18748 6400 18754 6452
rect 19978 6400 19984 6452
rect 20036 6440 20042 6452
rect 24210 6440 24216 6452
rect 20036 6412 22094 6440
rect 24171 6412 24216 6440
rect 20036 6400 20042 6412
rect 9766 6332 9772 6384
rect 9824 6372 9830 6384
rect 9824 6344 12434 6372
rect 9824 6332 9830 6344
rect 12406 6168 12434 6344
rect 13814 6332 13820 6384
rect 13872 6372 13878 6384
rect 19426 6372 19432 6384
rect 13872 6344 19432 6372
rect 13872 6332 13878 6344
rect 19426 6332 19432 6344
rect 19484 6332 19490 6384
rect 21726 6372 21732 6384
rect 21206 6344 21732 6372
rect 21726 6332 21732 6344
rect 21784 6332 21790 6384
rect 22066 6372 22094 6412
rect 24210 6400 24216 6412
rect 24268 6400 24274 6452
rect 24302 6400 24308 6452
rect 24360 6440 24366 6452
rect 26602 6440 26608 6452
rect 24360 6412 26608 6440
rect 24360 6400 24366 6412
rect 26602 6400 26608 6412
rect 26660 6440 26666 6452
rect 26660 6412 27016 6440
rect 26660 6400 26666 6412
rect 22741 6375 22799 6381
rect 22741 6372 22753 6375
rect 22066 6344 22753 6372
rect 22741 6341 22753 6344
rect 22787 6341 22799 6375
rect 22741 6335 22799 6341
rect 23198 6332 23204 6384
rect 23256 6332 23262 6384
rect 24949 6375 25007 6381
rect 24949 6341 24961 6375
rect 24995 6372 25007 6375
rect 25222 6372 25228 6384
rect 24995 6344 25228 6372
rect 24995 6341 25007 6344
rect 24949 6335 25007 6341
rect 25222 6332 25228 6344
rect 25280 6332 25286 6384
rect 26418 6332 26424 6384
rect 26476 6372 26482 6384
rect 26878 6372 26884 6384
rect 26476 6344 26884 6372
rect 26476 6332 26482 6344
rect 26878 6332 26884 6344
rect 26936 6332 26942 6384
rect 26988 6372 27016 6412
rect 28350 6400 28356 6452
rect 28408 6440 28414 6452
rect 28994 6440 29000 6452
rect 28408 6412 29000 6440
rect 28408 6400 28414 6412
rect 28994 6400 29000 6412
rect 29052 6400 29058 6452
rect 29730 6400 29736 6452
rect 29788 6440 29794 6452
rect 29788 6412 30236 6440
rect 29788 6400 29794 6412
rect 27062 6372 27068 6384
rect 26988 6344 27068 6372
rect 27062 6332 27068 6344
rect 27120 6332 27126 6384
rect 28718 6332 28724 6384
rect 28776 6372 28782 6384
rect 28813 6375 28871 6381
rect 28813 6372 28825 6375
rect 28776 6344 28825 6372
rect 28776 6332 28782 6344
rect 28813 6341 28825 6344
rect 28859 6341 28871 6375
rect 28813 6335 28871 6341
rect 29086 6332 29092 6384
rect 29144 6372 29150 6384
rect 30208 6372 30236 6412
rect 30558 6400 30564 6452
rect 30616 6440 30622 6452
rect 32674 6440 32680 6452
rect 30616 6412 31754 6440
rect 32635 6412 32680 6440
rect 30616 6400 30622 6412
rect 30282 6372 30288 6384
rect 29144 6344 29394 6372
rect 30208 6344 30288 6372
rect 29144 6332 29150 6344
rect 30282 6332 30288 6344
rect 30340 6372 30346 6384
rect 31297 6375 31355 6381
rect 31297 6372 31309 6375
rect 30340 6344 31309 6372
rect 30340 6332 30346 6344
rect 17313 6307 17371 6313
rect 17313 6273 17325 6307
rect 17359 6304 17371 6307
rect 19518 6304 19524 6316
rect 17359 6276 19524 6304
rect 17359 6273 17371 6276
rect 17313 6267 17371 6273
rect 19518 6264 19524 6276
rect 19576 6264 19582 6316
rect 21634 6264 21640 6316
rect 21692 6304 21698 6316
rect 22462 6304 22468 6316
rect 21692 6276 22468 6304
rect 21692 6264 21698 6276
rect 22462 6264 22468 6276
rect 22520 6264 22526 6316
rect 26050 6264 26056 6316
rect 26108 6264 26114 6316
rect 26602 6264 26608 6316
rect 26660 6304 26666 6316
rect 29270 6304 29276 6316
rect 26660 6276 29276 6304
rect 26660 6264 26666 6276
rect 29270 6264 29276 6276
rect 29328 6264 29334 6316
rect 30852 6313 30880 6344
rect 31297 6341 31309 6344
rect 31343 6341 31355 6375
rect 31726 6372 31754 6412
rect 32674 6400 32680 6412
rect 32732 6400 32738 6452
rect 33318 6440 33324 6452
rect 33279 6412 33324 6440
rect 33318 6400 33324 6412
rect 33376 6400 33382 6452
rect 33502 6400 33508 6452
rect 33560 6440 33566 6452
rect 34606 6440 34612 6452
rect 33560 6412 34100 6440
rect 34567 6412 34612 6440
rect 33560 6400 33566 6412
rect 33965 6375 34023 6381
rect 33965 6372 33977 6375
rect 31726 6344 33977 6372
rect 31297 6335 31355 6341
rect 33965 6341 33977 6344
rect 34011 6341 34023 6375
rect 34072 6372 34100 6412
rect 34606 6400 34612 6412
rect 34664 6400 34670 6452
rect 34790 6400 34796 6452
rect 34848 6440 34854 6452
rect 35253 6443 35311 6449
rect 35253 6440 35265 6443
rect 34848 6412 35265 6440
rect 34848 6400 34854 6412
rect 35253 6409 35265 6412
rect 35299 6409 35311 6443
rect 35253 6403 35311 6409
rect 36538 6400 36544 6452
rect 36596 6440 36602 6452
rect 36633 6443 36691 6449
rect 36633 6440 36645 6443
rect 36596 6412 36645 6440
rect 36596 6400 36602 6412
rect 36633 6409 36645 6412
rect 36679 6409 36691 6443
rect 36633 6403 36691 6409
rect 34422 6372 34428 6384
rect 34072 6344 34428 6372
rect 33965 6335 34023 6341
rect 34422 6332 34428 6344
rect 34480 6372 34486 6384
rect 34480 6344 35480 6372
rect 34480 6332 34486 6344
rect 30837 6307 30895 6313
rect 30837 6273 30849 6307
rect 30883 6304 30895 6307
rect 30883 6276 30917 6304
rect 30883 6273 30895 6276
rect 30837 6267 30895 6273
rect 31110 6264 31116 6316
rect 31168 6304 31174 6316
rect 32769 6307 32827 6313
rect 32769 6304 32781 6307
rect 31168 6276 32781 6304
rect 31168 6264 31174 6276
rect 32769 6273 32781 6276
rect 32815 6273 32827 6307
rect 32769 6267 32827 6273
rect 15657 6239 15715 6245
rect 15657 6205 15669 6239
rect 15703 6236 15715 6239
rect 17034 6236 17040 6248
rect 15703 6208 17040 6236
rect 15703 6205 15715 6208
rect 15657 6199 15715 6205
rect 17034 6196 17040 6208
rect 17092 6236 17098 6248
rect 19610 6236 19616 6248
rect 17092 6208 19616 6236
rect 17092 6196 17098 6208
rect 19610 6196 19616 6208
rect 19668 6196 19674 6248
rect 19705 6239 19763 6245
rect 19705 6205 19717 6239
rect 19751 6205 19763 6239
rect 19978 6236 19984 6248
rect 19939 6208 19984 6236
rect 19705 6199 19763 6205
rect 16301 6171 16359 6177
rect 16301 6168 16313 6171
rect 12406 6140 16313 6168
rect 16301 6137 16313 6140
rect 16347 6168 16359 6171
rect 16942 6168 16948 6180
rect 16347 6140 16948 6168
rect 16347 6137 16359 6140
rect 16301 6131 16359 6137
rect 16942 6128 16948 6140
rect 17000 6168 17006 6180
rect 19426 6168 19432 6180
rect 17000 6140 19432 6168
rect 17000 6128 17006 6140
rect 19426 6128 19432 6140
rect 19484 6128 19490 6180
rect 13265 6103 13323 6109
rect 13265 6069 13277 6103
rect 13311 6100 13323 6103
rect 13909 6103 13967 6109
rect 13909 6100 13921 6103
rect 13311 6072 13921 6100
rect 13311 6069 13323 6072
rect 13265 6063 13323 6069
rect 13909 6069 13921 6072
rect 13955 6100 13967 6103
rect 14458 6100 14464 6112
rect 13955 6072 14464 6100
rect 13955 6069 13967 6072
rect 13909 6063 13967 6069
rect 14458 6060 14464 6072
rect 14516 6100 14522 6112
rect 14645 6103 14703 6109
rect 14645 6100 14657 6103
rect 14516 6072 14657 6100
rect 14516 6060 14522 6072
rect 14645 6069 14657 6072
rect 14691 6100 14703 6103
rect 15197 6103 15255 6109
rect 15197 6100 15209 6103
rect 14691 6072 15209 6100
rect 14691 6069 14703 6072
rect 14645 6063 14703 6069
rect 15197 6069 15209 6072
rect 15243 6100 15255 6103
rect 16114 6100 16120 6112
rect 15243 6072 16120 6100
rect 15243 6069 15255 6072
rect 15197 6063 15255 6069
rect 16114 6060 16120 6072
rect 16172 6060 16178 6112
rect 17770 6060 17776 6112
rect 17828 6100 17834 6112
rect 17865 6103 17923 6109
rect 17865 6100 17877 6103
rect 17828 6072 17877 6100
rect 17828 6060 17834 6072
rect 17865 6069 17877 6072
rect 17911 6069 17923 6103
rect 17865 6063 17923 6069
rect 19061 6103 19119 6109
rect 19061 6069 19073 6103
rect 19107 6100 19119 6103
rect 19242 6100 19248 6112
rect 19107 6072 19248 6100
rect 19107 6069 19119 6072
rect 19061 6063 19119 6069
rect 19242 6060 19248 6072
rect 19300 6060 19306 6112
rect 19334 6060 19340 6112
rect 19392 6100 19398 6112
rect 19610 6100 19616 6112
rect 19392 6072 19616 6100
rect 19392 6060 19398 6072
rect 19610 6060 19616 6072
rect 19668 6060 19674 6112
rect 19720 6100 19748 6199
rect 19978 6196 19984 6208
rect 20036 6196 20042 6248
rect 24578 6196 24584 6248
rect 24636 6236 24642 6248
rect 24673 6239 24731 6245
rect 24673 6236 24685 6239
rect 24636 6208 24685 6236
rect 24636 6196 24642 6208
rect 24673 6205 24685 6208
rect 24719 6205 24731 6239
rect 29822 6236 29828 6248
rect 24673 6199 24731 6205
rect 24780 6208 29828 6236
rect 20990 6128 20996 6180
rect 21048 6168 21054 6180
rect 21453 6171 21511 6177
rect 21453 6168 21465 6171
rect 21048 6140 21465 6168
rect 21048 6128 21054 6140
rect 21453 6137 21465 6140
rect 21499 6137 21511 6171
rect 21453 6131 21511 6137
rect 21542 6128 21548 6180
rect 21600 6168 21606 6180
rect 22186 6168 22192 6180
rect 21600 6140 22192 6168
rect 21600 6128 21606 6140
rect 22186 6128 22192 6140
rect 22244 6128 22250 6180
rect 23934 6128 23940 6180
rect 23992 6168 23998 6180
rect 24780 6168 24808 6208
rect 29822 6196 29828 6208
rect 29880 6196 29886 6248
rect 30190 6196 30196 6248
rect 30248 6236 30254 6248
rect 30561 6239 30619 6245
rect 30561 6236 30573 6239
rect 30248 6208 30573 6236
rect 30248 6196 30254 6208
rect 30561 6205 30573 6208
rect 30607 6205 30619 6239
rect 32784 6236 32812 6267
rect 33134 6264 33140 6316
rect 33192 6304 33198 6316
rect 33413 6307 33471 6313
rect 33413 6304 33425 6307
rect 33192 6276 33425 6304
rect 33192 6264 33198 6276
rect 33413 6273 33425 6276
rect 33459 6304 33471 6307
rect 34057 6307 34115 6313
rect 34057 6304 34069 6307
rect 33459 6276 34069 6304
rect 33459 6273 33471 6276
rect 33413 6267 33471 6273
rect 34057 6273 34069 6276
rect 34103 6304 34115 6307
rect 34606 6304 34612 6316
rect 34103 6276 34612 6304
rect 34103 6273 34115 6276
rect 34057 6267 34115 6273
rect 34606 6264 34612 6276
rect 34664 6264 34670 6316
rect 34716 6313 34744 6344
rect 34701 6307 34759 6313
rect 35345 6310 35403 6313
rect 34701 6273 34713 6307
rect 34747 6273 34759 6307
rect 34701 6267 34759 6273
rect 35268 6307 35403 6310
rect 35268 6282 35357 6307
rect 35268 6236 35296 6282
rect 35345 6273 35357 6282
rect 35391 6273 35403 6307
rect 35452 6304 35480 6344
rect 35618 6332 35624 6384
rect 35676 6372 35682 6384
rect 35989 6375 36047 6381
rect 35989 6372 36001 6375
rect 35676 6344 36001 6372
rect 35676 6332 35682 6344
rect 35989 6341 36001 6344
rect 36035 6341 36047 6375
rect 35989 6335 36047 6341
rect 36081 6307 36139 6313
rect 36081 6304 36093 6307
rect 35452 6276 36093 6304
rect 35345 6267 35403 6273
rect 36081 6273 36093 6276
rect 36127 6304 36139 6307
rect 36630 6304 36636 6316
rect 36127 6276 36636 6304
rect 36127 6273 36139 6276
rect 36081 6267 36139 6273
rect 36630 6264 36636 6276
rect 36688 6304 36694 6316
rect 36725 6307 36783 6313
rect 36725 6304 36737 6307
rect 36688 6276 36737 6304
rect 36688 6264 36694 6276
rect 36725 6273 36737 6276
rect 36771 6273 36783 6307
rect 36725 6267 36783 6273
rect 37550 6264 37556 6316
rect 37608 6304 37614 6316
rect 38013 6307 38071 6313
rect 38013 6304 38025 6307
rect 37608 6276 38025 6304
rect 37608 6264 37614 6276
rect 38013 6273 38025 6276
rect 38059 6273 38071 6307
rect 38013 6267 38071 6273
rect 38194 6264 38200 6316
rect 38252 6304 38258 6316
rect 38289 6307 38347 6313
rect 38289 6304 38301 6307
rect 38252 6276 38301 6304
rect 38252 6264 38258 6276
rect 38289 6273 38301 6276
rect 38335 6273 38347 6307
rect 38289 6267 38347 6273
rect 36262 6236 36268 6248
rect 32784 6208 36268 6236
rect 30561 6199 30619 6205
rect 36262 6196 36268 6208
rect 36320 6196 36326 6248
rect 27154 6168 27160 6180
rect 23992 6140 24808 6168
rect 25976 6140 27160 6168
rect 23992 6128 23998 6140
rect 21634 6100 21640 6112
rect 19720 6072 21640 6100
rect 21634 6060 21640 6072
rect 21692 6060 21698 6112
rect 21818 6060 21824 6112
rect 21876 6100 21882 6112
rect 23750 6100 23756 6112
rect 21876 6072 23756 6100
rect 21876 6060 21882 6072
rect 23750 6060 23756 6072
rect 23808 6060 23814 6112
rect 24578 6060 24584 6112
rect 24636 6100 24642 6112
rect 25976 6100 26004 6140
rect 27154 6128 27160 6140
rect 27212 6168 27218 6180
rect 27709 6171 27767 6177
rect 27709 6168 27721 6171
rect 27212 6140 27721 6168
rect 27212 6128 27218 6140
rect 27709 6137 27721 6140
rect 27755 6168 27767 6171
rect 28261 6171 28319 6177
rect 28261 6168 28273 6171
rect 27755 6140 28273 6168
rect 27755 6137 27767 6140
rect 27709 6131 27767 6137
rect 28261 6137 28273 6140
rect 28307 6168 28319 6171
rect 28350 6168 28356 6180
rect 28307 6140 28356 6168
rect 28307 6137 28319 6140
rect 28261 6131 28319 6137
rect 28350 6128 28356 6140
rect 28408 6128 28414 6180
rect 34238 6168 34244 6180
rect 30760 6140 34244 6168
rect 26418 6100 26424 6112
rect 24636 6072 26004 6100
rect 26379 6072 26424 6100
rect 24636 6060 24642 6072
rect 26418 6060 26424 6072
rect 26476 6060 26482 6112
rect 26510 6060 26516 6112
rect 26568 6100 26574 6112
rect 30760 6100 30788 6140
rect 34238 6128 34244 6140
rect 34296 6128 34302 6180
rect 34606 6128 34612 6180
rect 34664 6168 34670 6180
rect 35526 6168 35532 6180
rect 34664 6140 35532 6168
rect 34664 6128 34670 6140
rect 35526 6128 35532 6140
rect 35584 6128 35590 6180
rect 26568 6072 30788 6100
rect 26568 6060 26574 6072
rect 30926 6060 30932 6112
rect 30984 6100 30990 6112
rect 32582 6100 32588 6112
rect 30984 6072 32588 6100
rect 30984 6060 30990 6072
rect 32582 6060 32588 6072
rect 32640 6060 32646 6112
rect 32950 6060 32956 6112
rect 33008 6100 33014 6112
rect 34790 6100 34796 6112
rect 33008 6072 34796 6100
rect 33008 6060 33014 6072
rect 34790 6060 34796 6072
rect 34848 6060 34854 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 14553 5899 14611 5905
rect 14553 5865 14565 5899
rect 14599 5896 14611 5899
rect 14826 5896 14832 5908
rect 14599 5868 14832 5896
rect 14599 5865 14611 5868
rect 14553 5859 14611 5865
rect 14826 5856 14832 5868
rect 14884 5856 14890 5908
rect 16669 5899 16727 5905
rect 16669 5865 16681 5899
rect 16715 5896 16727 5899
rect 17402 5896 17408 5908
rect 16715 5868 17408 5896
rect 16715 5865 16727 5868
rect 16669 5859 16727 5865
rect 17402 5856 17408 5868
rect 17460 5856 17466 5908
rect 18877 5899 18935 5905
rect 18877 5865 18889 5899
rect 18923 5896 18935 5899
rect 19058 5896 19064 5908
rect 18923 5868 19064 5896
rect 18923 5865 18935 5868
rect 18877 5859 18935 5865
rect 19058 5856 19064 5868
rect 19116 5856 19122 5908
rect 19242 5856 19248 5908
rect 19300 5896 19306 5908
rect 20898 5896 20904 5908
rect 19300 5868 20904 5896
rect 19300 5856 19306 5868
rect 20898 5856 20904 5868
rect 20956 5856 20962 5908
rect 20993 5899 21051 5905
rect 20993 5865 21005 5899
rect 21039 5896 21051 5899
rect 21174 5896 21180 5908
rect 21039 5868 21180 5896
rect 21039 5865 21051 5868
rect 20993 5859 21051 5865
rect 21174 5856 21180 5868
rect 21232 5856 21238 5908
rect 21542 5856 21548 5908
rect 21600 5856 21606 5908
rect 22094 5856 22100 5908
rect 22152 5896 22158 5908
rect 23658 5896 23664 5908
rect 22152 5868 23664 5896
rect 22152 5856 22158 5868
rect 23658 5856 23664 5868
rect 23716 5856 23722 5908
rect 23750 5856 23756 5908
rect 23808 5896 23814 5908
rect 25958 5896 25964 5908
rect 23808 5868 25964 5896
rect 23808 5856 23814 5868
rect 25958 5856 25964 5868
rect 26016 5856 26022 5908
rect 26050 5856 26056 5908
rect 26108 5896 26114 5908
rect 26108 5868 31432 5896
rect 26108 5856 26114 5868
rect 17218 5788 17224 5840
rect 17276 5828 17282 5840
rect 17313 5831 17371 5837
rect 17313 5828 17325 5831
rect 17276 5800 17325 5828
rect 17276 5788 17282 5800
rect 17313 5797 17325 5800
rect 17359 5797 17371 5831
rect 21560 5828 21588 5856
rect 17313 5791 17371 5797
rect 17420 5800 21588 5828
rect 23201 5831 23259 5837
rect 14642 5760 14648 5772
rect 6886 5732 14648 5760
rect 2869 5695 2927 5701
rect 2869 5661 2881 5695
rect 2915 5692 2927 5695
rect 6886 5692 6914 5732
rect 14642 5720 14648 5732
rect 14700 5760 14706 5772
rect 15381 5763 15439 5769
rect 15381 5760 15393 5763
rect 14700 5732 15393 5760
rect 14700 5720 14706 5732
rect 15381 5729 15393 5732
rect 15427 5729 15439 5763
rect 16022 5760 16028 5772
rect 15983 5732 16028 5760
rect 15381 5723 15439 5729
rect 16022 5720 16028 5732
rect 16080 5720 16086 5772
rect 16298 5720 16304 5772
rect 16356 5760 16362 5772
rect 17420 5760 17448 5800
rect 23201 5797 23213 5831
rect 23247 5828 23259 5831
rect 23290 5828 23296 5840
rect 23247 5800 23296 5828
rect 23247 5797 23259 5800
rect 23201 5791 23259 5797
rect 23290 5788 23296 5800
rect 23348 5788 23354 5840
rect 24762 5788 24768 5840
rect 24820 5828 24826 5840
rect 24820 5800 25084 5828
rect 24820 5788 24826 5800
rect 16356 5732 17448 5760
rect 16356 5720 16362 5732
rect 19334 5720 19340 5772
rect 19392 5760 19398 5772
rect 25056 5760 25084 5800
rect 26252 5800 27844 5828
rect 26252 5760 26280 5800
rect 19392 5732 24992 5760
rect 25056 5732 26280 5760
rect 19392 5720 19398 5732
rect 2915 5664 6914 5692
rect 13173 5695 13231 5701
rect 2915 5661 2927 5664
rect 2869 5655 2927 5661
rect 13173 5661 13185 5695
rect 13219 5692 13231 5695
rect 13446 5692 13452 5704
rect 13219 5664 13452 5692
rect 13219 5661 13231 5664
rect 13173 5655 13231 5661
rect 13446 5652 13452 5664
rect 13504 5692 13510 5704
rect 13725 5695 13783 5701
rect 13725 5692 13737 5695
rect 13504 5664 13737 5692
rect 13504 5652 13510 5664
rect 13725 5661 13737 5664
rect 13771 5692 13783 5695
rect 14458 5692 14464 5704
rect 13771 5664 14464 5692
rect 13771 5661 13783 5664
rect 13725 5655 13783 5661
rect 14458 5652 14464 5664
rect 14516 5652 14522 5704
rect 16761 5695 16819 5701
rect 16761 5661 16773 5695
rect 16807 5661 16819 5695
rect 16761 5655 16819 5661
rect 17405 5695 17463 5701
rect 17405 5661 17417 5695
rect 17451 5692 17463 5695
rect 20162 5692 20168 5704
rect 17451 5664 20168 5692
rect 17451 5661 17463 5664
rect 17405 5655 17463 5661
rect 15930 5624 15936 5636
rect 15891 5596 15936 5624
rect 15930 5584 15936 5596
rect 15988 5584 15994 5636
rect 16776 5624 16804 5655
rect 20162 5652 20168 5664
rect 20220 5652 20226 5704
rect 20254 5652 20260 5704
rect 20312 5692 20318 5704
rect 20622 5692 20628 5704
rect 20312 5664 20628 5692
rect 20312 5652 20318 5664
rect 20622 5652 20628 5664
rect 20680 5652 20686 5704
rect 21450 5692 21456 5704
rect 21411 5664 21456 5692
rect 21450 5652 21456 5664
rect 21508 5652 21514 5704
rect 22862 5664 23244 5692
rect 24964 5678 24992 5732
rect 26418 5720 26424 5772
rect 26476 5760 26482 5772
rect 26789 5763 26847 5769
rect 26789 5760 26801 5763
rect 26476 5732 26801 5760
rect 26476 5720 26482 5732
rect 26789 5729 26801 5732
rect 26835 5729 26847 5763
rect 26789 5723 26847 5729
rect 27433 5763 27491 5769
rect 27433 5729 27445 5763
rect 27479 5760 27491 5763
rect 27522 5760 27528 5772
rect 27479 5732 27528 5760
rect 27479 5729 27491 5732
rect 27433 5723 27491 5729
rect 27522 5720 27528 5732
rect 27580 5720 27586 5772
rect 19058 5624 19064 5636
rect 16776 5596 19064 5624
rect 19058 5584 19064 5596
rect 19116 5584 19122 5636
rect 20898 5584 20904 5636
rect 20956 5624 20962 5636
rect 21729 5627 21787 5633
rect 20956 5596 21680 5624
rect 20956 5584 20962 5596
rect 2774 5556 2780 5568
rect 2735 5528 2780 5556
rect 2774 5516 2780 5528
rect 2832 5516 2838 5568
rect 13078 5516 13084 5568
rect 13136 5556 13142 5568
rect 16666 5556 16672 5568
rect 13136 5528 16672 5556
rect 13136 5516 13142 5528
rect 16666 5516 16672 5528
rect 16724 5516 16730 5568
rect 18325 5559 18383 5565
rect 18325 5525 18337 5559
rect 18371 5556 18383 5559
rect 18598 5556 18604 5568
rect 18371 5528 18604 5556
rect 18371 5525 18383 5528
rect 18325 5519 18383 5525
rect 18598 5516 18604 5528
rect 18656 5516 18662 5568
rect 19610 5516 19616 5568
rect 19668 5556 19674 5568
rect 19705 5559 19763 5565
rect 19705 5556 19717 5559
rect 19668 5528 19717 5556
rect 19668 5516 19674 5528
rect 19705 5525 19717 5528
rect 19751 5556 19763 5559
rect 19978 5556 19984 5568
rect 19751 5528 19984 5556
rect 19751 5525 19763 5528
rect 19705 5519 19763 5525
rect 19978 5516 19984 5528
rect 20036 5516 20042 5568
rect 21652 5556 21680 5596
rect 21729 5593 21741 5627
rect 21775 5624 21787 5627
rect 23216 5624 23244 5664
rect 26326 5652 26332 5704
rect 26384 5692 26390 5704
rect 27154 5692 27160 5704
rect 26384 5664 27160 5692
rect 26384 5652 26390 5664
rect 27154 5652 27160 5664
rect 27212 5652 27218 5704
rect 27816 5678 27844 5800
rect 29638 5788 29644 5840
rect 29696 5828 29702 5840
rect 29733 5831 29791 5837
rect 29733 5828 29745 5831
rect 29696 5800 29745 5828
rect 29696 5788 29702 5800
rect 29733 5797 29745 5800
rect 29779 5828 29791 5831
rect 30190 5828 30196 5840
rect 29779 5800 30196 5828
rect 29779 5797 29791 5800
rect 29733 5791 29791 5797
rect 30190 5788 30196 5800
rect 30248 5788 30254 5840
rect 31404 5828 31432 5868
rect 31478 5856 31484 5908
rect 31536 5896 31542 5908
rect 32861 5899 32919 5905
rect 32861 5896 32873 5899
rect 31536 5868 32873 5896
rect 31536 5856 31542 5868
rect 32861 5865 32873 5868
rect 32907 5865 32919 5899
rect 32861 5859 32919 5865
rect 33318 5856 33324 5908
rect 33376 5896 33382 5908
rect 36265 5899 36323 5905
rect 36265 5896 36277 5899
rect 33376 5868 36277 5896
rect 33376 5856 33382 5868
rect 36265 5865 36277 5868
rect 36311 5865 36323 5899
rect 36265 5859 36323 5865
rect 34977 5831 35035 5837
rect 34977 5828 34989 5831
rect 31404 5800 34989 5828
rect 34977 5797 34989 5800
rect 35023 5797 35035 5831
rect 34977 5791 35035 5797
rect 28902 5760 28908 5772
rect 28863 5732 28908 5760
rect 28902 5720 28908 5732
rect 28960 5720 28966 5772
rect 30650 5720 30656 5772
rect 30708 5760 30714 5772
rect 31205 5763 31263 5769
rect 31205 5760 31217 5763
rect 30708 5732 31217 5760
rect 30708 5720 30714 5732
rect 31205 5729 31217 5732
rect 31251 5729 31263 5763
rect 31205 5723 31263 5729
rect 31481 5763 31539 5769
rect 31481 5729 31493 5763
rect 31527 5760 31539 5763
rect 31662 5760 31668 5772
rect 31527 5732 31668 5760
rect 31527 5729 31539 5732
rect 31481 5723 31539 5729
rect 31662 5720 31668 5732
rect 31720 5760 31726 5772
rect 31941 5763 31999 5769
rect 31941 5760 31953 5763
rect 31720 5732 31953 5760
rect 31720 5720 31726 5732
rect 31941 5729 31953 5732
rect 31987 5729 31999 5763
rect 31941 5723 31999 5729
rect 32582 5720 32588 5772
rect 32640 5760 32646 5772
rect 37093 5763 37151 5769
rect 37093 5760 37105 5763
rect 32640 5732 37105 5760
rect 32640 5720 32646 5732
rect 37093 5729 37105 5732
rect 37139 5729 37151 5763
rect 37093 5723 37151 5729
rect 29181 5695 29239 5701
rect 29181 5661 29193 5695
rect 29227 5661 29239 5695
rect 32950 5692 32956 5704
rect 32911 5664 32956 5692
rect 29181 5655 29239 5661
rect 26050 5624 26056 5636
rect 21775 5596 22094 5624
rect 23216 5596 24808 5624
rect 26011 5596 26056 5624
rect 21775 5593 21787 5596
rect 21729 5587 21787 5593
rect 21818 5556 21824 5568
rect 21652 5528 21824 5556
rect 21818 5516 21824 5528
rect 21876 5516 21882 5568
rect 22066 5556 22094 5596
rect 23842 5556 23848 5568
rect 22066 5528 23848 5556
rect 23842 5516 23848 5528
rect 23900 5556 23906 5568
rect 24302 5556 24308 5568
rect 23900 5528 24308 5556
rect 23900 5516 23906 5528
rect 24302 5516 24308 5528
rect 24360 5516 24366 5568
rect 24578 5556 24584 5568
rect 24539 5528 24584 5556
rect 24578 5516 24584 5528
rect 24636 5516 24642 5568
rect 24780 5556 24808 5596
rect 26050 5584 26056 5596
rect 26108 5584 26114 5636
rect 28994 5584 29000 5636
rect 29052 5624 29058 5636
rect 29196 5624 29224 5655
rect 32950 5652 32956 5664
rect 33008 5652 33014 5704
rect 33134 5652 33140 5704
rect 33192 5692 33198 5704
rect 33597 5695 33655 5701
rect 33597 5692 33609 5695
rect 33192 5664 33609 5692
rect 33192 5652 33198 5664
rect 33597 5661 33609 5664
rect 33643 5661 33655 5695
rect 34146 5692 34152 5704
rect 34107 5664 34152 5692
rect 33597 5655 33655 5661
rect 34146 5652 34152 5664
rect 34204 5652 34210 5704
rect 34241 5695 34299 5701
rect 34241 5661 34253 5695
rect 34287 5692 34299 5695
rect 35066 5692 35072 5704
rect 34287 5664 35072 5692
rect 34287 5661 34299 5664
rect 34241 5655 34299 5661
rect 35066 5652 35072 5664
rect 35124 5652 35130 5704
rect 35713 5695 35771 5701
rect 35713 5661 35725 5695
rect 35759 5694 35771 5695
rect 35802 5694 35808 5704
rect 35759 5666 35808 5694
rect 35759 5661 35771 5666
rect 35713 5655 35771 5661
rect 35802 5652 35808 5666
rect 35860 5652 35866 5704
rect 36262 5652 36268 5704
rect 36320 5692 36326 5704
rect 36357 5695 36415 5701
rect 36357 5692 36369 5695
rect 36320 5664 36369 5692
rect 36320 5652 36326 5664
rect 36357 5661 36369 5664
rect 36403 5661 36415 5695
rect 36357 5655 36415 5661
rect 37185 5695 37243 5701
rect 37185 5661 37197 5695
rect 37231 5692 37243 5695
rect 37274 5692 37280 5704
rect 37231 5664 37280 5692
rect 37231 5661 37243 5664
rect 37185 5655 37243 5661
rect 37274 5652 37280 5664
rect 37332 5692 37338 5704
rect 37829 5695 37887 5701
rect 37829 5692 37841 5695
rect 37332 5664 37841 5692
rect 37332 5652 37338 5664
rect 37829 5661 37841 5664
rect 37875 5692 37887 5695
rect 38010 5692 38016 5704
rect 37875 5664 38016 5692
rect 37875 5661 37887 5664
rect 37829 5655 37887 5661
rect 38010 5652 38016 5664
rect 38068 5652 38074 5704
rect 29052 5596 29224 5624
rect 29052 5584 29058 5596
rect 29914 5584 29920 5636
rect 29972 5624 29978 5636
rect 33505 5627 33563 5633
rect 33505 5624 33517 5627
rect 29972 5596 30038 5624
rect 31726 5596 33517 5624
rect 29972 5584 29978 5596
rect 31726 5556 31754 5596
rect 33505 5593 33517 5596
rect 33551 5593 33563 5627
rect 33505 5587 33563 5593
rect 35621 5627 35679 5633
rect 35621 5593 35633 5627
rect 35667 5593 35679 5627
rect 35621 5587 35679 5593
rect 24780 5528 31754 5556
rect 32490 5516 32496 5568
rect 32548 5556 32554 5568
rect 35636 5556 35664 5587
rect 32548 5528 35664 5556
rect 32548 5516 32554 5528
rect 37274 5516 37280 5568
rect 37332 5556 37338 5568
rect 37737 5559 37795 5565
rect 37737 5556 37749 5559
rect 37332 5528 37749 5556
rect 37332 5516 37338 5528
rect 37737 5525 37749 5528
rect 37783 5525 37795 5559
rect 37737 5519 37795 5525
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 10505 5355 10563 5361
rect 10505 5321 10517 5355
rect 10551 5352 10563 5355
rect 13538 5352 13544 5364
rect 10551 5324 13544 5352
rect 10551 5321 10563 5324
rect 10505 5315 10563 5321
rect 1854 5216 1860 5228
rect 1815 5188 1860 5216
rect 1854 5176 1860 5188
rect 1912 5216 1918 5228
rect 2317 5219 2375 5225
rect 2317 5216 2329 5219
rect 1912 5188 2329 5216
rect 1912 5176 1918 5188
rect 2317 5185 2329 5188
rect 2363 5185 2375 5219
rect 2317 5179 2375 5185
rect 9953 5219 10011 5225
rect 9953 5185 9965 5219
rect 9999 5216 10011 5219
rect 10520 5216 10548 5315
rect 13538 5312 13544 5324
rect 13596 5312 13602 5364
rect 15010 5352 15016 5364
rect 14971 5324 15016 5352
rect 15010 5312 15016 5324
rect 15068 5312 15074 5364
rect 16574 5352 16580 5364
rect 15856 5324 16580 5352
rect 13078 5284 13084 5296
rect 13039 5256 13084 5284
rect 13078 5244 13084 5256
rect 13136 5244 13142 5296
rect 13725 5287 13783 5293
rect 13725 5253 13737 5287
rect 13771 5284 13783 5287
rect 15856 5284 15884 5324
rect 16574 5312 16580 5324
rect 16632 5312 16638 5364
rect 16758 5312 16764 5364
rect 16816 5352 16822 5364
rect 16816 5324 20852 5352
rect 16816 5312 16822 5324
rect 13771 5256 15884 5284
rect 15948 5256 17172 5284
rect 13771 5253 13783 5256
rect 13725 5247 13783 5253
rect 11882 5216 11888 5228
rect 9999 5188 10548 5216
rect 11843 5188 11888 5216
rect 9999 5185 10011 5188
rect 9953 5179 10011 5185
rect 11882 5176 11888 5188
rect 11940 5216 11946 5228
rect 12345 5219 12403 5225
rect 12345 5216 12357 5219
rect 11940 5188 12357 5216
rect 11940 5176 11946 5188
rect 12345 5185 12357 5188
rect 12391 5185 12403 5219
rect 12345 5179 12403 5185
rect 12989 5219 13047 5225
rect 12989 5185 13001 5219
rect 13035 5216 13047 5219
rect 13446 5216 13452 5228
rect 13035 5188 13452 5216
rect 13035 5185 13047 5188
rect 12989 5179 13047 5185
rect 13446 5176 13452 5188
rect 13504 5176 13510 5228
rect 13817 5219 13875 5225
rect 13817 5185 13829 5219
rect 13863 5216 13875 5219
rect 13906 5216 13912 5228
rect 13863 5188 13912 5216
rect 13863 5185 13875 5188
rect 13817 5179 13875 5185
rect 13906 5176 13912 5188
rect 13964 5176 13970 5228
rect 14277 5219 14335 5225
rect 14277 5185 14289 5219
rect 14323 5216 14335 5219
rect 14458 5216 14464 5228
rect 14323 5188 14464 5216
rect 14323 5185 14335 5188
rect 14277 5179 14335 5185
rect 14458 5176 14464 5188
rect 14516 5176 14522 5228
rect 14918 5216 14924 5228
rect 14879 5188 14924 5216
rect 14918 5176 14924 5188
rect 14976 5176 14982 5228
rect 15838 5216 15844 5228
rect 15799 5188 15844 5216
rect 15838 5176 15844 5188
rect 15896 5176 15902 5228
rect 15948 5225 15976 5256
rect 15933 5219 15991 5225
rect 15933 5185 15945 5219
rect 15979 5185 15991 5219
rect 17034 5216 17040 5228
rect 16995 5188 17040 5216
rect 15933 5179 15991 5185
rect 17034 5176 17040 5188
rect 17092 5176 17098 5228
rect 17144 5216 17172 5256
rect 17402 5244 17408 5296
rect 17460 5284 17466 5296
rect 20824 5284 20852 5324
rect 21450 5312 21456 5364
rect 21508 5352 21514 5364
rect 22097 5355 22155 5361
rect 22097 5352 22109 5355
rect 21508 5324 22109 5352
rect 21508 5312 21514 5324
rect 22097 5321 22109 5324
rect 22143 5352 22155 5355
rect 22462 5352 22468 5364
rect 22143 5324 22468 5352
rect 22143 5321 22155 5324
rect 22097 5315 22155 5321
rect 22462 5312 22468 5324
rect 22520 5312 22526 5364
rect 29638 5352 29644 5364
rect 22664 5324 29644 5352
rect 17460 5256 20010 5284
rect 20824 5256 22094 5284
rect 17460 5244 17466 5256
rect 19886 5216 19892 5228
rect 17144 5188 19892 5216
rect 19886 5176 19892 5188
rect 19944 5176 19950 5228
rect 21450 5176 21456 5228
rect 21508 5216 21514 5228
rect 22066 5216 22094 5256
rect 22186 5244 22192 5296
rect 22244 5284 22250 5296
rect 22664 5284 22692 5324
rect 29638 5312 29644 5324
rect 29696 5312 29702 5364
rect 29914 5352 29920 5364
rect 29840 5324 29920 5352
rect 23106 5284 23112 5296
rect 22244 5256 22692 5284
rect 23067 5256 23112 5284
rect 22244 5244 22250 5256
rect 23106 5244 23112 5256
rect 23164 5244 23170 5296
rect 24026 5244 24032 5296
rect 24084 5284 24090 5296
rect 24394 5284 24400 5296
rect 24084 5256 24400 5284
rect 24084 5244 24090 5256
rect 24394 5244 24400 5256
rect 24452 5244 24458 5296
rect 25774 5244 25780 5296
rect 25832 5284 25838 5296
rect 26145 5287 26203 5293
rect 26145 5284 26157 5287
rect 25832 5256 26157 5284
rect 25832 5244 25838 5256
rect 26145 5253 26157 5256
rect 26191 5253 26203 5287
rect 26145 5247 26203 5253
rect 26510 5244 26516 5296
rect 26568 5284 26574 5296
rect 29840 5293 29868 5324
rect 29914 5312 29920 5324
rect 29972 5312 29978 5364
rect 30282 5312 30288 5364
rect 30340 5352 30346 5364
rect 30561 5355 30619 5361
rect 30561 5352 30573 5355
rect 30340 5324 30573 5352
rect 30340 5312 30346 5324
rect 30561 5321 30573 5324
rect 30607 5321 30619 5355
rect 30561 5315 30619 5321
rect 29825 5287 29883 5293
rect 26568 5256 28658 5284
rect 26568 5244 26574 5256
rect 29825 5253 29837 5287
rect 29871 5253 29883 5287
rect 29825 5247 29883 5253
rect 32030 5244 32036 5296
rect 32088 5284 32094 5296
rect 33778 5284 33784 5296
rect 32088 5256 32614 5284
rect 33739 5256 33784 5284
rect 32088 5244 32094 5256
rect 33778 5244 33784 5256
rect 33836 5244 33842 5296
rect 37918 5244 37924 5296
rect 37976 5284 37982 5296
rect 38013 5287 38071 5293
rect 38013 5284 38025 5287
rect 37976 5256 38025 5284
rect 37976 5244 37982 5256
rect 38013 5253 38025 5256
rect 38059 5253 38071 5287
rect 38013 5247 38071 5253
rect 38102 5244 38108 5296
rect 38160 5284 38166 5296
rect 38197 5287 38255 5293
rect 38197 5284 38209 5287
rect 38160 5256 38209 5284
rect 38160 5244 38166 5256
rect 38197 5253 38209 5256
rect 38243 5253 38255 5287
rect 38197 5247 38255 5253
rect 23198 5216 23204 5228
rect 21508 5188 21553 5216
rect 22066 5188 23204 5216
rect 21508 5176 21514 5188
rect 23198 5176 23204 5188
rect 23256 5176 23262 5228
rect 24118 5216 24124 5228
rect 24079 5188 24124 5216
rect 24118 5176 24124 5188
rect 24176 5176 24182 5228
rect 16758 5148 16764 5160
rect 14292 5120 16764 5148
rect 12434 5040 12440 5092
rect 12492 5080 12498 5092
rect 12492 5052 12537 5080
rect 12492 5040 12498 5052
rect 1670 5012 1676 5024
rect 1631 4984 1676 5012
rect 1670 4972 1676 4984
rect 1728 4972 1734 5024
rect 9766 5012 9772 5024
rect 9727 4984 9772 5012
rect 9766 4972 9772 4984
rect 9824 4972 9830 5024
rect 11793 5015 11851 5021
rect 11793 4981 11805 5015
rect 11839 5012 11851 5015
rect 14292 5012 14320 5120
rect 16758 5108 16764 5120
rect 16816 5108 16822 5160
rect 18322 5108 18328 5160
rect 18380 5148 18386 5160
rect 18693 5151 18751 5157
rect 18693 5148 18705 5151
rect 18380 5120 18705 5148
rect 18380 5108 18386 5120
rect 18693 5117 18705 5120
rect 18739 5148 18751 5151
rect 19242 5148 19248 5160
rect 18739 5120 19248 5148
rect 18739 5117 18751 5120
rect 18693 5111 18751 5117
rect 19242 5108 19248 5120
rect 19300 5108 19306 5160
rect 20806 5108 20812 5160
rect 20864 5148 20870 5160
rect 21177 5151 21235 5157
rect 21177 5148 21189 5151
rect 20864 5120 21189 5148
rect 20864 5108 20870 5120
rect 21177 5117 21189 5120
rect 21223 5117 21235 5151
rect 21177 5111 21235 5117
rect 21634 5108 21640 5160
rect 21692 5148 21698 5160
rect 22186 5148 22192 5160
rect 21692 5120 22192 5148
rect 21692 5108 21698 5120
rect 22186 5108 22192 5120
rect 22244 5108 22250 5160
rect 24946 5148 24952 5160
rect 22296 5120 24952 5148
rect 14642 5040 14648 5092
rect 14700 5080 14706 5092
rect 14700 5052 19840 5080
rect 14700 5040 14706 5052
rect 11839 4984 14320 5012
rect 11839 4981 11851 4984
rect 11793 4975 11851 4981
rect 14366 4972 14372 5024
rect 14424 5012 14430 5024
rect 16850 5012 16856 5024
rect 14424 4984 14469 5012
rect 16811 4984 16856 5012
rect 14424 4972 14430 4984
rect 16850 4972 16856 4984
rect 16908 4972 16914 5024
rect 17589 5015 17647 5021
rect 17589 4981 17601 5015
rect 17635 5012 17647 5015
rect 17770 5012 17776 5024
rect 17635 4984 17776 5012
rect 17635 4981 17647 4984
rect 17589 4975 17647 4981
rect 17770 4972 17776 4984
rect 17828 4972 17834 5024
rect 18138 5012 18144 5024
rect 18099 4984 18144 5012
rect 18138 4972 18144 4984
rect 18196 4972 18202 5024
rect 19242 5012 19248 5024
rect 19203 4984 19248 5012
rect 19242 4972 19248 4984
rect 19300 4972 19306 5024
rect 19702 5012 19708 5024
rect 19663 4984 19708 5012
rect 19702 4972 19708 4984
rect 19760 4972 19766 5024
rect 19812 5012 19840 5052
rect 19886 5040 19892 5092
rect 19944 5080 19950 5092
rect 20070 5080 20076 5092
rect 19944 5052 20076 5080
rect 19944 5040 19950 5052
rect 20070 5040 20076 5052
rect 20128 5040 20134 5092
rect 22296 5080 22324 5120
rect 24946 5108 24952 5120
rect 25004 5108 25010 5160
rect 25130 5108 25136 5160
rect 25188 5148 25194 5160
rect 25188 5120 25452 5148
rect 25188 5108 25194 5120
rect 22554 5080 22560 5092
rect 21376 5052 22324 5080
rect 22388 5052 22560 5080
rect 21376 5012 21404 5052
rect 19812 4984 21404 5012
rect 22186 4972 22192 5024
rect 22244 5012 22250 5024
rect 22388 5012 22416 5052
rect 22554 5040 22560 5052
rect 22612 5080 22618 5092
rect 24026 5080 24032 5092
rect 22612 5052 24032 5080
rect 22612 5040 22618 5052
rect 24026 5040 24032 5052
rect 24084 5040 24090 5092
rect 22244 4984 22416 5012
rect 22244 4972 22250 4984
rect 22462 4972 22468 5024
rect 22520 5012 22526 5024
rect 22649 5015 22707 5021
rect 22649 5012 22661 5015
rect 22520 4984 22661 5012
rect 22520 4972 22526 4984
rect 22649 4981 22661 4984
rect 22695 5012 22707 5015
rect 23014 5012 23020 5024
rect 22695 4984 23020 5012
rect 22695 4981 22707 4984
rect 22649 4975 22707 4981
rect 23014 4972 23020 4984
rect 23072 4972 23078 5024
rect 25424 5012 25452 5120
rect 25516 5080 25544 5202
rect 26878 5176 26884 5228
rect 26936 5216 26942 5228
rect 30101 5219 30159 5225
rect 26936 5188 28672 5216
rect 26936 5176 26942 5188
rect 27982 5108 27988 5160
rect 28040 5148 28046 5160
rect 28077 5151 28135 5157
rect 28077 5148 28089 5151
rect 28040 5120 28089 5148
rect 28040 5108 28046 5120
rect 28077 5117 28089 5120
rect 28123 5117 28135 5151
rect 28644 5148 28672 5188
rect 30101 5185 30113 5219
rect 30147 5216 30159 5219
rect 30282 5216 30288 5228
rect 30147 5188 30288 5216
rect 30147 5185 30159 5188
rect 30101 5179 30159 5185
rect 30282 5176 30288 5188
rect 30340 5176 30346 5228
rect 31294 5176 31300 5228
rect 31352 5216 31358 5228
rect 31573 5219 31631 5225
rect 31573 5216 31585 5219
rect 31352 5188 31585 5216
rect 31352 5176 31358 5188
rect 31573 5185 31585 5188
rect 31619 5185 31631 5219
rect 31573 5179 31631 5185
rect 34146 5176 34152 5228
rect 34204 5216 34210 5228
rect 34330 5216 34336 5228
rect 34204 5188 34336 5216
rect 34204 5176 34210 5188
rect 34330 5176 34336 5188
rect 34388 5176 34394 5228
rect 34514 5176 34520 5228
rect 34572 5216 34578 5228
rect 34609 5219 34667 5225
rect 34609 5216 34621 5219
rect 34572 5188 34621 5216
rect 34572 5176 34578 5188
rect 34609 5185 34621 5188
rect 34655 5185 34667 5219
rect 34609 5179 34667 5185
rect 34701 5219 34759 5225
rect 34701 5185 34713 5219
rect 34747 5216 34759 5219
rect 34790 5216 34796 5228
rect 34747 5188 34796 5216
rect 34747 5185 34759 5188
rect 34701 5179 34759 5185
rect 34790 5176 34796 5188
rect 34848 5176 34854 5228
rect 35066 5176 35072 5228
rect 35124 5216 35130 5228
rect 35345 5219 35403 5225
rect 35345 5216 35357 5219
rect 35124 5188 35357 5216
rect 35124 5176 35130 5188
rect 35345 5185 35357 5188
rect 35391 5216 35403 5219
rect 35989 5219 36047 5225
rect 35989 5216 36001 5219
rect 35391 5188 36001 5216
rect 35391 5185 35403 5188
rect 35345 5179 35403 5185
rect 35989 5185 36001 5188
rect 36035 5216 36047 5219
rect 36262 5216 36268 5228
rect 36035 5188 36268 5216
rect 36035 5185 36047 5188
rect 35989 5179 36047 5185
rect 36262 5176 36268 5188
rect 36320 5216 36326 5228
rect 36633 5219 36691 5225
rect 36633 5216 36645 5219
rect 36320 5188 36645 5216
rect 36320 5176 36326 5188
rect 36633 5185 36645 5188
rect 36679 5185 36691 5219
rect 36633 5179 36691 5185
rect 29454 5148 29460 5160
rect 28644 5120 29460 5148
rect 28077 5111 28135 5117
rect 29454 5108 29460 5120
rect 29512 5108 29518 5160
rect 31665 5151 31723 5157
rect 31665 5117 31677 5151
rect 31711 5148 31723 5151
rect 33686 5148 33692 5160
rect 31711 5120 33692 5148
rect 31711 5117 31723 5120
rect 31665 5111 31723 5117
rect 33686 5108 33692 5120
rect 33744 5108 33750 5160
rect 34054 5148 34060 5160
rect 34015 5120 34060 5148
rect 34054 5108 34060 5120
rect 34112 5148 34118 5160
rect 34422 5148 34428 5160
rect 34112 5120 34428 5148
rect 34112 5108 34118 5120
rect 34422 5108 34428 5120
rect 34480 5108 34486 5160
rect 25516 5052 28856 5080
rect 27157 5015 27215 5021
rect 27157 5012 27169 5015
rect 25424 4984 27169 5012
rect 27157 4981 27169 4984
rect 27203 4981 27215 5015
rect 28828 5012 28856 5052
rect 34330 5040 34336 5092
rect 34388 5080 34394 5092
rect 35253 5083 35311 5089
rect 35253 5080 35265 5083
rect 34388 5052 35265 5080
rect 34388 5040 34394 5052
rect 35253 5049 35265 5052
rect 35299 5049 35311 5083
rect 35253 5043 35311 5049
rect 31570 5012 31576 5024
rect 28828 4984 31576 5012
rect 27157 4975 27215 4981
rect 31570 4972 31576 4984
rect 31628 4972 31634 5024
rect 32306 5012 32312 5024
rect 32267 4984 32312 5012
rect 32306 4972 32312 4984
rect 32364 4972 32370 5024
rect 35894 5012 35900 5024
rect 35855 4984 35900 5012
rect 35894 4972 35900 4984
rect 35952 4972 35958 5024
rect 36538 5012 36544 5024
rect 36499 4984 36544 5012
rect 36538 4972 36544 4984
rect 36596 4972 36602 5024
rect 37550 5012 37556 5024
rect 37511 4984 37556 5012
rect 37550 4972 37556 4984
rect 37608 4972 37614 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 12342 4808 12348 4820
rect 12303 4780 12348 4808
rect 12342 4768 12348 4780
rect 12400 4768 12406 4820
rect 13633 4811 13691 4817
rect 13633 4777 13645 4811
rect 13679 4808 13691 4811
rect 13814 4808 13820 4820
rect 13679 4780 13820 4808
rect 13679 4777 13691 4780
rect 13633 4771 13691 4777
rect 13814 4768 13820 4780
rect 13872 4768 13878 4820
rect 14642 4808 14648 4820
rect 14603 4780 14648 4808
rect 14642 4768 14648 4780
rect 14700 4768 14706 4820
rect 15289 4811 15347 4817
rect 15289 4777 15301 4811
rect 15335 4808 15347 4811
rect 15930 4808 15936 4820
rect 15335 4780 15936 4808
rect 15335 4777 15347 4780
rect 15289 4771 15347 4777
rect 15930 4768 15936 4780
rect 15988 4768 15994 4820
rect 16022 4768 16028 4820
rect 16080 4808 16086 4820
rect 22830 4808 22836 4820
rect 16080 4780 22836 4808
rect 16080 4768 16086 4780
rect 22830 4768 22836 4780
rect 22888 4768 22894 4820
rect 22925 4811 22983 4817
rect 22925 4777 22937 4811
rect 22971 4808 22983 4811
rect 23014 4808 23020 4820
rect 22971 4780 23020 4808
rect 22971 4777 22983 4780
rect 22925 4771 22983 4777
rect 23014 4768 23020 4780
rect 23072 4808 23078 4820
rect 24118 4808 24124 4820
rect 23072 4780 24124 4808
rect 23072 4768 23078 4780
rect 24118 4768 24124 4780
rect 24176 4768 24182 4820
rect 24210 4768 24216 4820
rect 24268 4808 24274 4820
rect 24268 4780 24808 4808
rect 24268 4768 24274 4780
rect 12989 4743 13047 4749
rect 12989 4709 13001 4743
rect 13035 4740 13047 4743
rect 19334 4740 19340 4752
rect 13035 4712 19340 4740
rect 13035 4709 13047 4712
rect 12989 4703 13047 4709
rect 19334 4700 19340 4712
rect 19392 4700 19398 4752
rect 19702 4700 19708 4752
rect 19760 4740 19766 4752
rect 20346 4740 20352 4752
rect 19760 4712 20352 4740
rect 19760 4700 19766 4712
rect 20346 4700 20352 4712
rect 20404 4700 20410 4752
rect 22370 4740 22376 4752
rect 22331 4712 22376 4740
rect 22370 4700 22376 4712
rect 22428 4700 22434 4752
rect 23937 4743 23995 4749
rect 23937 4709 23949 4743
rect 23983 4740 23995 4743
rect 24670 4740 24676 4752
rect 23983 4712 24676 4740
rect 23983 4709 23995 4712
rect 23937 4703 23995 4709
rect 24670 4700 24676 4712
rect 24728 4700 24734 4752
rect 24780 4740 24808 4780
rect 24854 4768 24860 4820
rect 24912 4808 24918 4820
rect 26418 4808 26424 4820
rect 24912 4780 26424 4808
rect 24912 4768 24918 4780
rect 26418 4768 26424 4780
rect 26476 4768 26482 4820
rect 26694 4768 26700 4820
rect 26752 4808 26758 4820
rect 26789 4811 26847 4817
rect 26789 4808 26801 4811
rect 26752 4780 26801 4808
rect 26752 4768 26758 4780
rect 26789 4777 26801 4780
rect 26835 4808 26847 4811
rect 31294 4808 31300 4820
rect 26835 4780 31300 4808
rect 26835 4777 26847 4780
rect 26789 4771 26847 4777
rect 31294 4768 31300 4780
rect 31352 4768 31358 4820
rect 31386 4768 31392 4820
rect 31444 4808 31450 4820
rect 32214 4817 32220 4820
rect 31481 4811 31539 4817
rect 31481 4808 31493 4811
rect 31444 4780 31493 4808
rect 31444 4768 31450 4780
rect 31481 4777 31493 4780
rect 31527 4777 31539 4811
rect 31481 4771 31539 4777
rect 32204 4811 32220 4817
rect 32204 4777 32216 4811
rect 32204 4771 32220 4777
rect 32214 4768 32220 4771
rect 32272 4768 32278 4820
rect 33244 4780 37596 4808
rect 24780 4712 24992 4740
rect 20254 4672 20260 4684
rect 15672 4644 20260 4672
rect 11790 4604 11796 4616
rect 11751 4576 11796 4604
rect 11790 4564 11796 4576
rect 11848 4604 11854 4616
rect 12253 4607 12311 4613
rect 12253 4604 12265 4607
rect 11848 4576 12265 4604
rect 11848 4564 11854 4576
rect 12253 4573 12265 4576
rect 12299 4573 12311 4607
rect 12253 4567 12311 4573
rect 12897 4607 12955 4613
rect 12897 4573 12909 4607
rect 12943 4604 12955 4607
rect 13446 4604 13452 4616
rect 12943 4576 13452 4604
rect 12943 4573 12955 4576
rect 12897 4567 12955 4573
rect 13446 4564 13452 4576
rect 13504 4604 13510 4616
rect 13541 4607 13599 4613
rect 13541 4604 13553 4607
rect 13504 4576 13553 4604
rect 13504 4564 13510 4576
rect 13541 4573 13553 4576
rect 13587 4573 13599 4607
rect 13541 4567 13599 4573
rect 13906 4564 13912 4616
rect 13964 4604 13970 4616
rect 14553 4607 14611 4613
rect 14553 4604 14565 4607
rect 13964 4576 14565 4604
rect 13964 4564 13970 4576
rect 14553 4573 14565 4576
rect 14599 4604 14611 4607
rect 14918 4604 14924 4616
rect 14599 4576 14924 4604
rect 14599 4573 14611 4576
rect 14553 4567 14611 4573
rect 14918 4564 14924 4576
rect 14976 4604 14982 4616
rect 15286 4604 15292 4616
rect 14976 4576 15292 4604
rect 14976 4564 14982 4576
rect 15286 4564 15292 4576
rect 15344 4564 15350 4616
rect 15381 4607 15439 4613
rect 15381 4573 15393 4607
rect 15427 4604 15439 4607
rect 15672 4604 15700 4644
rect 20254 4632 20260 4644
rect 20312 4632 20318 4684
rect 20625 4675 20683 4681
rect 20625 4641 20637 4675
rect 20671 4672 20683 4675
rect 21450 4672 21456 4684
rect 20671 4644 21456 4672
rect 20671 4641 20683 4644
rect 20625 4635 20683 4641
rect 15838 4604 15844 4616
rect 15427 4576 15700 4604
rect 15799 4576 15844 4604
rect 15427 4573 15439 4576
rect 15381 4567 15439 4573
rect 15838 4564 15844 4576
rect 15896 4564 15902 4616
rect 16477 4601 16535 4607
rect 16477 4598 16489 4601
rect 16408 4570 16489 4598
rect 11701 4539 11759 4545
rect 11701 4505 11713 4539
rect 11747 4536 11759 4539
rect 16022 4536 16028 4548
rect 11747 4508 16028 4536
rect 11747 4505 11759 4508
rect 11701 4499 11759 4505
rect 16022 4496 16028 4508
rect 16080 4496 16086 4548
rect 15930 4468 15936 4480
rect 15891 4440 15936 4468
rect 15930 4428 15936 4440
rect 15988 4428 15994 4480
rect 16114 4428 16120 4480
rect 16172 4468 16178 4480
rect 16408 4468 16436 4570
rect 16477 4567 16489 4570
rect 16523 4567 16535 4601
rect 16477 4561 16535 4567
rect 16666 4564 16672 4616
rect 16724 4604 16730 4616
rect 17129 4607 17187 4613
rect 17129 4604 17141 4607
rect 16724 4576 17141 4604
rect 16724 4564 16730 4576
rect 17129 4573 17141 4576
rect 17175 4604 17187 4607
rect 17586 4604 17592 4616
rect 17175 4576 17592 4604
rect 17175 4573 17187 4576
rect 17129 4567 17187 4573
rect 17586 4564 17592 4576
rect 17644 4564 17650 4616
rect 19426 4604 19432 4616
rect 19306 4576 19432 4604
rect 17218 4536 17224 4548
rect 17179 4508 17224 4536
rect 17218 4496 17224 4508
rect 17276 4496 17282 4548
rect 19306 4536 19334 4576
rect 19426 4564 19432 4576
rect 19484 4564 19490 4616
rect 19613 4607 19671 4613
rect 19613 4573 19625 4607
rect 19659 4604 19671 4607
rect 20165 4607 20223 4613
rect 20165 4604 20177 4607
rect 19659 4576 20177 4604
rect 19659 4573 19671 4576
rect 19613 4567 19671 4573
rect 20165 4573 20177 4576
rect 20211 4604 20223 4607
rect 20456 4604 20576 4606
rect 20640 4604 20668 4635
rect 21450 4632 21456 4644
rect 21508 4632 21514 4684
rect 23750 4632 23756 4684
rect 23808 4672 23814 4684
rect 24486 4672 24492 4684
rect 23808 4644 24492 4672
rect 23808 4632 23814 4644
rect 24486 4632 24492 4644
rect 24544 4672 24550 4684
rect 24581 4675 24639 4681
rect 24581 4672 24593 4675
rect 24544 4644 24593 4672
rect 24544 4632 24550 4644
rect 24581 4641 24593 4644
rect 24627 4641 24639 4675
rect 24581 4635 24639 4641
rect 24854 4632 24860 4684
rect 24912 4632 24918 4684
rect 24964 4672 24992 4712
rect 26053 4675 26111 4681
rect 26053 4672 26065 4675
rect 24964 4644 26065 4672
rect 26053 4641 26065 4644
rect 26099 4641 26111 4675
rect 28258 4672 28264 4684
rect 28219 4644 28264 4672
rect 26053 4635 26111 4641
rect 28258 4632 28264 4644
rect 28316 4632 28322 4684
rect 28537 4675 28595 4681
rect 28537 4641 28549 4675
rect 28583 4672 28595 4675
rect 28994 4672 29000 4684
rect 28583 4644 29000 4672
rect 28583 4641 28595 4644
rect 28537 4635 28595 4641
rect 28994 4632 29000 4644
rect 29052 4672 29058 4684
rect 29733 4675 29791 4681
rect 29733 4672 29745 4675
rect 29052 4644 29745 4672
rect 29052 4632 29058 4644
rect 29733 4641 29745 4644
rect 29779 4641 29791 4675
rect 29733 4635 29791 4641
rect 31294 4632 31300 4684
rect 31352 4672 31358 4684
rect 33244 4672 33272 4780
rect 33502 4700 33508 4752
rect 33560 4740 33566 4752
rect 37568 4749 37596 4780
rect 33689 4743 33747 4749
rect 33689 4740 33701 4743
rect 33560 4712 33701 4740
rect 33560 4700 33566 4712
rect 33689 4709 33701 4712
rect 33735 4709 33747 4743
rect 33689 4703 33747 4709
rect 37553 4743 37611 4749
rect 37553 4709 37565 4743
rect 37599 4709 37611 4743
rect 37553 4703 37611 4709
rect 35894 4672 35900 4684
rect 31352 4644 33272 4672
rect 34072 4644 35900 4672
rect 31352 4632 31358 4644
rect 20211 4578 20668 4604
rect 20211 4576 20484 4578
rect 20548 4576 20668 4578
rect 20211 4573 20223 4576
rect 20165 4567 20223 4573
rect 18248 4508 19334 4536
rect 16172 4440 16436 4468
rect 16577 4471 16635 4477
rect 16172 4428 16178 4440
rect 16577 4437 16589 4471
rect 16623 4468 16635 4471
rect 18248 4468 18276 4508
rect 16623 4440 18276 4468
rect 18325 4471 18383 4477
rect 16623 4437 16635 4440
rect 16577 4431 16635 4437
rect 18325 4437 18337 4471
rect 18371 4468 18383 4471
rect 18598 4468 18604 4480
rect 18371 4440 18604 4468
rect 18371 4437 18383 4440
rect 18325 4431 18383 4437
rect 18598 4428 18604 4440
rect 18656 4468 18662 4480
rect 18785 4471 18843 4477
rect 18785 4468 18797 4471
rect 18656 4440 18797 4468
rect 18656 4428 18662 4440
rect 18785 4437 18797 4440
rect 18831 4468 18843 4471
rect 19242 4468 19248 4480
rect 18831 4440 19248 4468
rect 18831 4437 18843 4440
rect 18785 4431 18843 4437
rect 19242 4428 19248 4440
rect 19300 4468 19306 4480
rect 19628 4468 19656 4567
rect 23014 4564 23020 4616
rect 23072 4604 23078 4616
rect 23845 4607 23903 4613
rect 23845 4604 23857 4607
rect 23072 4576 23857 4604
rect 23072 4564 23078 4576
rect 23845 4573 23857 4576
rect 23891 4604 23903 4607
rect 24872 4604 24900 4632
rect 23891 4576 24900 4604
rect 23891 4573 23903 4576
rect 23845 4567 23903 4573
rect 26326 4564 26332 4616
rect 26384 4604 26390 4616
rect 26384 4576 26429 4604
rect 31142 4576 31432 4604
rect 26384 4564 26390 4576
rect 20254 4496 20260 4548
rect 20312 4536 20318 4548
rect 20898 4536 20904 4548
rect 20312 4508 20904 4536
rect 20312 4496 20318 4508
rect 20898 4496 20904 4508
rect 20956 4496 20962 4548
rect 21634 4496 21640 4548
rect 21692 4496 21698 4548
rect 22296 4508 22784 4536
rect 19300 4440 19656 4468
rect 19300 4428 19306 4440
rect 20162 4428 20168 4480
rect 20220 4468 20226 4480
rect 22296 4468 22324 4508
rect 20220 4440 22324 4468
rect 22756 4468 22784 4508
rect 22830 4496 22836 4548
rect 22888 4536 22894 4548
rect 22888 4508 24886 4536
rect 26160 4508 27094 4536
rect 22888 4496 22894 4508
rect 23750 4468 23756 4480
rect 22756 4440 23756 4468
rect 20220 4428 20226 4440
rect 23750 4428 23756 4440
rect 23808 4428 23814 4480
rect 24670 4428 24676 4480
rect 24728 4468 24734 4480
rect 26160 4468 26188 4508
rect 28902 4496 28908 4548
rect 28960 4536 28966 4548
rect 28960 4508 29132 4536
rect 28960 4496 28966 4508
rect 28994 4468 29000 4480
rect 24728 4440 26188 4468
rect 28955 4440 29000 4468
rect 24728 4428 24734 4440
rect 28994 4428 29000 4440
rect 29052 4428 29058 4480
rect 29104 4468 29132 4508
rect 29178 4496 29184 4548
rect 29236 4536 29242 4548
rect 30009 4539 30067 4545
rect 30009 4536 30021 4539
rect 29236 4508 30021 4536
rect 29236 4496 29242 4508
rect 30009 4505 30021 4508
rect 30055 4505 30067 4539
rect 31404 4536 31432 4576
rect 31662 4564 31668 4616
rect 31720 4604 31726 4616
rect 31941 4607 31999 4613
rect 31941 4604 31953 4607
rect 31720 4576 31953 4604
rect 31720 4564 31726 4576
rect 31941 4573 31953 4576
rect 31987 4573 31999 4607
rect 33428 4604 33640 4606
rect 34072 4604 34100 4644
rect 35894 4632 35900 4644
rect 35952 4632 35958 4684
rect 36280 4644 37044 4672
rect 33350 4578 34100 4604
rect 33350 4576 33456 4578
rect 33612 4576 34100 4578
rect 31941 4567 31999 4573
rect 34146 4564 34152 4616
rect 34204 4604 34210 4616
rect 34333 4607 34391 4613
rect 34333 4604 34345 4607
rect 34204 4576 34345 4604
rect 34204 4564 34210 4576
rect 34333 4573 34345 4576
rect 34379 4573 34391 4607
rect 34333 4567 34391 4573
rect 34606 4564 34612 4616
rect 34664 4604 34670 4616
rect 35069 4607 35127 4613
rect 35069 4604 35081 4607
rect 34664 4576 35081 4604
rect 34664 4564 34670 4576
rect 35069 4573 35081 4576
rect 35115 4604 35127 4607
rect 35713 4607 35771 4613
rect 35713 4604 35725 4607
rect 35115 4576 35725 4604
rect 35115 4573 35127 4576
rect 35069 4567 35127 4573
rect 35713 4573 35725 4576
rect 35759 4573 35771 4607
rect 35713 4567 35771 4573
rect 35802 4564 35808 4616
rect 35860 4604 35866 4616
rect 36280 4604 36308 4644
rect 35860 4576 36308 4604
rect 35860 4564 35866 4576
rect 36354 4564 36360 4616
rect 36412 4604 36418 4616
rect 37016 4613 37044 4644
rect 37001 4607 37059 4613
rect 36412 4576 36457 4604
rect 36412 4564 36418 4576
rect 37001 4573 37013 4607
rect 37047 4573 37059 4607
rect 37642 4604 37648 4616
rect 37603 4576 37648 4604
rect 37001 4567 37059 4573
rect 37642 4564 37648 4576
rect 37700 4564 37706 4616
rect 38010 4564 38016 4616
rect 38068 4604 38074 4616
rect 38105 4607 38163 4613
rect 38105 4604 38117 4607
rect 38068 4576 38117 4604
rect 38068 4564 38074 4576
rect 38105 4573 38117 4576
rect 38151 4573 38163 4607
rect 38105 4567 38163 4573
rect 32490 4536 32496 4548
rect 31404 4508 32496 4536
rect 30009 4499 30067 4505
rect 32490 4496 32496 4508
rect 32548 4496 32554 4548
rect 36909 4539 36967 4545
rect 36909 4536 36921 4539
rect 33612 4508 36921 4536
rect 33612 4468 33640 4508
rect 36909 4505 36921 4508
rect 36955 4505 36967 4539
rect 38197 4539 38255 4545
rect 38197 4536 38209 4539
rect 36909 4499 36967 4505
rect 37016 4508 38209 4536
rect 37016 4480 37044 4508
rect 38197 4505 38209 4508
rect 38243 4505 38255 4539
rect 38197 4499 38255 4505
rect 29104 4440 33640 4468
rect 33778 4428 33784 4480
rect 33836 4468 33842 4480
rect 34149 4471 34207 4477
rect 34149 4468 34161 4471
rect 33836 4440 34161 4468
rect 33836 4428 33842 4440
rect 34149 4437 34161 4440
rect 34195 4437 34207 4471
rect 34974 4468 34980 4480
rect 34935 4440 34980 4468
rect 34149 4431 34207 4437
rect 34974 4428 34980 4440
rect 35032 4428 35038 4480
rect 35342 4428 35348 4480
rect 35400 4468 35406 4480
rect 35621 4471 35679 4477
rect 35621 4468 35633 4471
rect 35400 4440 35633 4468
rect 35400 4428 35406 4440
rect 35621 4437 35633 4440
rect 35667 4437 35679 4471
rect 35621 4431 35679 4437
rect 35986 4428 35992 4480
rect 36044 4468 36050 4480
rect 36265 4471 36323 4477
rect 36265 4468 36277 4471
rect 36044 4440 36277 4468
rect 36044 4428 36050 4440
rect 36265 4437 36277 4440
rect 36311 4437 36323 4471
rect 36265 4431 36323 4437
rect 36998 4428 37004 4480
rect 37056 4428 37062 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 15746 4264 15752 4276
rect 12912 4236 15752 4264
rect 11606 4156 11612 4208
rect 11664 4196 11670 4208
rect 12912 4205 12940 4236
rect 15746 4224 15752 4236
rect 15804 4224 15810 4276
rect 15930 4224 15936 4276
rect 15988 4264 15994 4276
rect 24670 4264 24676 4276
rect 15988 4236 24676 4264
rect 15988 4224 15994 4236
rect 24670 4224 24676 4236
rect 24728 4224 24734 4276
rect 33870 4264 33876 4276
rect 24872 4236 33876 4264
rect 12897 4199 12955 4205
rect 12897 4196 12909 4199
rect 11664 4168 12909 4196
rect 11664 4156 11670 4168
rect 12897 4165 12909 4168
rect 12943 4165 12955 4199
rect 14274 4196 14280 4208
rect 14235 4168 14280 4196
rect 12897 4159 12955 4165
rect 14274 4156 14280 4168
rect 14332 4156 14338 4208
rect 17954 4196 17960 4208
rect 16224 4168 17960 4196
rect 11149 4131 11207 4137
rect 11149 4097 11161 4131
rect 11195 4128 11207 4131
rect 11885 4131 11943 4137
rect 11885 4128 11897 4131
rect 11195 4100 11897 4128
rect 11195 4097 11207 4100
rect 11149 4091 11207 4097
rect 11885 4097 11897 4100
rect 11931 4128 11943 4131
rect 12437 4131 12495 4137
rect 12437 4128 12449 4131
rect 11931 4100 12449 4128
rect 11931 4097 11943 4100
rect 11885 4091 11943 4097
rect 12437 4097 12449 4100
rect 12483 4128 12495 4131
rect 13446 4128 13452 4140
rect 12483 4100 13452 4128
rect 12483 4097 12495 4100
rect 12437 4091 12495 4097
rect 13446 4088 13452 4100
rect 13504 4088 13510 4140
rect 15286 4128 15292 4140
rect 15199 4100 15292 4128
rect 15286 4088 15292 4100
rect 15344 4128 15350 4140
rect 15838 4128 15844 4140
rect 15344 4100 15844 4128
rect 15344 4088 15350 4100
rect 15838 4088 15844 4100
rect 15896 4088 15902 4140
rect 16114 4128 16120 4140
rect 16075 4100 16120 4128
rect 16114 4088 16120 4100
rect 16172 4088 16178 4140
rect 16224 4137 16252 4168
rect 17954 4156 17960 4168
rect 18012 4156 18018 4208
rect 18598 4156 18604 4208
rect 18656 4196 18662 4208
rect 21818 4196 21824 4208
rect 18656 4168 19748 4196
rect 21206 4168 21824 4196
rect 18656 4156 18662 4168
rect 16209 4131 16267 4137
rect 16209 4097 16221 4131
rect 16255 4097 16267 4131
rect 17034 4128 17040 4140
rect 16995 4100 17040 4128
rect 16209 4091 16267 4097
rect 17034 4088 17040 4100
rect 17092 4088 17098 4140
rect 17129 4131 17187 4137
rect 17129 4097 17141 4131
rect 17175 4128 17187 4131
rect 17310 4128 17316 4140
rect 17175 4100 17316 4128
rect 17175 4097 17187 4100
rect 17129 4091 17187 4097
rect 17310 4088 17316 4100
rect 17368 4088 17374 4140
rect 17586 4088 17592 4140
rect 17644 4137 17650 4140
rect 17644 4128 17655 4137
rect 18506 4128 18512 4140
rect 17644 4100 18512 4128
rect 17644 4091 17655 4100
rect 17644 4088 17650 4091
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 18782 4088 18788 4140
rect 18840 4128 18846 4140
rect 19242 4128 19248 4140
rect 18840 4100 19248 4128
rect 18840 4088 18846 4100
rect 19242 4088 19248 4100
rect 19300 4128 19306 4140
rect 19720 4137 19748 4168
rect 21818 4156 21824 4168
rect 21876 4156 21882 4208
rect 24872 4196 24900 4236
rect 33870 4224 33876 4236
rect 33928 4224 33934 4276
rect 36538 4264 36544 4276
rect 33980 4236 36544 4264
rect 23506 4168 24900 4196
rect 24946 4156 24952 4208
rect 25004 4156 25010 4208
rect 29546 4196 29552 4208
rect 29026 4168 29552 4196
rect 29546 4156 29552 4168
rect 29604 4156 29610 4208
rect 31294 4196 31300 4208
rect 30774 4168 31300 4196
rect 31294 4156 31300 4168
rect 31352 4156 31358 4208
rect 33980 4196 34008 4236
rect 36538 4224 36544 4236
rect 36596 4224 36602 4276
rect 33810 4168 34008 4196
rect 34882 4156 34888 4208
rect 34940 4196 34946 4208
rect 34940 4168 35848 4196
rect 34940 4156 34946 4168
rect 19705 4131 19763 4137
rect 19300 4100 19472 4128
rect 19300 4088 19306 4100
rect 12526 4020 12532 4072
rect 12584 4060 12590 4072
rect 14185 4063 14243 4069
rect 14185 4060 14197 4063
rect 12584 4032 14197 4060
rect 12584 4020 12590 4032
rect 14185 4029 14197 4032
rect 14231 4029 14243 4063
rect 14550 4060 14556 4072
rect 14511 4032 14556 4060
rect 14185 4023 14243 4029
rect 14550 4020 14556 4032
rect 14608 4020 14614 4072
rect 15381 4063 15439 4069
rect 15381 4029 15393 4063
rect 15427 4060 15439 4063
rect 16298 4060 16304 4072
rect 15427 4032 16304 4060
rect 15427 4029 15439 4032
rect 15381 4023 15439 4029
rect 16298 4020 16304 4032
rect 16356 4020 16362 4072
rect 16574 4020 16580 4072
rect 16632 4060 16638 4072
rect 17402 4060 17408 4072
rect 16632 4032 17408 4060
rect 16632 4020 16638 4032
rect 17402 4020 17408 4032
rect 17460 4020 17466 4072
rect 17678 4020 17684 4072
rect 17736 4060 17742 4072
rect 17736 4032 17781 4060
rect 17880 4032 19380 4060
rect 17736 4020 17742 4032
rect 13541 3995 13599 4001
rect 13541 3961 13553 3995
rect 13587 3961 13599 3995
rect 13541 3955 13599 3961
rect 13556 3924 13584 3955
rect 13630 3952 13636 4004
rect 13688 3992 13694 4004
rect 17880 3992 17908 4032
rect 19245 3995 19303 4001
rect 19245 3992 19257 3995
rect 13688 3964 17908 3992
rect 18616 3964 19257 3992
rect 13688 3952 13694 3964
rect 18616 3936 18644 3964
rect 19245 3961 19257 3964
rect 19291 3961 19303 3995
rect 19245 3955 19303 3961
rect 18046 3924 18052 3936
rect 13556 3896 18052 3924
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 18598 3924 18604 3936
rect 18559 3896 18604 3924
rect 18598 3884 18604 3896
rect 18656 3884 18662 3936
rect 19352 3924 19380 4032
rect 19444 3992 19472 4100
rect 19705 4097 19717 4131
rect 19751 4097 19763 4131
rect 22002 4128 22008 4140
rect 21963 4100 22008 4128
rect 19705 4091 19763 4097
rect 22002 4088 22008 4100
rect 22060 4088 22066 4140
rect 24210 4128 24216 4140
rect 24171 4100 24216 4128
rect 24210 4088 24216 4100
rect 24268 4088 24274 4140
rect 26418 4128 26424 4140
rect 26379 4100 26424 4128
rect 26418 4088 26424 4100
rect 26476 4088 26482 4140
rect 26510 4088 26516 4140
rect 26568 4128 26574 4140
rect 26568 4100 26613 4128
rect 29288 4100 30052 4128
rect 26568 4088 26574 4100
rect 19981 4063 20039 4069
rect 19981 4060 19993 4063
rect 19812 4032 19993 4060
rect 19812 3992 19840 4032
rect 19981 4029 19993 4032
rect 20027 4029 20039 4063
rect 19981 4023 20039 4029
rect 20714 4020 20720 4072
rect 20772 4060 20778 4072
rect 22281 4063 22339 4069
rect 22281 4060 22293 4063
rect 20772 4032 22293 4060
rect 20772 4020 20778 4032
rect 21468 4001 21496 4032
rect 22281 4029 22293 4032
rect 22327 4029 22339 4063
rect 22281 4023 22339 4029
rect 22370 4020 22376 4072
rect 22428 4060 22434 4072
rect 24486 4060 24492 4072
rect 22428 4032 24348 4060
rect 24447 4032 24492 4060
rect 22428 4020 22434 4032
rect 19444 3964 19840 3992
rect 21453 3995 21511 4001
rect 21453 3961 21465 3995
rect 21499 3992 21511 3995
rect 21499 3964 21533 3992
rect 21499 3961 21511 3964
rect 21453 3955 21511 3961
rect 23658 3952 23664 4004
rect 23716 3992 23722 4004
rect 23753 3995 23811 4001
rect 23753 3992 23765 3995
rect 23716 3964 23765 3992
rect 23716 3952 23722 3964
rect 23753 3961 23765 3964
rect 23799 3992 23811 3995
rect 24210 3992 24216 4004
rect 23799 3964 24216 3992
rect 23799 3961 23811 3964
rect 23753 3955 23811 3961
rect 24210 3952 24216 3964
rect 24268 3952 24274 4004
rect 22094 3924 22100 3936
rect 19352 3896 22100 3924
rect 22094 3884 22100 3896
rect 22152 3884 22158 3936
rect 22462 3884 22468 3936
rect 22520 3924 22526 3936
rect 24026 3924 24032 3936
rect 22520 3896 24032 3924
rect 22520 3884 22526 3896
rect 24026 3884 24032 3896
rect 24084 3884 24090 3936
rect 24320 3924 24348 4032
rect 24486 4020 24492 4032
rect 24544 4020 24550 4072
rect 26326 4020 26332 4072
rect 26384 4060 26390 4072
rect 27430 4060 27436 4072
rect 26384 4032 27436 4060
rect 26384 4020 26390 4032
rect 27430 4020 27436 4032
rect 27488 4060 27494 4072
rect 27525 4063 27583 4069
rect 27525 4060 27537 4063
rect 27488 4032 27537 4060
rect 27488 4020 27494 4032
rect 27525 4029 27537 4032
rect 27571 4029 27583 4063
rect 27525 4023 27583 4029
rect 27801 4063 27859 4069
rect 27801 4029 27813 4063
rect 27847 4060 27859 4063
rect 29288 4060 29316 4100
rect 27847 4032 29316 4060
rect 27847 4029 27859 4032
rect 27801 4023 27859 4029
rect 29362 4020 29368 4072
rect 29420 4060 29426 4072
rect 29733 4063 29791 4069
rect 29733 4060 29745 4063
rect 29420 4032 29745 4060
rect 29420 4020 29426 4032
rect 29733 4029 29745 4032
rect 29779 4029 29791 4063
rect 30024 4060 30052 4100
rect 31478 4088 31484 4140
rect 31536 4128 31542 4140
rect 31662 4128 31668 4140
rect 31536 4100 31668 4128
rect 31536 4088 31542 4100
rect 31662 4088 31668 4100
rect 31720 4128 31726 4140
rect 31720 4088 31754 4128
rect 33870 4088 33876 4140
rect 33928 4128 33934 4140
rect 34606 4128 34612 4140
rect 33928 4100 34612 4128
rect 33928 4088 33934 4100
rect 34606 4088 34612 4100
rect 34664 4088 34670 4140
rect 34701 4131 34759 4137
rect 34701 4097 34713 4131
rect 34747 4126 34759 4131
rect 34900 4126 34928 4156
rect 35820 4140 35848 4168
rect 36354 4156 36360 4208
rect 36412 4196 36418 4208
rect 36412 4168 36768 4196
rect 36412 4156 36418 4168
rect 34747 4098 34928 4126
rect 34747 4097 34759 4098
rect 34701 4091 34759 4097
rect 34974 4088 34980 4140
rect 35032 4128 35038 4140
rect 35345 4131 35403 4137
rect 35345 4128 35357 4131
rect 35032 4100 35357 4128
rect 35032 4088 35038 4100
rect 35345 4097 35357 4100
rect 35391 4128 35403 4131
rect 35434 4128 35440 4140
rect 35391 4100 35440 4128
rect 35391 4097 35403 4100
rect 35345 4091 35403 4097
rect 35434 4088 35440 4100
rect 35492 4088 35498 4140
rect 35802 4088 35808 4140
rect 35860 4128 35866 4140
rect 35989 4131 36047 4137
rect 35989 4128 36001 4131
rect 35860 4100 36001 4128
rect 35860 4088 35866 4100
rect 35989 4097 36001 4100
rect 36035 4128 36047 4131
rect 36633 4131 36691 4137
rect 36633 4128 36645 4131
rect 36035 4100 36645 4128
rect 36035 4097 36047 4100
rect 35989 4091 36047 4097
rect 36633 4097 36645 4100
rect 36679 4097 36691 4131
rect 36740 4128 36768 4168
rect 37645 4131 37703 4137
rect 37645 4128 37657 4131
rect 36740 4100 37657 4128
rect 36633 4091 36691 4097
rect 37645 4097 37657 4100
rect 37691 4097 37703 4131
rect 37645 4091 37703 4097
rect 38105 4131 38163 4137
rect 38105 4097 38117 4131
rect 38151 4097 38163 4131
rect 38105 4091 38163 4097
rect 30742 4060 30748 4072
rect 30024 4032 30748 4060
rect 29733 4023 29791 4029
rect 30742 4020 30748 4032
rect 30800 4020 30806 4072
rect 30834 4020 30840 4072
rect 30892 4060 30898 4072
rect 31110 4060 31116 4072
rect 30892 4032 31116 4060
rect 30892 4020 30898 4032
rect 31110 4020 31116 4032
rect 31168 4060 31174 4072
rect 31205 4063 31263 4069
rect 31205 4060 31217 4063
rect 31168 4032 31217 4060
rect 31168 4020 31174 4032
rect 31205 4029 31217 4032
rect 31251 4029 31263 4063
rect 31726 4060 31754 4088
rect 32309 4063 32367 4069
rect 32309 4060 32321 4063
rect 31726 4032 32321 4060
rect 31205 4023 31263 4029
rect 32309 4029 32321 4032
rect 32355 4029 32367 4063
rect 32582 4060 32588 4072
rect 32309 4023 32367 4029
rect 32416 4032 32588 4060
rect 26142 3952 26148 4004
rect 26200 3992 26206 4004
rect 26418 3992 26424 4004
rect 26200 3964 26424 3992
rect 26200 3952 26206 3964
rect 26418 3952 26424 3964
rect 26476 3952 26482 4004
rect 28810 3952 28816 4004
rect 28868 3992 28874 4004
rect 28868 3964 29408 3992
rect 28868 3952 28874 3964
rect 25958 3924 25964 3936
rect 24320 3896 25964 3924
rect 25958 3884 25964 3896
rect 26016 3884 26022 3936
rect 26694 3884 26700 3936
rect 26752 3924 26758 3936
rect 28994 3924 29000 3936
rect 26752 3896 29000 3924
rect 26752 3884 26758 3896
rect 28994 3884 29000 3896
rect 29052 3884 29058 3936
rect 29270 3924 29276 3936
rect 29231 3896 29276 3924
rect 29270 3884 29276 3896
rect 29328 3884 29334 3936
rect 29380 3924 29408 3964
rect 32122 3952 32128 4004
rect 32180 3992 32186 4004
rect 32416 3992 32444 4032
rect 32582 4020 32588 4032
rect 32640 4020 32646 4072
rect 33134 4020 33140 4072
rect 33192 4060 33198 4072
rect 37553 4063 37611 4069
rect 37553 4060 37565 4063
rect 33192 4032 37565 4060
rect 33192 4020 33198 4032
rect 37553 4029 37565 4032
rect 37599 4029 37611 4063
rect 37553 4023 37611 4029
rect 32180 3964 32444 3992
rect 32180 3952 32186 3964
rect 34514 3952 34520 4004
rect 34572 3992 34578 4004
rect 36541 3995 36599 4001
rect 36541 3992 36553 3995
rect 34572 3964 36553 3992
rect 34572 3952 34578 3964
rect 36541 3961 36553 3964
rect 36587 3961 36599 3995
rect 36541 3955 36599 3961
rect 36630 3952 36636 4004
rect 36688 3992 36694 4004
rect 37642 3992 37648 4004
rect 36688 3964 37648 3992
rect 36688 3952 36694 3964
rect 37642 3952 37648 3964
rect 37700 3992 37706 4004
rect 38120 3992 38148 4091
rect 37700 3964 38148 3992
rect 37700 3952 37706 3964
rect 33778 3924 33784 3936
rect 29380 3896 33784 3924
rect 33778 3884 33784 3896
rect 33836 3884 33842 3936
rect 33870 3884 33876 3936
rect 33928 3924 33934 3936
rect 34057 3927 34115 3933
rect 34057 3924 34069 3927
rect 33928 3896 34069 3924
rect 33928 3884 33934 3896
rect 34057 3893 34069 3896
rect 34103 3893 34115 3927
rect 34057 3887 34115 3893
rect 34146 3884 34152 3936
rect 34204 3924 34210 3936
rect 34609 3927 34667 3933
rect 34609 3924 34621 3927
rect 34204 3896 34621 3924
rect 34204 3884 34210 3896
rect 34609 3893 34621 3896
rect 34655 3893 34667 3927
rect 34609 3887 34667 3893
rect 34698 3884 34704 3936
rect 34756 3924 34762 3936
rect 35253 3927 35311 3933
rect 35253 3924 35265 3927
rect 34756 3896 35265 3924
rect 34756 3884 34762 3896
rect 35253 3893 35265 3896
rect 35299 3893 35311 3927
rect 35894 3924 35900 3936
rect 35855 3896 35900 3924
rect 35253 3887 35311 3893
rect 35894 3884 35900 3896
rect 35952 3884 35958 3936
rect 36170 3884 36176 3936
rect 36228 3924 36234 3936
rect 38197 3927 38255 3933
rect 38197 3924 38209 3927
rect 36228 3896 38209 3924
rect 36228 3884 36234 3896
rect 38197 3893 38209 3896
rect 38243 3893 38255 3927
rect 38197 3887 38255 3893
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 2314 3720 2320 3732
rect 2275 3692 2320 3720
rect 2314 3680 2320 3692
rect 2372 3680 2378 3732
rect 10597 3723 10655 3729
rect 10597 3689 10609 3723
rect 10643 3720 10655 3723
rect 10962 3720 10968 3732
rect 10643 3692 10968 3720
rect 10643 3689 10655 3692
rect 10597 3683 10655 3689
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 11606 3720 11612 3732
rect 11567 3692 11612 3720
rect 11606 3680 11612 3692
rect 11664 3680 11670 3732
rect 12250 3720 12256 3732
rect 12211 3692 12256 3720
rect 12250 3680 12256 3692
rect 12308 3680 12314 3732
rect 13633 3723 13691 3729
rect 13633 3689 13645 3723
rect 13679 3720 13691 3723
rect 14274 3720 14280 3732
rect 13679 3692 14280 3720
rect 13679 3689 13691 3692
rect 13633 3683 13691 3689
rect 14274 3680 14280 3692
rect 14332 3680 14338 3732
rect 14384 3692 21864 3720
rect 14182 3612 14188 3664
rect 14240 3652 14246 3664
rect 14384 3652 14412 3692
rect 14240 3624 14412 3652
rect 14568 3624 20668 3652
rect 14240 3612 14246 3624
rect 12176 3556 12848 3584
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3516 1915 3519
rect 2774 3516 2780 3528
rect 1903 3488 2780 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 2774 3476 2780 3488
rect 2832 3476 2838 3528
rect 11790 3476 11796 3528
rect 11848 3516 11854 3528
rect 12176 3525 12204 3556
rect 12161 3519 12219 3525
rect 12161 3516 12173 3519
rect 11848 3488 12173 3516
rect 11848 3476 11854 3488
rect 12161 3485 12173 3488
rect 12207 3485 12219 3519
rect 12161 3479 12219 3485
rect 11149 3451 11207 3457
rect 11149 3417 11161 3451
rect 11195 3448 11207 3451
rect 12820 3448 12848 3556
rect 12894 3544 12900 3596
rect 12952 3584 12958 3596
rect 12952 3556 14504 3584
rect 12952 3544 12958 3556
rect 12986 3476 12992 3528
rect 13044 3516 13050 3528
rect 13541 3519 13599 3525
rect 13541 3516 13553 3519
rect 13044 3488 13553 3516
rect 13044 3476 13050 3488
rect 13541 3485 13553 3488
rect 13587 3516 13599 3519
rect 13722 3516 13728 3528
rect 13587 3488 13728 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 14274 3516 14280 3528
rect 14235 3488 14280 3516
rect 14274 3476 14280 3488
rect 14332 3476 14338 3528
rect 14292 3448 14320 3476
rect 11195 3420 12434 3448
rect 12820 3420 14320 3448
rect 14476 3448 14504 3556
rect 14568 3525 14596 3624
rect 17494 3584 17500 3596
rect 15212 3556 17500 3584
rect 14553 3519 14611 3525
rect 14553 3485 14565 3519
rect 14599 3485 14611 3519
rect 14553 3479 14611 3485
rect 15212 3457 15240 3556
rect 17494 3544 17500 3556
rect 17552 3584 17558 3596
rect 18598 3584 18604 3596
rect 17552 3556 18604 3584
rect 17552 3544 17558 3556
rect 18598 3544 18604 3556
rect 18656 3584 18662 3596
rect 19150 3584 19156 3596
rect 18656 3556 19156 3584
rect 18656 3544 18662 3556
rect 19150 3544 19156 3556
rect 19208 3584 19214 3596
rect 20533 3587 20591 3593
rect 20533 3584 20545 3587
rect 19208 3556 20545 3584
rect 19208 3544 19214 3556
rect 20533 3553 20545 3556
rect 20579 3553 20591 3587
rect 20640 3584 20668 3624
rect 21542 3584 21548 3596
rect 20640 3556 21548 3584
rect 20533 3547 20591 3553
rect 21542 3544 21548 3556
rect 21600 3544 21606 3596
rect 21836 3584 21864 3692
rect 22094 3680 22100 3732
rect 22152 3720 22158 3732
rect 23014 3720 23020 3732
rect 22152 3692 23020 3720
rect 22152 3680 22158 3692
rect 23014 3680 23020 3692
rect 23072 3680 23078 3732
rect 23198 3720 23204 3732
rect 23159 3692 23204 3720
rect 23198 3680 23204 3692
rect 23256 3680 23262 3732
rect 28810 3720 28816 3732
rect 24044 3692 28816 3720
rect 21910 3612 21916 3664
rect 21968 3652 21974 3664
rect 21968 3624 23152 3652
rect 21968 3612 21974 3624
rect 22922 3584 22928 3596
rect 21836 3556 22928 3584
rect 22922 3544 22928 3556
rect 22980 3544 22986 3596
rect 17126 3476 17132 3528
rect 17184 3516 17190 3528
rect 17184 3488 17229 3516
rect 17184 3476 17190 3488
rect 17402 3476 17408 3528
rect 17460 3516 17466 3528
rect 17589 3519 17647 3525
rect 17589 3516 17601 3519
rect 17460 3488 17601 3516
rect 17460 3476 17466 3488
rect 17589 3485 17601 3488
rect 17635 3485 17647 3519
rect 17862 3516 17868 3528
rect 17823 3488 17868 3516
rect 17589 3479 17647 3485
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 18506 3516 18512 3528
rect 18419 3488 18512 3516
rect 18506 3476 18512 3488
rect 18564 3516 18570 3528
rect 23124 3525 23152 3624
rect 23109 3519 23167 3525
rect 18564 3488 19748 3516
rect 18564 3476 18570 3488
rect 15197 3451 15255 3457
rect 15197 3448 15209 3451
rect 14476 3420 15209 3448
rect 11195 3417 11207 3420
rect 11149 3411 11207 3417
rect 1670 3380 1676 3392
rect 1631 3352 1676 3380
rect 1670 3340 1676 3352
rect 1728 3340 1734 3392
rect 12406 3380 12434 3420
rect 15197 3417 15209 3420
rect 15243 3417 15255 3451
rect 15197 3411 15255 3417
rect 15933 3451 15991 3457
rect 15933 3417 15945 3451
rect 15979 3448 15991 3451
rect 16485 3451 16543 3457
rect 16485 3448 16497 3451
rect 15979 3420 16497 3448
rect 15979 3417 15991 3420
rect 15933 3411 15991 3417
rect 16485 3417 16497 3420
rect 16531 3417 16543 3451
rect 16485 3411 16543 3417
rect 16577 3451 16635 3457
rect 16577 3417 16589 3451
rect 16623 3448 16635 3451
rect 16942 3448 16948 3460
rect 16623 3420 16948 3448
rect 16623 3417 16635 3420
rect 16577 3411 16635 3417
rect 16942 3408 16948 3420
rect 17000 3408 17006 3460
rect 18138 3408 18144 3460
rect 18196 3448 18202 3460
rect 18690 3448 18696 3460
rect 18196 3420 18696 3448
rect 18196 3408 18202 3420
rect 18690 3408 18696 3420
rect 18748 3448 18754 3460
rect 19613 3451 19671 3457
rect 19613 3448 19625 3451
rect 18748 3420 19625 3448
rect 18748 3408 18754 3420
rect 19613 3417 19625 3420
rect 19659 3417 19671 3451
rect 19613 3411 19671 3417
rect 12986 3380 12992 3392
rect 12406 3352 12992 3380
rect 12986 3340 12992 3352
rect 13044 3340 13050 3392
rect 13081 3383 13139 3389
rect 13081 3349 13093 3383
rect 13127 3380 13139 3383
rect 16758 3380 16764 3392
rect 13127 3352 16764 3380
rect 13127 3349 13139 3352
rect 13081 3343 13139 3349
rect 16758 3340 16764 3352
rect 16816 3340 16822 3392
rect 18601 3383 18659 3389
rect 18601 3349 18613 3383
rect 18647 3380 18659 3383
rect 18874 3380 18880 3392
rect 18647 3352 18880 3380
rect 18647 3349 18659 3352
rect 18601 3343 18659 3349
rect 18874 3340 18880 3352
rect 18932 3340 18938 3392
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 19521 3383 19579 3389
rect 19521 3380 19533 3383
rect 19484 3352 19533 3380
rect 19484 3340 19490 3352
rect 19521 3349 19533 3352
rect 19567 3349 19579 3383
rect 19720 3380 19748 3488
rect 23109 3485 23121 3519
rect 23155 3516 23167 3519
rect 23934 3516 23940 3528
rect 23155 3488 23940 3516
rect 23155 3485 23167 3488
rect 23109 3479 23167 3485
rect 23934 3476 23940 3488
rect 23992 3476 23998 3528
rect 24044 3525 24072 3692
rect 28810 3680 28816 3692
rect 28868 3680 28874 3732
rect 29181 3723 29239 3729
rect 29181 3689 29193 3723
rect 29227 3720 29239 3723
rect 31662 3720 31668 3732
rect 29227 3692 31668 3720
rect 29227 3689 29239 3692
rect 29181 3683 29239 3689
rect 31662 3680 31668 3692
rect 31720 3680 31726 3732
rect 31938 3720 31944 3732
rect 31899 3692 31944 3720
rect 31938 3680 31944 3692
rect 31996 3680 32002 3732
rect 32030 3680 32036 3732
rect 32088 3720 32094 3732
rect 33226 3720 33232 3732
rect 32088 3692 33232 3720
rect 32088 3680 32094 3692
rect 33226 3680 33232 3692
rect 33284 3680 33290 3732
rect 34238 3720 34244 3732
rect 34199 3692 34244 3720
rect 34238 3680 34244 3692
rect 34296 3680 34302 3732
rect 26418 3612 26424 3664
rect 26476 3652 26482 3664
rect 27525 3655 27583 3661
rect 27525 3652 27537 3655
rect 26476 3624 27537 3652
rect 26476 3612 26482 3624
rect 27525 3621 27537 3624
rect 27571 3621 27583 3655
rect 27525 3615 27583 3621
rect 27890 3612 27896 3664
rect 27948 3652 27954 3664
rect 29638 3652 29644 3664
rect 27948 3624 29644 3652
rect 27948 3612 27954 3624
rect 29638 3612 29644 3624
rect 29696 3612 29702 3664
rect 29733 3655 29791 3661
rect 29733 3621 29745 3655
rect 29779 3652 29791 3655
rect 29914 3652 29920 3664
rect 29779 3624 29920 3652
rect 29779 3621 29791 3624
rect 29733 3615 29791 3621
rect 29914 3612 29920 3624
rect 29972 3612 29978 3664
rect 31570 3612 31576 3664
rect 31628 3652 31634 3664
rect 32306 3652 32312 3664
rect 31628 3624 32312 3652
rect 31628 3612 31634 3624
rect 32306 3612 32312 3624
rect 32364 3612 32370 3664
rect 33778 3612 33784 3664
rect 33836 3652 33842 3664
rect 36814 3652 36820 3664
rect 33836 3624 36820 3652
rect 33836 3612 33842 3624
rect 36814 3612 36820 3624
rect 36872 3612 36878 3664
rect 24302 3544 24308 3596
rect 24360 3584 24366 3596
rect 24578 3584 24584 3596
rect 24360 3556 24584 3584
rect 24360 3544 24366 3556
rect 24578 3544 24584 3556
rect 24636 3584 24642 3596
rect 25041 3587 25099 3593
rect 25041 3584 25053 3587
rect 24636 3556 25053 3584
rect 24636 3544 24642 3556
rect 25041 3553 25053 3556
rect 25087 3584 25099 3587
rect 26326 3584 26332 3596
rect 25087 3556 26332 3584
rect 25087 3553 25099 3556
rect 25041 3547 25099 3553
rect 26326 3544 26332 3556
rect 26384 3544 26390 3596
rect 26510 3544 26516 3596
rect 26568 3584 26574 3596
rect 31202 3584 31208 3596
rect 26568 3556 31208 3584
rect 26568 3544 26574 3556
rect 31202 3544 31208 3556
rect 31260 3544 31266 3596
rect 31478 3584 31484 3596
rect 31439 3556 31484 3584
rect 31478 3544 31484 3556
rect 31536 3584 31542 3596
rect 33689 3587 33747 3593
rect 33689 3584 33701 3587
rect 31536 3556 33701 3584
rect 31536 3544 31542 3556
rect 33689 3553 33701 3556
rect 33735 3584 33747 3587
rect 34054 3584 34060 3596
rect 33735 3556 34060 3584
rect 33735 3553 33747 3556
rect 33689 3547 33747 3553
rect 34054 3544 34060 3556
rect 34112 3584 34118 3596
rect 37550 3584 37556 3596
rect 34112 3556 37556 3584
rect 34112 3544 34118 3556
rect 37550 3544 37556 3556
rect 37608 3544 37614 3596
rect 24029 3519 24087 3525
rect 24029 3485 24041 3519
rect 24075 3485 24087 3519
rect 24029 3479 24087 3485
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 28994 3516 29000 3528
rect 24268 3488 24992 3516
rect 24268 3476 24274 3488
rect 19978 3408 19984 3460
rect 20036 3448 20042 3460
rect 20809 3451 20867 3457
rect 20809 3448 20821 3451
rect 20036 3420 20821 3448
rect 20036 3408 20042 3420
rect 20809 3417 20821 3420
rect 20855 3448 20867 3451
rect 20898 3448 20904 3460
rect 20855 3420 20904 3448
rect 20855 3417 20867 3420
rect 20809 3411 20867 3417
rect 20898 3408 20904 3420
rect 20956 3408 20962 3460
rect 22186 3448 22192 3460
rect 22034 3420 22192 3448
rect 22186 3408 22192 3420
rect 22244 3408 22250 3460
rect 22554 3448 22560 3460
rect 22515 3420 22560 3448
rect 22554 3408 22560 3420
rect 22612 3408 22618 3460
rect 24964 3448 24992 3488
rect 26988 3488 28304 3516
rect 28907 3488 29000 3516
rect 25317 3451 25375 3457
rect 25317 3448 25329 3451
rect 24964 3420 25329 3448
rect 25317 3417 25329 3420
rect 25363 3417 25375 3451
rect 26988 3448 27016 3488
rect 26542 3420 27016 3448
rect 25317 3411 25375 3417
rect 27062 3408 27068 3460
rect 27120 3448 27126 3460
rect 27120 3420 27165 3448
rect 27120 3408 27126 3420
rect 27246 3408 27252 3460
rect 27304 3448 27310 3460
rect 28276 3448 28304 3488
rect 28994 3476 29000 3488
rect 29052 3516 29058 3528
rect 29822 3516 29828 3528
rect 29052 3488 29828 3516
rect 29052 3476 29058 3488
rect 29822 3476 29828 3488
rect 29880 3476 29886 3528
rect 34238 3476 34244 3528
rect 34296 3516 34302 3528
rect 34333 3519 34391 3525
rect 34333 3516 34345 3519
rect 34296 3488 34345 3516
rect 34296 3476 34302 3488
rect 34333 3485 34345 3488
rect 34379 3516 34391 3519
rect 35069 3519 35127 3525
rect 35069 3516 35081 3519
rect 34379 3488 35081 3516
rect 34379 3485 34391 3488
rect 34333 3479 34391 3485
rect 35069 3485 35081 3488
rect 35115 3516 35127 3519
rect 35713 3519 35771 3525
rect 35713 3516 35725 3519
rect 35115 3488 35725 3516
rect 35115 3485 35127 3488
rect 35069 3479 35127 3485
rect 35713 3485 35725 3488
rect 35759 3516 35771 3519
rect 36357 3519 36415 3525
rect 36357 3516 36369 3519
rect 35759 3488 36369 3516
rect 35759 3485 35771 3488
rect 35713 3479 35771 3485
rect 36357 3485 36369 3488
rect 36403 3516 36415 3519
rect 36630 3516 36636 3528
rect 36403 3488 36636 3516
rect 36403 3485 36415 3488
rect 36357 3479 36415 3485
rect 36630 3476 36636 3488
rect 36688 3476 36694 3528
rect 36814 3516 36820 3528
rect 36775 3488 36820 3516
rect 36814 3476 36820 3488
rect 36872 3476 36878 3528
rect 38013 3519 38071 3525
rect 38013 3516 38025 3519
rect 37016 3488 38025 3516
rect 27304 3420 28212 3448
rect 28276 3420 29868 3448
rect 30774 3420 30880 3448
rect 27304 3408 27310 3420
rect 21174 3380 21180 3392
rect 19720 3352 21180 3380
rect 19521 3343 19579 3349
rect 21174 3340 21180 3352
rect 21232 3340 21238 3392
rect 23842 3380 23848 3392
rect 23803 3352 23848 3380
rect 23842 3340 23848 3352
rect 23900 3340 23906 3392
rect 23934 3340 23940 3392
rect 23992 3380 23998 3392
rect 26694 3380 26700 3392
rect 23992 3352 26700 3380
rect 23992 3340 23998 3352
rect 26694 3340 26700 3352
rect 26752 3340 26758 3392
rect 28074 3380 28080 3392
rect 28035 3352 28080 3380
rect 28074 3340 28080 3352
rect 28132 3340 28138 3392
rect 28184 3380 28212 3420
rect 29730 3380 29736 3392
rect 28184 3352 29736 3380
rect 29730 3340 29736 3352
rect 29788 3340 29794 3392
rect 29840 3380 29868 3420
rect 30558 3380 30564 3392
rect 29840 3352 30564 3380
rect 30558 3340 30564 3352
rect 30616 3340 30622 3392
rect 30852 3380 30880 3420
rect 30926 3408 30932 3460
rect 30984 3448 30990 3460
rect 31205 3451 31263 3457
rect 31205 3448 31217 3451
rect 30984 3420 31217 3448
rect 30984 3408 30990 3420
rect 31205 3417 31217 3420
rect 31251 3417 31263 3451
rect 31205 3411 31263 3417
rect 31294 3408 31300 3460
rect 31352 3448 31358 3460
rect 31570 3448 31576 3460
rect 31352 3420 31576 3448
rect 31352 3408 31358 3420
rect 31570 3408 31576 3420
rect 31628 3408 31634 3460
rect 33318 3448 33324 3460
rect 31726 3420 32076 3448
rect 32982 3420 33324 3448
rect 31726 3380 31754 3420
rect 30852 3352 31754 3380
rect 32048 3380 32076 3420
rect 33318 3408 33324 3420
rect 33376 3408 33382 3460
rect 33410 3408 33416 3460
rect 33468 3448 33474 3460
rect 33870 3448 33876 3460
rect 33468 3420 33876 3448
rect 33468 3408 33474 3420
rect 33870 3408 33876 3420
rect 33928 3408 33934 3460
rect 35986 3448 35992 3460
rect 33980 3420 35992 3448
rect 33980 3380 34008 3420
rect 35986 3408 35992 3420
rect 36044 3408 36050 3460
rect 34974 3380 34980 3392
rect 32048 3352 34008 3380
rect 34935 3352 34980 3380
rect 34974 3340 34980 3352
rect 35032 3340 35038 3392
rect 35618 3380 35624 3392
rect 35579 3352 35624 3380
rect 35618 3340 35624 3352
rect 35676 3340 35682 3392
rect 36262 3380 36268 3392
rect 36223 3352 36268 3380
rect 36262 3340 36268 3352
rect 36320 3340 36326 3392
rect 37016 3389 37044 3488
rect 38013 3485 38025 3488
rect 38059 3485 38071 3519
rect 38013 3479 38071 3485
rect 37001 3383 37059 3389
rect 37001 3349 37013 3383
rect 37047 3349 37059 3383
rect 37550 3380 37556 3392
rect 37511 3352 37556 3380
rect 37001 3343 37059 3349
rect 37550 3340 37556 3352
rect 37608 3340 37614 3392
rect 38194 3380 38200 3392
rect 38155 3352 38200 3380
rect 38194 3340 38200 3352
rect 38252 3340 38258 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 5077 3179 5135 3185
rect 5077 3145 5089 3179
rect 5123 3145 5135 3179
rect 5077 3139 5135 3145
rect 11149 3179 11207 3185
rect 11149 3145 11161 3179
rect 11195 3176 11207 3179
rect 11606 3176 11612 3188
rect 11195 3148 11612 3176
rect 11195 3145 11207 3148
rect 11149 3139 11207 3145
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 2314 3040 2320 3052
rect 1903 3012 2320 3040
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 2314 3000 2320 3012
rect 2372 3000 2378 3052
rect 2593 3043 2651 3049
rect 2593 3009 2605 3043
rect 2639 3040 2651 3043
rect 5092 3040 5120 3139
rect 11606 3136 11612 3148
rect 11664 3136 11670 3188
rect 12526 3176 12532 3188
rect 12487 3148 12532 3176
rect 12526 3136 12532 3148
rect 12584 3136 12590 3188
rect 15289 3179 15347 3185
rect 15289 3145 15301 3179
rect 15335 3176 15347 3179
rect 16574 3176 16580 3188
rect 15335 3148 16580 3176
rect 15335 3145 15347 3148
rect 15289 3139 15347 3145
rect 16574 3136 16580 3148
rect 16632 3136 16638 3188
rect 16942 3176 16948 3188
rect 16903 3148 16948 3176
rect 16942 3136 16948 3148
rect 17000 3136 17006 3188
rect 21266 3176 21272 3188
rect 17052 3148 21272 3176
rect 10594 3108 10600 3120
rect 10507 3080 10600 3108
rect 10594 3068 10600 3080
rect 10652 3108 10658 3120
rect 13357 3111 13415 3117
rect 10652 3080 12480 3108
rect 10652 3068 10658 3080
rect 12452 3052 12480 3080
rect 13357 3077 13369 3111
rect 13403 3108 13415 3111
rect 13630 3108 13636 3120
rect 13403 3080 13636 3108
rect 13403 3077 13415 3080
rect 13357 3071 13415 3077
rect 13630 3068 13636 3080
rect 13688 3068 13694 3120
rect 16114 3108 16120 3120
rect 15212 3080 16120 3108
rect 2639 3012 5120 3040
rect 5261 3043 5319 3049
rect 2639 3009 2651 3012
rect 2593 3003 2651 3009
rect 5261 3009 5273 3043
rect 5307 3040 5319 3043
rect 10042 3040 10048 3052
rect 5307 3012 10048 3040
rect 5307 3009 5319 3012
rect 5261 3003 5319 3009
rect 10042 3000 10048 3012
rect 10100 3000 10106 3052
rect 11790 3040 11796 3052
rect 11751 3012 11796 3040
rect 11790 3000 11796 3012
rect 11848 3000 11854 3052
rect 12434 3040 12440 3052
rect 12395 3012 12440 3040
rect 12434 3000 12440 3012
rect 12492 3000 12498 3052
rect 13081 3043 13139 3049
rect 13081 3009 13093 3043
rect 13127 3040 13139 3043
rect 13998 3040 14004 3052
rect 13127 3012 14004 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 13998 3000 14004 3012
rect 14056 3040 14062 3052
rect 14274 3040 14280 3052
rect 14056 3012 14280 3040
rect 14056 3000 14062 3012
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 15212 3049 15240 3080
rect 16114 3068 16120 3080
rect 16172 3068 16178 3120
rect 15197 3043 15255 3049
rect 15197 3009 15209 3043
rect 15243 3009 15255 3043
rect 15197 3003 15255 3009
rect 15746 3000 15752 3052
rect 15804 3040 15810 3052
rect 17052 3049 17080 3148
rect 21266 3136 21272 3148
rect 21324 3136 21330 3188
rect 21358 3136 21364 3188
rect 21416 3176 21422 3188
rect 21453 3179 21511 3185
rect 21453 3176 21465 3179
rect 21416 3148 21465 3176
rect 21416 3136 21422 3148
rect 21453 3145 21465 3148
rect 21499 3145 21511 3179
rect 21453 3139 21511 3145
rect 22186 3136 22192 3188
rect 22244 3176 22250 3188
rect 28074 3176 28080 3188
rect 22244 3148 28080 3176
rect 22244 3136 22250 3148
rect 17770 3108 17776 3120
rect 17731 3080 17776 3108
rect 17770 3068 17776 3080
rect 17828 3068 17834 3120
rect 19058 3108 19064 3120
rect 18998 3080 19064 3108
rect 19058 3068 19064 3080
rect 19116 3068 19122 3120
rect 19981 3111 20039 3117
rect 19981 3077 19993 3111
rect 20027 3108 20039 3111
rect 20254 3108 20260 3120
rect 20027 3080 20260 3108
rect 20027 3077 20039 3080
rect 19981 3071 20039 3077
rect 20254 3068 20260 3080
rect 20312 3068 20318 3120
rect 24026 3068 24032 3120
rect 24084 3108 24090 3120
rect 24857 3111 24915 3117
rect 24857 3108 24869 3111
rect 24084 3080 24869 3108
rect 24084 3068 24090 3080
rect 24857 3077 24869 3080
rect 24903 3077 24915 3111
rect 27798 3108 27804 3120
rect 26082 3080 27804 3108
rect 24857 3071 24915 3077
rect 27798 3068 27804 3080
rect 27856 3068 27862 3120
rect 27908 3117 27936 3148
rect 28074 3136 28080 3148
rect 28132 3136 28138 3188
rect 29270 3136 29276 3188
rect 29328 3176 29334 3188
rect 29328 3148 31754 3176
rect 29328 3136 29334 3148
rect 27893 3111 27951 3117
rect 27893 3077 27905 3111
rect 27939 3077 27951 3111
rect 27893 3071 27951 3077
rect 28902 3068 28908 3120
rect 28960 3068 28966 3120
rect 29362 3068 29368 3120
rect 29420 3108 29426 3120
rect 29641 3111 29699 3117
rect 29641 3108 29653 3111
rect 29420 3080 29653 3108
rect 29420 3068 29426 3080
rect 29641 3077 29653 3080
rect 29687 3077 29699 3111
rect 29641 3071 29699 3077
rect 29730 3068 29736 3120
rect 29788 3108 29794 3120
rect 31478 3108 31484 3120
rect 29788 3080 31484 3108
rect 29788 3068 29794 3080
rect 16209 3043 16267 3049
rect 16209 3040 16221 3043
rect 15804 3012 16221 3040
rect 15804 3000 15810 3012
rect 16209 3009 16221 3012
rect 16255 3009 16267 3043
rect 16209 3003 16267 3009
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3009 17095 3043
rect 17494 3040 17500 3052
rect 17455 3012 17500 3040
rect 17037 3003 17095 3009
rect 14182 2972 14188 2984
rect 14143 2944 14188 2972
rect 14182 2932 14188 2944
rect 14240 2932 14246 2984
rect 14292 2972 14320 3000
rect 15933 2975 15991 2981
rect 15933 2972 15945 2975
rect 14292 2944 15945 2972
rect 15933 2941 15945 2944
rect 15979 2941 15991 2975
rect 16224 2972 16252 3003
rect 17494 3000 17500 3012
rect 17552 3000 17558 3052
rect 19150 3000 19156 3052
rect 19208 3040 19214 3052
rect 19705 3043 19763 3049
rect 19705 3040 19717 3043
rect 19208 3012 19717 3040
rect 19208 3000 19214 3012
rect 19705 3009 19717 3012
rect 19751 3009 19763 3043
rect 19705 3003 19763 3009
rect 21082 3000 21088 3052
rect 21140 3000 21146 3052
rect 22002 3040 22008 3052
rect 21963 3012 22008 3040
rect 22002 3000 22008 3012
rect 22060 3000 22066 3052
rect 23382 3000 23388 3052
rect 23440 3000 23446 3052
rect 24578 3040 24584 3052
rect 24539 3012 24584 3040
rect 24578 3000 24584 3012
rect 24636 3000 24642 3052
rect 26234 3000 26240 3052
rect 26292 3040 26298 3052
rect 26605 3043 26663 3049
rect 26605 3040 26617 3043
rect 26292 3012 26617 3040
rect 26292 3000 26298 3012
rect 26605 3009 26617 3012
rect 26651 3009 26663 3043
rect 27246 3040 27252 3052
rect 26605 3003 26663 3009
rect 26712 3012 27252 3040
rect 17402 2972 17408 2984
rect 16224 2944 17408 2972
rect 15933 2935 15991 2941
rect 17402 2932 17408 2944
rect 17460 2932 17466 2984
rect 17862 2932 17868 2984
rect 17920 2972 17926 2984
rect 19978 2972 19984 2984
rect 17920 2944 19984 2972
rect 17920 2932 17926 2944
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 21266 2932 21272 2984
rect 21324 2972 21330 2984
rect 22281 2975 22339 2981
rect 22281 2972 22293 2975
rect 21324 2944 22293 2972
rect 21324 2932 21330 2944
rect 22281 2941 22293 2944
rect 22327 2972 22339 2975
rect 23658 2972 23664 2984
rect 22327 2944 23664 2972
rect 22327 2941 22339 2944
rect 22281 2935 22339 2941
rect 23658 2932 23664 2944
rect 23716 2932 23722 2984
rect 25222 2932 25228 2984
rect 25280 2972 25286 2984
rect 26712 2972 26740 3012
rect 27246 3000 27252 3012
rect 27304 3000 27310 3052
rect 27433 3043 27491 3049
rect 27433 3009 27445 3043
rect 27479 3040 27491 3043
rect 27982 3040 27988 3052
rect 27479 3012 27988 3040
rect 27479 3009 27491 3012
rect 27433 3003 27491 3009
rect 27982 3000 27988 3012
rect 28040 3000 28046 3052
rect 29932 3049 29960 3080
rect 31478 3068 31484 3080
rect 31536 3068 31542 3120
rect 31726 3108 31754 3148
rect 32214 3136 32220 3188
rect 32272 3176 32278 3188
rect 36078 3176 36084 3188
rect 32272 3148 36084 3176
rect 32272 3136 32278 3148
rect 36078 3136 36084 3148
rect 36136 3136 36142 3188
rect 37550 3136 37556 3188
rect 37608 3176 37614 3188
rect 38197 3179 38255 3185
rect 38197 3176 38209 3179
rect 37608 3148 38209 3176
rect 37608 3136 37614 3148
rect 38197 3145 38209 3148
rect 38243 3145 38255 3179
rect 38197 3139 38255 3145
rect 32585 3111 32643 3117
rect 32585 3108 32597 3111
rect 31726 3080 32597 3108
rect 32585 3077 32597 3080
rect 32631 3108 32643 3111
rect 32674 3108 32680 3120
rect 32631 3080 32680 3108
rect 32631 3077 32643 3080
rect 32585 3071 32643 3077
rect 32674 3068 32680 3080
rect 32732 3068 32738 3120
rect 37274 3108 37280 3120
rect 33810 3080 37280 3108
rect 37274 3068 37280 3080
rect 37332 3068 37338 3120
rect 37461 3111 37519 3117
rect 37461 3077 37473 3111
rect 37507 3108 37519 3111
rect 37734 3108 37740 3120
rect 37507 3080 37740 3108
rect 37507 3077 37519 3080
rect 37461 3071 37519 3077
rect 37734 3068 37740 3080
rect 37792 3068 37798 3120
rect 29917 3043 29975 3049
rect 29917 3009 29929 3043
rect 29963 3009 29975 3043
rect 29917 3003 29975 3009
rect 30653 3043 30711 3049
rect 30653 3009 30665 3043
rect 30699 3040 30711 3043
rect 31754 3040 31760 3052
rect 30699 3012 31432 3040
rect 31715 3012 31760 3040
rect 30699 3009 30711 3012
rect 30653 3003 30711 3009
rect 25280 2944 26740 2972
rect 25280 2932 25286 2944
rect 26786 2932 26792 2984
rect 26844 2972 26850 2984
rect 31294 2972 31300 2984
rect 26844 2944 31300 2972
rect 26844 2932 26850 2944
rect 31294 2932 31300 2944
rect 31352 2932 31358 2984
rect 19242 2904 19248 2916
rect 19203 2876 19248 2904
rect 19242 2864 19248 2876
rect 19300 2864 19306 2916
rect 23566 2864 23572 2916
rect 23624 2904 23630 2916
rect 23753 2907 23811 2913
rect 23753 2904 23765 2907
rect 23624 2876 23765 2904
rect 23624 2864 23630 2876
rect 23753 2873 23765 2876
rect 23799 2873 23811 2907
rect 31404 2904 31432 3012
rect 31754 3000 31760 3012
rect 31812 3000 31818 3052
rect 34606 3000 34612 3052
rect 34664 3040 34670 3052
rect 34701 3043 34759 3049
rect 34701 3040 34713 3043
rect 34664 3012 34713 3040
rect 34664 3000 34670 3012
rect 34701 3009 34713 3012
rect 34747 3040 34759 3043
rect 35345 3043 35403 3049
rect 35345 3040 35357 3043
rect 34747 3012 35357 3040
rect 34747 3009 34759 3012
rect 34701 3003 34759 3009
rect 35345 3009 35357 3012
rect 35391 3040 35403 3043
rect 35802 3040 35808 3052
rect 35391 3012 35808 3040
rect 35391 3009 35403 3012
rect 35345 3003 35403 3009
rect 35802 3000 35808 3012
rect 35860 3000 35866 3052
rect 35989 3043 36047 3049
rect 35989 3009 36001 3043
rect 36035 3040 36047 3043
rect 36078 3040 36084 3052
rect 36035 3012 36084 3040
rect 36035 3009 36047 3012
rect 35989 3003 36047 3009
rect 36078 3000 36084 3012
rect 36136 3000 36142 3052
rect 36449 3043 36507 3049
rect 36449 3040 36461 3043
rect 36188 3012 36461 3040
rect 31478 2932 31484 2984
rect 31536 2972 31542 2984
rect 32309 2975 32367 2981
rect 32309 2972 32321 2975
rect 31536 2944 32321 2972
rect 31536 2932 31542 2944
rect 32309 2941 32321 2944
rect 32355 2941 32367 2975
rect 32309 2935 32367 2941
rect 32416 2944 35848 2972
rect 31573 2907 31631 2913
rect 31573 2904 31585 2907
rect 31404 2876 31585 2904
rect 23753 2867 23811 2873
rect 31573 2873 31585 2876
rect 31619 2873 31631 2907
rect 31573 2867 31631 2873
rect 31754 2864 31760 2916
rect 31812 2904 31818 2916
rect 32416 2904 32444 2944
rect 34330 2904 34336 2916
rect 31812 2876 32444 2904
rect 33612 2876 34336 2904
rect 31812 2864 31818 2876
rect 1302 2796 1308 2848
rect 1360 2836 1366 2848
rect 1673 2839 1731 2845
rect 1673 2836 1685 2839
rect 1360 2808 1685 2836
rect 1360 2796 1366 2808
rect 1673 2805 1685 2808
rect 1719 2805 1731 2839
rect 1673 2799 1731 2805
rect 2409 2839 2467 2845
rect 2409 2805 2421 2839
rect 2455 2836 2467 2839
rect 2774 2836 2780 2848
rect 2455 2808 2780 2836
rect 2455 2805 2467 2808
rect 2409 2799 2467 2805
rect 2774 2796 2780 2808
rect 2832 2796 2838 2848
rect 3050 2836 3056 2848
rect 3011 2808 3056 2836
rect 3050 2796 3056 2808
rect 3108 2796 3114 2848
rect 9674 2836 9680 2848
rect 9635 2808 9680 2836
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 11882 2836 11888 2848
rect 11843 2808 11888 2836
rect 11882 2796 11888 2808
rect 11940 2796 11946 2848
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 21358 2836 21364 2848
rect 12492 2808 21364 2836
rect 12492 2796 12498 2808
rect 21358 2796 21364 2808
rect 21416 2796 21422 2848
rect 21542 2796 21548 2848
rect 21600 2836 21606 2848
rect 30190 2836 30196 2848
rect 21600 2808 30196 2836
rect 21600 2796 21606 2808
rect 30190 2796 30196 2808
rect 30248 2796 30254 2848
rect 30282 2796 30288 2848
rect 30340 2836 30346 2848
rect 30469 2839 30527 2845
rect 30469 2836 30481 2839
rect 30340 2808 30481 2836
rect 30340 2796 30346 2808
rect 30469 2805 30481 2808
rect 30515 2805 30527 2839
rect 30469 2799 30527 2805
rect 30558 2796 30564 2848
rect 30616 2836 30622 2848
rect 33612 2836 33640 2876
rect 34330 2864 34336 2876
rect 34388 2864 34394 2916
rect 34422 2864 34428 2916
rect 34480 2904 34486 2916
rect 35820 2913 35848 2944
rect 35805 2907 35863 2913
rect 34480 2876 35756 2904
rect 34480 2864 34486 2876
rect 30616 2808 33640 2836
rect 34057 2839 34115 2845
rect 30616 2796 30622 2808
rect 34057 2805 34069 2839
rect 34103 2836 34115 2839
rect 34238 2836 34244 2848
rect 34103 2808 34244 2836
rect 34103 2805 34115 2808
rect 34057 2799 34115 2805
rect 34238 2796 34244 2808
rect 34296 2796 34302 2848
rect 34514 2796 34520 2848
rect 34572 2836 34578 2848
rect 34609 2839 34667 2845
rect 34609 2836 34621 2839
rect 34572 2808 34621 2836
rect 34572 2796 34578 2808
rect 34609 2805 34621 2808
rect 34655 2805 34667 2839
rect 34609 2799 34667 2805
rect 34698 2796 34704 2848
rect 34756 2836 34762 2848
rect 35253 2839 35311 2845
rect 35253 2836 35265 2839
rect 34756 2808 35265 2836
rect 34756 2796 34762 2808
rect 35253 2805 35265 2808
rect 35299 2805 35311 2839
rect 35728 2836 35756 2876
rect 35805 2873 35817 2907
rect 35851 2873 35863 2907
rect 35805 2867 35863 2873
rect 36188 2836 36216 3012
rect 36449 3009 36461 3012
rect 36495 3009 36507 3043
rect 36449 3003 36507 3009
rect 37366 3000 37372 3052
rect 37424 3040 37430 3052
rect 37645 3043 37703 3049
rect 37645 3040 37657 3043
rect 37424 3012 37657 3040
rect 37424 3000 37430 3012
rect 37645 3009 37657 3012
rect 37691 3009 37703 3043
rect 37645 3003 37703 3009
rect 36630 2836 36636 2848
rect 35728 2808 36216 2836
rect 36591 2808 36636 2836
rect 35253 2799 35311 2805
rect 36630 2796 36636 2808
rect 36688 2796 36694 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 10042 2632 10048 2644
rect 10003 2604 10048 2632
rect 10042 2592 10048 2604
rect 10100 2592 10106 2644
rect 11149 2635 11207 2641
rect 11149 2601 11161 2635
rect 11195 2632 11207 2635
rect 12894 2632 12900 2644
rect 11195 2604 12900 2632
rect 11195 2601 11207 2604
rect 11149 2595 11207 2601
rect 12894 2592 12900 2604
rect 12952 2592 12958 2644
rect 16758 2592 16764 2644
rect 16816 2632 16822 2644
rect 19058 2632 19064 2644
rect 16816 2604 19064 2632
rect 16816 2592 16822 2604
rect 19058 2592 19064 2604
rect 19116 2592 19122 2644
rect 19705 2635 19763 2641
rect 19705 2601 19717 2635
rect 19751 2632 19763 2635
rect 20070 2632 20076 2644
rect 19751 2604 20076 2632
rect 19751 2601 19763 2604
rect 19705 2595 19763 2601
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 20990 2592 20996 2644
rect 21048 2632 21054 2644
rect 22005 2635 22063 2641
rect 22005 2632 22017 2635
rect 21048 2604 22017 2632
rect 21048 2592 21054 2604
rect 22005 2601 22017 2604
rect 22051 2601 22063 2635
rect 22005 2595 22063 2601
rect 23658 2592 23664 2644
rect 23716 2632 23722 2644
rect 24581 2635 24639 2641
rect 24581 2632 24593 2635
rect 23716 2604 24593 2632
rect 23716 2592 23722 2604
rect 24581 2601 24593 2604
rect 24627 2601 24639 2635
rect 24581 2595 24639 2601
rect 29181 2635 29239 2641
rect 29181 2601 29193 2635
rect 29227 2632 29239 2635
rect 30374 2632 30380 2644
rect 29227 2604 30380 2632
rect 29227 2601 29239 2604
rect 29181 2595 29239 2601
rect 30374 2592 30380 2604
rect 30432 2592 30438 2644
rect 31110 2592 31116 2644
rect 31168 2632 31174 2644
rect 31481 2635 31539 2641
rect 31481 2632 31493 2635
rect 31168 2604 31493 2632
rect 31168 2592 31174 2604
rect 31481 2601 31493 2604
rect 31527 2601 31539 2635
rect 34698 2632 34704 2644
rect 31481 2595 31539 2601
rect 32140 2604 34704 2632
rect 9401 2567 9459 2573
rect 9401 2533 9413 2567
rect 9447 2564 9459 2567
rect 10594 2564 10600 2576
rect 9447 2536 10600 2564
rect 9447 2533 9459 2536
rect 9401 2527 9459 2533
rect 10594 2524 10600 2536
rect 10652 2524 10658 2576
rect 13354 2524 13360 2576
rect 13412 2564 13418 2576
rect 13449 2567 13507 2573
rect 13449 2564 13461 2567
rect 13412 2536 13461 2564
rect 13412 2524 13418 2536
rect 13449 2533 13461 2536
rect 13495 2533 13507 2567
rect 13449 2527 13507 2533
rect 18693 2567 18751 2573
rect 18693 2533 18705 2567
rect 18739 2564 18751 2567
rect 19978 2564 19984 2576
rect 18739 2536 19984 2564
rect 18739 2533 18751 2536
rect 18693 2527 18751 2533
rect 19978 2524 19984 2536
rect 20036 2524 20042 2576
rect 2133 2499 2191 2505
rect 2133 2465 2145 2499
rect 2179 2496 2191 2499
rect 2498 2496 2504 2508
rect 2179 2468 2504 2496
rect 2179 2465 2191 2468
rect 2133 2459 2191 2465
rect 2498 2456 2504 2468
rect 2556 2456 2562 2508
rect 4062 2496 4068 2508
rect 4023 2468 4068 2496
rect 4062 2456 4068 2468
rect 4120 2456 4126 2508
rect 9766 2496 9772 2508
rect 4908 2468 9772 2496
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 2409 2431 2467 2437
rect 2409 2428 2421 2431
rect 72 2400 2421 2428
rect 72 2388 78 2400
rect 2409 2397 2421 2400
rect 2455 2428 2467 2431
rect 3050 2428 3056 2440
rect 2455 2400 3056 2428
rect 2455 2397 2467 2400
rect 2409 2391 2467 2397
rect 3050 2388 3056 2400
rect 3108 2388 3114 2440
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2428 3479 2431
rect 4080 2428 4108 2456
rect 4908 2437 4936 2468
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 17034 2496 17040 2508
rect 15488 2468 17040 2496
rect 3467 2400 4108 2428
rect 4893 2431 4951 2437
rect 3467 2397 3479 2400
rect 3421 2391 3479 2397
rect 4893 2397 4905 2431
rect 4939 2397 4951 2431
rect 6546 2428 6552 2440
rect 6507 2400 6552 2428
rect 4893 2391 4951 2397
rect 6546 2388 6552 2400
rect 6604 2388 6610 2440
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 9732 2400 9873 2428
rect 9732 2388 9738 2400
rect 9861 2397 9873 2400
rect 9907 2397 9919 2431
rect 9861 2391 9919 2397
rect 11054 2388 11060 2440
rect 11112 2428 11118 2440
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 11112 2400 11989 2428
rect 11112 2388 11118 2400
rect 11977 2397 11989 2400
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 13998 2388 14004 2440
rect 14056 2428 14062 2440
rect 15488 2437 15516 2468
rect 17034 2456 17040 2468
rect 17092 2456 17098 2508
rect 17586 2496 17592 2508
rect 17547 2468 17592 2496
rect 17586 2456 17592 2468
rect 17644 2456 17650 2508
rect 21453 2499 21511 2505
rect 21453 2465 21465 2499
rect 21499 2496 21511 2499
rect 22002 2496 22008 2508
rect 21499 2468 22008 2496
rect 21499 2465 21511 2468
rect 21453 2459 21511 2465
rect 22002 2456 22008 2468
rect 22060 2496 22066 2508
rect 23753 2499 23811 2505
rect 23753 2496 23765 2499
rect 22060 2468 23765 2496
rect 22060 2456 22066 2468
rect 23753 2465 23765 2468
rect 23799 2496 23811 2499
rect 24578 2496 24584 2508
rect 23799 2468 24584 2496
rect 23799 2465 23811 2468
rect 23753 2459 23811 2465
rect 24578 2456 24584 2468
rect 24636 2456 24642 2508
rect 25958 2456 25964 2508
rect 26016 2496 26022 2508
rect 26053 2499 26111 2505
rect 26053 2496 26065 2499
rect 26016 2468 26065 2496
rect 26016 2456 26022 2468
rect 26053 2465 26065 2468
rect 26099 2465 26111 2499
rect 29730 2496 29736 2508
rect 29691 2468 29736 2496
rect 26053 2459 26111 2465
rect 29730 2456 29736 2468
rect 29788 2456 29794 2508
rect 30009 2499 30067 2505
rect 30009 2465 30021 2499
rect 30055 2496 30067 2499
rect 31386 2496 31392 2508
rect 30055 2468 31392 2496
rect 30055 2465 30067 2468
rect 30009 2459 30067 2465
rect 31386 2456 31392 2468
rect 31444 2456 31450 2508
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 14056 2400 14289 2428
rect 14056 2388 14062 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 15473 2431 15531 2437
rect 15473 2397 15485 2431
rect 15519 2397 15531 2431
rect 15473 2391 15531 2397
rect 16301 2431 16359 2437
rect 16301 2397 16313 2431
rect 16347 2428 16359 2431
rect 16850 2428 16856 2440
rect 16347 2400 16856 2428
rect 16347 2397 16359 2400
rect 16301 2391 16359 2397
rect 16850 2388 16856 2400
rect 16908 2388 16914 2440
rect 17402 2428 17408 2440
rect 17363 2400 17408 2428
rect 17402 2388 17408 2400
rect 17460 2388 17466 2440
rect 18874 2428 18880 2440
rect 18835 2400 18880 2428
rect 18874 2388 18880 2400
rect 18932 2388 18938 2440
rect 26329 2431 26387 2437
rect 26329 2397 26341 2431
rect 26375 2428 26387 2431
rect 27062 2428 27068 2440
rect 26375 2400 27068 2428
rect 26375 2397 26387 2400
rect 26329 2391 26387 2397
rect 27062 2388 27068 2400
rect 27120 2428 27126 2440
rect 27430 2428 27436 2440
rect 27120 2400 27436 2428
rect 27120 2388 27126 2400
rect 27430 2388 27436 2400
rect 27488 2388 27494 2440
rect 9217 2363 9275 2369
rect 9217 2329 9229 2363
rect 9263 2329 9275 2363
rect 9217 2323 9275 2329
rect 10597 2363 10655 2369
rect 10597 2329 10609 2363
rect 10643 2360 10655 2363
rect 13538 2360 13544 2372
rect 10643 2332 13544 2360
rect 10643 2329 10655 2332
rect 10597 2323 10655 2329
rect 3234 2292 3240 2304
rect 3195 2264 3240 2292
rect 3234 2252 3240 2264
rect 3292 2252 3298 2304
rect 4522 2252 4528 2304
rect 4580 2292 4586 2304
rect 4709 2295 4767 2301
rect 4709 2292 4721 2295
rect 4580 2264 4721 2292
rect 4580 2252 4586 2264
rect 4709 2261 4721 2264
rect 4755 2261 4767 2295
rect 4709 2255 4767 2261
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 6512 2264 6745 2292
rect 6512 2252 6518 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 8481 2295 8539 2301
rect 8481 2292 8493 2295
rect 8444 2264 8493 2292
rect 8444 2252 8450 2264
rect 8481 2261 8493 2264
rect 8527 2292 8539 2295
rect 9232 2292 9260 2323
rect 13538 2320 13544 2332
rect 13596 2360 13602 2372
rect 13633 2363 13691 2369
rect 13633 2360 13645 2363
rect 13596 2332 13645 2360
rect 13596 2320 13602 2332
rect 13633 2329 13645 2332
rect 13679 2329 13691 2363
rect 14550 2360 14556 2372
rect 14511 2332 14556 2360
rect 13633 2323 13691 2329
rect 14550 2320 14556 2332
rect 14608 2320 14614 2372
rect 20622 2320 20628 2372
rect 20680 2320 20686 2372
rect 21177 2363 21235 2369
rect 21177 2329 21189 2363
rect 21223 2329 21235 2363
rect 23046 2332 23336 2360
rect 21177 2323 21235 2329
rect 8527 2264 9260 2292
rect 8527 2261 8539 2264
rect 8481 2255 8539 2261
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11793 2295 11851 2301
rect 11793 2292 11805 2295
rect 11664 2264 11805 2292
rect 11664 2252 11670 2264
rect 11793 2261 11805 2264
rect 11839 2261 11851 2295
rect 11793 2255 11851 2261
rect 14826 2252 14832 2304
rect 14884 2292 14890 2304
rect 15289 2295 15347 2301
rect 15289 2292 15301 2295
rect 14884 2264 15301 2292
rect 14884 2252 14890 2264
rect 15289 2261 15301 2264
rect 15335 2261 15347 2295
rect 15289 2255 15347 2261
rect 16117 2295 16175 2301
rect 16117 2261 16129 2295
rect 16163 2292 16175 2295
rect 16758 2292 16764 2304
rect 16163 2264 16764 2292
rect 16163 2261 16175 2264
rect 16117 2255 16175 2261
rect 16758 2252 16764 2264
rect 16816 2252 16822 2304
rect 16945 2295 17003 2301
rect 16945 2261 16957 2295
rect 16991 2292 17003 2295
rect 18966 2292 18972 2304
rect 16991 2264 18972 2292
rect 16991 2261 17003 2264
rect 16945 2255 17003 2261
rect 18966 2252 18972 2264
rect 19024 2292 19030 2304
rect 21192 2292 21220 2323
rect 19024 2264 21220 2292
rect 23308 2292 23336 2332
rect 23382 2320 23388 2372
rect 23440 2360 23446 2372
rect 23477 2363 23535 2369
rect 23477 2360 23489 2363
rect 23440 2332 23489 2360
rect 23440 2320 23446 2332
rect 23477 2329 23489 2332
rect 23523 2329 23535 2363
rect 23477 2323 23535 2329
rect 23566 2320 23572 2372
rect 23624 2360 23630 2372
rect 23624 2332 24886 2360
rect 23624 2320 23630 2332
rect 26786 2320 26792 2372
rect 26844 2360 26850 2372
rect 27706 2360 27712 2372
rect 26844 2332 27108 2360
rect 27667 2332 27712 2360
rect 26844 2320 26850 2332
rect 26970 2292 26976 2304
rect 23308 2264 26976 2292
rect 19024 2252 19030 2264
rect 26970 2252 26976 2264
rect 27028 2252 27034 2304
rect 27080 2292 27108 2332
rect 27706 2320 27712 2332
rect 27764 2320 27770 2372
rect 29914 2360 29920 2372
rect 28934 2332 29920 2360
rect 29914 2320 29920 2332
rect 29972 2320 29978 2372
rect 31294 2360 31300 2372
rect 31234 2332 31300 2360
rect 31294 2320 31300 2332
rect 31352 2320 31358 2372
rect 32140 2292 32168 2604
rect 34698 2592 34704 2604
rect 34756 2592 34762 2644
rect 32309 2567 32367 2573
rect 32309 2533 32321 2567
rect 32355 2564 32367 2567
rect 32582 2564 32588 2576
rect 32355 2536 32588 2564
rect 32355 2533 32367 2536
rect 32309 2527 32367 2533
rect 32582 2524 32588 2536
rect 32640 2524 32646 2576
rect 33778 2496 33784 2508
rect 33739 2468 33784 2496
rect 33778 2456 33784 2468
rect 33836 2456 33842 2508
rect 34054 2496 34060 2508
rect 34015 2468 34060 2496
rect 34054 2456 34060 2468
rect 34112 2456 34118 2508
rect 35802 2496 35808 2508
rect 35176 2468 35808 2496
rect 35176 2437 35204 2468
rect 35802 2456 35808 2468
rect 35860 2456 35866 2508
rect 37461 2499 37519 2505
rect 37461 2465 37473 2499
rect 37507 2496 37519 2499
rect 37642 2496 37648 2508
rect 37507 2468 37648 2496
rect 37507 2465 37519 2468
rect 37461 2459 37519 2465
rect 37642 2456 37648 2468
rect 37700 2456 37706 2508
rect 37737 2499 37795 2505
rect 37737 2465 37749 2499
rect 37783 2496 37795 2499
rect 38378 2496 38384 2508
rect 37783 2468 38384 2496
rect 37783 2465 37795 2468
rect 37737 2459 37795 2465
rect 38378 2456 38384 2468
rect 38436 2456 38442 2508
rect 35161 2431 35219 2437
rect 35161 2397 35173 2431
rect 35207 2397 35219 2431
rect 35161 2391 35219 2397
rect 35621 2431 35679 2437
rect 35621 2397 35633 2431
rect 35667 2397 35679 2431
rect 36630 2428 36636 2440
rect 36591 2400 36636 2428
rect 35621 2391 35679 2397
rect 33318 2320 33324 2372
rect 33376 2320 33382 2372
rect 33686 2320 33692 2372
rect 33744 2360 33750 2372
rect 35636 2360 35664 2391
rect 36630 2388 36636 2400
rect 36688 2388 36694 2440
rect 37660 2428 37688 2456
rect 39298 2428 39304 2440
rect 37660 2400 39304 2428
rect 39298 2388 39304 2400
rect 39356 2388 39362 2440
rect 33744 2332 35664 2360
rect 33744 2320 33750 2332
rect 27080 2264 32168 2292
rect 34146 2252 34152 2304
rect 34204 2292 34210 2304
rect 34977 2295 35035 2301
rect 34977 2292 34989 2295
rect 34204 2264 34989 2292
rect 34204 2252 34210 2264
rect 34977 2261 34989 2264
rect 35023 2261 35035 2295
rect 34977 2255 35035 2261
rect 35434 2252 35440 2304
rect 35492 2292 35498 2304
rect 35805 2295 35863 2301
rect 35805 2292 35817 2295
rect 35492 2264 35817 2292
rect 35492 2252 35498 2264
rect 35805 2261 35817 2264
rect 35851 2261 35863 2295
rect 35805 2255 35863 2261
rect 36817 2295 36875 2301
rect 36817 2261 36829 2295
rect 36863 2292 36875 2295
rect 37182 2292 37188 2304
rect 36863 2264 37188 2292
rect 36863 2261 36875 2264
rect 36817 2255 36875 2261
rect 37182 2252 37188 2264
rect 37240 2252 37246 2304
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 21818 2048 21824 2100
rect 21876 2088 21882 2100
rect 26786 2088 26792 2100
rect 21876 2060 26792 2088
rect 21876 2048 21882 2060
rect 26786 2048 26792 2060
rect 26844 2048 26850 2100
rect 26878 2048 26884 2100
rect 26936 2088 26942 2100
rect 35618 2088 35624 2100
rect 26936 2060 35624 2088
rect 26936 2048 26942 2060
rect 35618 2048 35624 2060
rect 35676 2048 35682 2100
rect 14550 1980 14556 2032
rect 14608 2020 14614 2032
rect 32398 2020 32404 2032
rect 14608 1992 32404 2020
rect 14608 1980 14614 1992
rect 32398 1980 32404 1992
rect 32456 1980 32462 2032
rect 21634 1912 21640 1964
rect 21692 1952 21698 1964
rect 26878 1952 26884 1964
rect 21692 1924 26884 1952
rect 21692 1912 21698 1924
rect 26878 1912 26884 1924
rect 26936 1912 26942 1964
rect 26970 1912 26976 1964
rect 27028 1952 27034 1964
rect 35342 1952 35348 1964
rect 27028 1924 35348 1952
rect 27028 1912 27034 1924
rect 35342 1912 35348 1924
rect 35400 1912 35406 1964
rect 11882 1844 11888 1896
rect 11940 1884 11946 1896
rect 23566 1884 23572 1896
rect 11940 1856 23572 1884
rect 11940 1844 11946 1856
rect 23566 1844 23572 1856
rect 23624 1844 23630 1896
rect 35894 1884 35900 1896
rect 24136 1856 35900 1884
rect 19058 1776 19064 1828
rect 19116 1816 19122 1828
rect 24136 1816 24164 1856
rect 35894 1844 35900 1856
rect 35952 1844 35958 1896
rect 19116 1788 24164 1816
rect 19116 1776 19122 1788
rect 29914 1776 29920 1828
rect 29972 1816 29978 1828
rect 36998 1816 37004 1828
rect 29972 1788 37004 1816
rect 29972 1776 29978 1788
rect 36998 1776 37004 1788
rect 37056 1776 37062 1828
rect 27706 1708 27712 1760
rect 27764 1748 27770 1760
rect 33502 1748 33508 1760
rect 27764 1720 33508 1748
rect 27764 1708 27770 1720
rect 33502 1708 33508 1720
rect 33560 1748 33566 1760
rect 34238 1748 34244 1760
rect 33560 1720 34244 1748
rect 33560 1708 33566 1720
rect 34238 1708 34244 1720
rect 34296 1708 34302 1760
rect 32398 1640 32404 1692
rect 32456 1680 32462 1692
rect 34606 1680 34612 1692
rect 32456 1652 34612 1680
rect 32456 1640 32462 1652
rect 34606 1640 34612 1652
rect 34664 1640 34670 1692
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 36820 37451 36872 37460
rect 36820 37417 36829 37451
rect 36829 37417 36863 37451
rect 36863 37417 36872 37451
rect 36820 37408 36872 37417
rect 17316 37340 17368 37392
rect 1400 37204 1452 37256
rect 6552 37272 6604 37324
rect 11520 37272 11572 37324
rect 12900 37272 12952 37324
rect 2504 37204 2556 37256
rect 6460 37204 6512 37256
rect 8116 37247 8168 37256
rect 8116 37213 8125 37247
rect 8125 37213 8159 37247
rect 8159 37213 8168 37247
rect 8116 37204 8168 37213
rect 9680 37204 9732 37256
rect 15200 37247 15252 37256
rect 10692 37136 10744 37188
rect 15200 37213 15209 37247
rect 15209 37213 15243 37247
rect 15243 37213 15252 37247
rect 15200 37204 15252 37213
rect 17132 37247 17184 37256
rect 17132 37213 17141 37247
rect 17141 37213 17175 37247
rect 17175 37213 17184 37247
rect 17132 37204 17184 37213
rect 18420 37247 18472 37256
rect 18420 37213 18429 37247
rect 18429 37213 18463 37247
rect 18463 37213 18472 37247
rect 18420 37204 18472 37213
rect 20352 37247 20404 37256
rect 20352 37213 20361 37247
rect 20361 37213 20395 37247
rect 20395 37213 20404 37247
rect 21916 37272 21968 37324
rect 22284 37247 22336 37256
rect 20352 37204 20404 37213
rect 22284 37213 22293 37247
rect 22293 37213 22327 37247
rect 22327 37213 22336 37247
rect 22284 37204 22336 37213
rect 23204 37204 23256 37256
rect 25136 37204 25188 37256
rect 27160 37247 27212 37256
rect 27160 37213 27169 37247
rect 27169 37213 27203 37247
rect 27203 37213 27212 37247
rect 27160 37204 27212 37213
rect 27344 37204 27396 37256
rect 30380 37247 30432 37256
rect 30380 37213 30389 37247
rect 30389 37213 30423 37247
rect 30423 37213 30432 37247
rect 30380 37204 30432 37213
rect 30656 37204 30708 37256
rect 33600 37247 33652 37256
rect 33600 37213 33609 37247
rect 33609 37213 33643 37247
rect 33643 37213 33652 37247
rect 33600 37204 33652 37213
rect 34796 37204 34848 37256
rect 15568 37136 15620 37188
rect 26332 37136 26384 37188
rect 36452 37136 36504 37188
rect 1768 37111 1820 37120
rect 1768 37077 1777 37111
rect 1777 37077 1811 37111
rect 1811 37077 1820 37111
rect 1768 37068 1820 37077
rect 2780 37068 2832 37120
rect 4620 37068 4672 37120
rect 5448 37111 5500 37120
rect 5448 37077 5457 37111
rect 5457 37077 5491 37111
rect 5491 37077 5500 37111
rect 5448 37068 5500 37077
rect 7748 37068 7800 37120
rect 14832 37068 14884 37120
rect 16764 37068 16816 37120
rect 18052 37068 18104 37120
rect 19984 37068 20036 37120
rect 25412 37111 25464 37120
rect 25412 37077 25421 37111
rect 25421 37077 25455 37111
rect 25455 37077 25464 37111
rect 25412 37068 25464 37077
rect 27068 37068 27120 37120
rect 28356 37068 28408 37120
rect 30288 37068 30340 37120
rect 32220 37068 32272 37120
rect 33508 37068 33560 37120
rect 34796 37068 34848 37120
rect 35440 37068 35492 37120
rect 36268 37068 36320 37120
rect 37372 37068 37424 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 2872 36864 2924 36916
rect 1676 36839 1728 36848
rect 1676 36805 1685 36839
rect 1685 36805 1719 36839
rect 1719 36805 1728 36839
rect 1676 36796 1728 36805
rect 8116 36864 8168 36916
rect 23204 36907 23256 36916
rect 23204 36873 23213 36907
rect 23213 36873 23247 36907
rect 23247 36873 23256 36907
rect 23204 36864 23256 36873
rect 33600 36864 33652 36916
rect 36268 36864 36320 36916
rect 36452 36907 36504 36916
rect 36452 36873 36461 36907
rect 36461 36873 36495 36907
rect 36495 36873 36504 36907
rect 36452 36864 36504 36873
rect 38200 36907 38252 36916
rect 38200 36873 38209 36907
rect 38209 36873 38243 36907
rect 38243 36873 38252 36907
rect 38200 36864 38252 36873
rect 10692 36771 10744 36780
rect 10692 36737 10701 36771
rect 10701 36737 10735 36771
rect 10735 36737 10744 36771
rect 10692 36728 10744 36737
rect 11612 36728 11664 36780
rect 22284 36728 22336 36780
rect 35532 36728 35584 36780
rect 37280 36728 37332 36780
rect 11980 36703 12032 36712
rect 11980 36669 11989 36703
rect 11989 36669 12023 36703
rect 12023 36669 12032 36703
rect 11980 36660 12032 36669
rect 2136 36592 2188 36644
rect 35532 36567 35584 36576
rect 35532 36533 35541 36567
rect 35541 36533 35575 36567
rect 35575 36533 35584 36567
rect 35532 36524 35584 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 11612 36363 11664 36372
rect 11612 36329 11621 36363
rect 11621 36329 11655 36363
rect 11655 36329 11664 36363
rect 11612 36320 11664 36329
rect 38660 36320 38712 36372
rect 1860 36159 1912 36168
rect 1860 36125 1869 36159
rect 1869 36125 1903 36159
rect 1903 36125 1912 36159
rect 1860 36116 1912 36125
rect 37372 36159 37424 36168
rect 37372 36125 37381 36159
rect 37381 36125 37415 36159
rect 37415 36125 37424 36159
rect 37372 36116 37424 36125
rect 1676 36023 1728 36032
rect 1676 35989 1685 36023
rect 1685 35989 1719 36023
rect 1719 35989 1728 36023
rect 1676 35980 1728 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 30380 35776 30432 35828
rect 28540 35640 28592 35692
rect 37372 35572 37424 35624
rect 38292 35615 38344 35624
rect 38292 35581 38301 35615
rect 38301 35581 38335 35615
rect 38335 35581 38344 35615
rect 38292 35572 38344 35581
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 38292 35275 38344 35284
rect 38292 35241 38301 35275
rect 38301 35241 38335 35275
rect 38335 35241 38344 35275
rect 38292 35232 38344 35241
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 1860 34688 1912 34740
rect 2044 34552 2096 34604
rect 13084 34484 13136 34536
rect 1676 34391 1728 34400
rect 1676 34357 1685 34391
rect 1685 34357 1719 34391
rect 1719 34357 1728 34391
rect 1676 34348 1728 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 25688 33464 25740 33516
rect 38200 33371 38252 33380
rect 38200 33337 38209 33371
rect 38209 33337 38243 33371
rect 38243 33337 38252 33371
rect 38200 33328 38252 33337
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 27344 32555 27396 32564
rect 27344 32521 27353 32555
rect 27353 32521 27387 32555
rect 27387 32521 27396 32555
rect 27344 32512 27396 32521
rect 9128 32376 9180 32428
rect 1676 32215 1728 32224
rect 1676 32181 1685 32215
rect 1685 32181 1719 32215
rect 1719 32181 1728 32215
rect 1676 32172 1728 32181
rect 28540 32308 28592 32360
rect 38292 32351 38344 32360
rect 38292 32317 38301 32351
rect 38301 32317 38335 32351
rect 38335 32317 38344 32351
rect 38292 32308 38344 32317
rect 28632 32172 28684 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 38292 32011 38344 32020
rect 38292 31977 38301 32011
rect 38301 31977 38335 32011
rect 38335 31977 38344 32011
rect 38292 31968 38344 31977
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 2504 30923 2556 30932
rect 2504 30889 2513 30923
rect 2513 30889 2547 30923
rect 2547 30889 2556 30923
rect 2504 30880 2556 30889
rect 30656 30880 30708 30932
rect 1952 30676 2004 30728
rect 26976 30676 27028 30728
rect 1676 30651 1728 30660
rect 1676 30617 1685 30651
rect 1685 30617 1719 30651
rect 1719 30617 1728 30651
rect 1676 30608 1728 30617
rect 2228 30608 2280 30660
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 1676 30379 1728 30388
rect 1676 30345 1685 30379
rect 1685 30345 1719 30379
rect 1719 30345 1728 30379
rect 1676 30336 1728 30345
rect 30196 30243 30248 30252
rect 30196 30209 30205 30243
rect 30205 30209 30239 30243
rect 30239 30209 30248 30243
rect 30196 30200 30248 30209
rect 38200 30243 38252 30252
rect 38200 30209 38209 30243
rect 38209 30209 38243 30243
rect 38243 30209 38252 30243
rect 38200 30200 38252 30209
rect 37280 30064 37332 30116
rect 38108 30039 38160 30048
rect 38108 30005 38117 30039
rect 38117 30005 38151 30039
rect 38151 30005 38160 30039
rect 38108 29996 38160 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 5448 29452 5500 29504
rect 23664 29495 23716 29504
rect 23664 29461 23673 29495
rect 23673 29461 23707 29495
rect 23707 29461 23716 29495
rect 23664 29452 23716 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 1584 29112 1636 29164
rect 25596 28976 25648 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 18420 28704 18472 28756
rect 1584 28679 1636 28688
rect 1584 28645 1593 28679
rect 1593 28645 1627 28679
rect 1627 28645 1636 28679
rect 1584 28636 1636 28645
rect 15568 28543 15620 28552
rect 15568 28509 15577 28543
rect 15577 28509 15611 28543
rect 15611 28509 15620 28543
rect 15568 28500 15620 28509
rect 15660 28407 15712 28416
rect 15660 28373 15669 28407
rect 15669 28373 15703 28407
rect 15703 28373 15712 28407
rect 15660 28364 15712 28373
rect 23112 28364 23164 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 17132 28160 17184 28212
rect 25596 28203 25648 28212
rect 25596 28169 25605 28203
rect 25605 28169 25639 28203
rect 25639 28169 25648 28203
rect 25596 28160 25648 28169
rect 26332 28203 26384 28212
rect 26332 28169 26341 28203
rect 26341 28169 26375 28203
rect 26375 28169 26384 28203
rect 26332 28160 26384 28169
rect 15200 28092 15252 28144
rect 18512 28067 18564 28076
rect 18512 28033 18521 28067
rect 18521 28033 18555 28067
rect 18555 28033 18564 28067
rect 18512 28024 18564 28033
rect 22284 28024 22336 28076
rect 28540 28067 28592 28076
rect 28540 28033 28549 28067
rect 28549 28033 28583 28067
rect 28583 28033 28592 28067
rect 28540 28024 28592 28033
rect 38200 28067 38252 28076
rect 38200 28033 38209 28067
rect 38209 28033 38243 28067
rect 38243 28033 38252 28067
rect 38200 28024 38252 28033
rect 24768 27956 24820 28008
rect 24860 27888 24912 27940
rect 37924 27888 37976 27940
rect 22928 27820 22980 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 11980 27412 12032 27464
rect 37372 27412 37424 27464
rect 15568 27276 15620 27328
rect 18512 27276 18564 27328
rect 21456 27276 21508 27328
rect 26424 27276 26476 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 6828 26936 6880 26988
rect 23664 26868 23716 26920
rect 38292 26911 38344 26920
rect 38292 26877 38301 26911
rect 38301 26877 38335 26911
rect 38335 26877 38344 26911
rect 38292 26868 38344 26877
rect 1676 26775 1728 26784
rect 1676 26741 1685 26775
rect 1685 26741 1719 26775
rect 1719 26741 1728 26775
rect 1676 26732 1728 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 38292 26571 38344 26580
rect 38292 26537 38301 26571
rect 38301 26537 38335 26571
rect 38335 26537 38344 26571
rect 38292 26528 38344 26537
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 2044 25440 2096 25492
rect 9128 25483 9180 25492
rect 9128 25449 9137 25483
rect 9137 25449 9171 25483
rect 9171 25449 9180 25483
rect 9128 25440 9180 25449
rect 1584 25279 1636 25288
rect 1584 25245 1593 25279
rect 1593 25245 1627 25279
rect 1627 25245 1636 25279
rect 1584 25236 1636 25245
rect 1952 25236 2004 25288
rect 7840 25143 7892 25152
rect 7840 25109 7849 25143
rect 7849 25109 7883 25143
rect 7883 25109 7892 25143
rect 7840 25100 7892 25109
rect 9772 25143 9824 25152
rect 9772 25109 9781 25143
rect 9781 25109 9815 25143
rect 9815 25109 9824 25143
rect 9772 25100 9824 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 1584 24939 1636 24948
rect 1584 24905 1593 24939
rect 1593 24905 1627 24939
rect 1627 24905 1636 24939
rect 1584 24896 1636 24905
rect 37832 24692 37884 24744
rect 38292 24735 38344 24744
rect 38292 24701 38301 24735
rect 38301 24701 38335 24735
rect 38335 24701 38344 24735
rect 38292 24692 38344 24701
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 38292 24395 38344 24404
rect 38292 24361 38301 24395
rect 38301 24361 38335 24395
rect 38335 24361 38344 24395
rect 38292 24352 38344 24361
rect 20352 24148 20404 24200
rect 27804 24148 27856 24200
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1584 23647 1636 23656
rect 1584 23613 1593 23647
rect 1593 23613 1627 23647
rect 1627 23613 1636 23647
rect 1584 23604 1636 23613
rect 1860 23647 1912 23656
rect 1860 23613 1869 23647
rect 1869 23613 1903 23647
rect 1903 23613 1912 23647
rect 1860 23604 1912 23613
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 23664 23264 23716 23316
rect 1584 23239 1636 23248
rect 1584 23205 1593 23239
rect 1593 23205 1627 23239
rect 1627 23205 1636 23239
rect 1584 23196 1636 23205
rect 23664 23060 23716 23112
rect 22836 22924 22888 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 35992 22584 36044 22636
rect 38200 22491 38252 22500
rect 38200 22457 38209 22491
rect 38209 22457 38243 22491
rect 38243 22457 38252 22491
rect 38200 22448 38252 22457
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 25596 22040 25648 22092
rect 22652 21836 22704 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 6828 21632 6880 21684
rect 25688 21675 25740 21684
rect 25688 21641 25697 21675
rect 25697 21641 25731 21675
rect 25731 21641 25740 21675
rect 25688 21632 25740 21641
rect 35992 21632 36044 21684
rect 1768 21496 1820 21548
rect 1676 21335 1728 21344
rect 1676 21301 1685 21335
rect 1685 21301 1719 21335
rect 1719 21301 1728 21335
rect 1676 21292 1728 21301
rect 13544 21292 13596 21344
rect 21272 21292 21324 21344
rect 30012 21496 30064 21548
rect 38016 21539 38068 21548
rect 38016 21505 38025 21539
rect 38025 21505 38059 21539
rect 38059 21505 38068 21539
rect 38016 21496 38068 21505
rect 38200 21335 38252 21344
rect 38200 21301 38209 21335
rect 38209 21301 38243 21335
rect 38243 21301 38252 21335
rect 38200 21292 38252 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1768 21131 1820 21140
rect 1768 21097 1777 21131
rect 1777 21097 1811 21131
rect 1811 21097 1820 21131
rect 1768 21088 1820 21097
rect 1952 20927 2004 20936
rect 1952 20893 1961 20927
rect 1961 20893 1995 20927
rect 1995 20893 2004 20927
rect 1952 20884 2004 20893
rect 24952 20884 25004 20936
rect 13084 20748 13136 20800
rect 20352 20748 20404 20800
rect 22008 20748 22060 20800
rect 25136 20748 25188 20800
rect 25412 20748 25464 20800
rect 27528 20748 27580 20800
rect 30012 20748 30064 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 2228 20408 2280 20460
rect 22008 20408 22060 20460
rect 23112 20408 23164 20460
rect 24860 20408 24912 20460
rect 24952 20408 25004 20460
rect 26148 20408 26200 20460
rect 22376 20247 22428 20256
rect 22376 20213 22385 20247
rect 22385 20213 22419 20247
rect 22419 20213 22428 20247
rect 22376 20204 22428 20213
rect 26056 20340 26108 20392
rect 38016 20272 38068 20324
rect 24860 20204 24912 20256
rect 25228 20204 25280 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 26056 20043 26108 20052
rect 26056 20009 26065 20043
rect 26065 20009 26099 20043
rect 26099 20009 26108 20043
rect 26056 20000 26108 20009
rect 23112 19932 23164 19984
rect 22376 19864 22428 19916
rect 24768 19932 24820 19984
rect 23756 19839 23808 19848
rect 1676 19771 1728 19780
rect 1676 19737 1685 19771
rect 1685 19737 1719 19771
rect 1719 19737 1728 19771
rect 1676 19728 1728 19737
rect 23756 19805 23765 19839
rect 23765 19805 23799 19839
rect 23799 19805 23808 19839
rect 23756 19796 23808 19805
rect 26148 19839 26200 19848
rect 26148 19805 26157 19839
rect 26157 19805 26191 19839
rect 26191 19805 26200 19839
rect 26148 19796 26200 19805
rect 19432 19660 19484 19712
rect 22192 19703 22244 19712
rect 22192 19669 22201 19703
rect 22201 19669 22235 19703
rect 22235 19669 22244 19703
rect 22192 19660 22244 19669
rect 23112 19703 23164 19712
rect 23112 19669 23121 19703
rect 23121 19669 23155 19703
rect 23155 19669 23164 19703
rect 23112 19660 23164 19669
rect 24032 19660 24084 19712
rect 24676 19660 24728 19712
rect 26608 19728 26660 19780
rect 26332 19660 26384 19712
rect 26700 19703 26752 19712
rect 26700 19669 26709 19703
rect 26709 19669 26743 19703
rect 26743 19669 26752 19703
rect 26700 19660 26752 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 1676 19499 1728 19508
rect 1676 19465 1685 19499
rect 1685 19465 1719 19499
rect 1719 19465 1728 19499
rect 1676 19456 1728 19465
rect 22100 19456 22152 19508
rect 24032 19431 24084 19440
rect 24032 19397 24041 19431
rect 24041 19397 24075 19431
rect 24075 19397 24084 19431
rect 24032 19388 24084 19397
rect 1952 19320 2004 19372
rect 16948 19320 17000 19372
rect 21916 19320 21968 19372
rect 22192 19363 22244 19372
rect 22192 19329 22201 19363
rect 22201 19329 22235 19363
rect 22235 19329 22244 19363
rect 22192 19320 22244 19329
rect 24308 19320 24360 19372
rect 21916 19184 21968 19236
rect 24768 19252 24820 19304
rect 25136 19295 25188 19304
rect 25136 19261 25145 19295
rect 25145 19261 25179 19295
rect 25179 19261 25188 19295
rect 25136 19252 25188 19261
rect 25780 19252 25832 19304
rect 26240 19320 26292 19372
rect 26700 19320 26752 19372
rect 27160 19320 27212 19372
rect 33600 19320 33652 19372
rect 26332 19252 26384 19304
rect 21364 19159 21416 19168
rect 21364 19125 21373 19159
rect 21373 19125 21407 19159
rect 21407 19125 21416 19159
rect 21364 19116 21416 19125
rect 27344 19116 27396 19168
rect 27620 19116 27672 19168
rect 38200 19159 38252 19168
rect 38200 19125 38209 19159
rect 38209 19125 38243 19159
rect 38243 19125 38252 19159
rect 38200 19116 38252 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 19432 18912 19484 18964
rect 1860 18708 1912 18760
rect 22100 18955 22152 18964
rect 22100 18921 22109 18955
rect 22109 18921 22143 18955
rect 22143 18921 22152 18955
rect 22100 18912 22152 18921
rect 26976 18912 27028 18964
rect 24860 18844 24912 18896
rect 21364 18776 21416 18828
rect 22652 18819 22704 18828
rect 22652 18785 22661 18819
rect 22661 18785 22695 18819
rect 22695 18785 22704 18819
rect 22652 18776 22704 18785
rect 23756 18819 23808 18828
rect 23756 18785 23765 18819
rect 23765 18785 23799 18819
rect 23799 18785 23808 18819
rect 23756 18776 23808 18785
rect 25228 18776 25280 18828
rect 26056 18844 26108 18896
rect 30196 18776 30248 18828
rect 18328 18640 18380 18692
rect 27252 18751 27304 18760
rect 22008 18640 22060 18692
rect 22468 18640 22520 18692
rect 22744 18683 22796 18692
rect 22744 18649 22753 18683
rect 22753 18649 22787 18683
rect 22787 18649 22796 18683
rect 23296 18683 23348 18692
rect 22744 18640 22796 18649
rect 23296 18649 23305 18683
rect 23305 18649 23339 18683
rect 23339 18649 23348 18683
rect 23296 18640 23348 18649
rect 17500 18572 17552 18624
rect 20260 18615 20312 18624
rect 20260 18581 20269 18615
rect 20269 18581 20303 18615
rect 20303 18581 20312 18615
rect 20260 18572 20312 18581
rect 21916 18572 21968 18624
rect 24952 18572 25004 18624
rect 25136 18640 25188 18692
rect 27252 18717 27261 18751
rect 27261 18717 27295 18751
rect 27295 18717 27304 18751
rect 27252 18708 27304 18717
rect 27620 18640 27672 18692
rect 26516 18615 26568 18624
rect 26516 18581 26525 18615
rect 26525 18581 26559 18615
rect 26559 18581 26568 18615
rect 26516 18572 26568 18581
rect 26700 18572 26752 18624
rect 29276 18572 29328 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 2136 18368 2188 18420
rect 17500 18343 17552 18352
rect 17500 18309 17509 18343
rect 17509 18309 17543 18343
rect 17543 18309 17552 18343
rect 17500 18300 17552 18309
rect 17592 18343 17644 18352
rect 17592 18309 17601 18343
rect 17601 18309 17635 18343
rect 17635 18309 17644 18343
rect 17592 18300 17644 18309
rect 4068 18232 4120 18284
rect 18144 18207 18196 18216
rect 18144 18173 18153 18207
rect 18153 18173 18187 18207
rect 18187 18173 18196 18207
rect 20168 18232 20220 18284
rect 22652 18300 22704 18352
rect 23388 18343 23440 18352
rect 19892 18207 19944 18216
rect 18144 18164 18196 18173
rect 19892 18173 19901 18207
rect 19901 18173 19935 18207
rect 19935 18173 19944 18207
rect 21548 18232 21600 18284
rect 22652 18207 22704 18216
rect 19892 18164 19944 18173
rect 22652 18173 22661 18207
rect 22661 18173 22695 18207
rect 22695 18173 22704 18207
rect 22652 18164 22704 18173
rect 22836 18164 22888 18216
rect 23388 18309 23397 18343
rect 23397 18309 23431 18343
rect 23431 18309 23440 18343
rect 23388 18300 23440 18309
rect 26700 18232 26752 18284
rect 24032 18164 24084 18216
rect 19984 18096 20036 18148
rect 20168 18096 20220 18148
rect 34428 18096 34480 18148
rect 1676 18071 1728 18080
rect 1676 18037 1685 18071
rect 1685 18037 1719 18071
rect 1719 18037 1728 18071
rect 1676 18028 1728 18037
rect 17868 18028 17920 18080
rect 19892 18028 19944 18080
rect 20904 18028 20956 18080
rect 24492 18071 24544 18080
rect 24492 18037 24501 18071
rect 24501 18037 24535 18071
rect 24535 18037 24544 18071
rect 24492 18028 24544 18037
rect 25964 18071 26016 18080
rect 25964 18037 25973 18071
rect 25973 18037 26007 18071
rect 26007 18037 26016 18071
rect 25964 18028 26016 18037
rect 29000 18071 29052 18080
rect 29000 18037 29009 18071
rect 29009 18037 29043 18071
rect 29043 18037 29052 18071
rect 29000 18028 29052 18037
rect 29460 18071 29512 18080
rect 29460 18037 29469 18071
rect 29469 18037 29503 18071
rect 29503 18037 29512 18071
rect 29460 18028 29512 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 17592 17824 17644 17876
rect 22744 17824 22796 17876
rect 23112 17824 23164 17876
rect 27528 17824 27580 17876
rect 15660 17756 15712 17808
rect 19432 17756 19484 17808
rect 20260 17756 20312 17808
rect 24216 17756 24268 17808
rect 16856 17620 16908 17672
rect 24492 17688 24544 17740
rect 26792 17688 26844 17740
rect 16580 17552 16632 17604
rect 20444 17620 20496 17672
rect 20812 17595 20864 17604
rect 20812 17561 20821 17595
rect 20821 17561 20855 17595
rect 20855 17561 20864 17595
rect 20812 17552 20864 17561
rect 20904 17595 20956 17604
rect 20904 17561 20913 17595
rect 20913 17561 20947 17595
rect 20947 17561 20956 17595
rect 20904 17552 20956 17561
rect 21088 17552 21140 17604
rect 21732 17552 21784 17604
rect 18236 17527 18288 17536
rect 18236 17493 18245 17527
rect 18245 17493 18279 17527
rect 18279 17493 18288 17527
rect 18236 17484 18288 17493
rect 19340 17484 19392 17536
rect 20168 17527 20220 17536
rect 20168 17493 20177 17527
rect 20177 17493 20211 17527
rect 20211 17493 20220 17527
rect 20168 17484 20220 17493
rect 24308 17620 24360 17672
rect 26056 17663 26108 17672
rect 26056 17629 26065 17663
rect 26065 17629 26099 17663
rect 26099 17629 26108 17663
rect 26056 17620 26108 17629
rect 26884 17663 26936 17672
rect 26884 17629 26893 17663
rect 26893 17629 26927 17663
rect 26927 17629 26936 17663
rect 26884 17620 26936 17629
rect 27528 17663 27580 17672
rect 27528 17629 27537 17663
rect 27537 17629 27571 17663
rect 27571 17629 27580 17663
rect 27528 17620 27580 17629
rect 28172 17663 28224 17672
rect 28172 17629 28181 17663
rect 28181 17629 28215 17663
rect 28215 17629 28224 17663
rect 28172 17620 28224 17629
rect 22652 17552 22704 17604
rect 25596 17595 25648 17604
rect 25596 17561 25605 17595
rect 25605 17561 25639 17595
rect 25639 17561 25648 17595
rect 25596 17552 25648 17561
rect 28724 17552 28776 17604
rect 25780 17484 25832 17536
rect 26332 17484 26384 17536
rect 27436 17527 27488 17536
rect 27436 17493 27445 17527
rect 27445 17493 27479 17527
rect 27479 17493 27488 17527
rect 27436 17484 27488 17493
rect 27528 17484 27580 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 13084 17280 13136 17332
rect 21640 17280 21692 17332
rect 21916 17280 21968 17332
rect 23388 17280 23440 17332
rect 25964 17280 26016 17332
rect 1584 17144 1636 17196
rect 11704 17144 11756 17196
rect 16856 17187 16908 17196
rect 16856 17153 16865 17187
rect 16865 17153 16899 17187
rect 16899 17153 16908 17187
rect 16856 17144 16908 17153
rect 22192 17255 22244 17264
rect 22192 17221 22201 17255
rect 22201 17221 22235 17255
rect 22235 17221 22244 17255
rect 22192 17212 22244 17221
rect 24584 17212 24636 17264
rect 30288 17280 30340 17332
rect 8300 17076 8352 17128
rect 17684 17076 17736 17128
rect 20536 17144 20588 17196
rect 20996 17076 21048 17128
rect 21272 17187 21324 17196
rect 21272 17153 21281 17187
rect 21281 17153 21315 17187
rect 21315 17153 21324 17187
rect 21272 17144 21324 17153
rect 26240 17187 26292 17196
rect 21732 17076 21784 17128
rect 21824 17076 21876 17128
rect 26240 17153 26249 17187
rect 26249 17153 26283 17187
rect 26283 17153 26292 17187
rect 26240 17144 26292 17153
rect 26424 17187 26476 17196
rect 26424 17153 26433 17187
rect 26433 17153 26467 17187
rect 26467 17153 26476 17187
rect 26424 17144 26476 17153
rect 26516 17144 26568 17196
rect 26884 17144 26936 17196
rect 29000 17212 29052 17264
rect 16672 17008 16724 17060
rect 17776 17051 17828 17060
rect 17776 17017 17785 17051
rect 17785 17017 17819 17051
rect 17819 17017 17828 17051
rect 17776 17008 17828 17017
rect 24768 17076 24820 17128
rect 24952 17119 25004 17128
rect 24952 17085 24961 17119
rect 24961 17085 24995 17119
rect 24995 17085 25004 17119
rect 24952 17076 25004 17085
rect 25504 17076 25556 17128
rect 27528 17076 27580 17128
rect 28080 17144 28132 17196
rect 28632 17187 28684 17196
rect 28632 17153 28641 17187
rect 28641 17153 28675 17187
rect 28675 17153 28684 17187
rect 28632 17144 28684 17153
rect 28908 17144 28960 17196
rect 28724 17076 28776 17128
rect 30012 17076 30064 17128
rect 38292 17119 38344 17128
rect 38292 17085 38301 17119
rect 38301 17085 38335 17119
rect 38335 17085 38344 17119
rect 38292 17076 38344 17085
rect 17408 16940 17460 16992
rect 18052 16940 18104 16992
rect 19340 16940 19392 16992
rect 20536 16940 20588 16992
rect 20720 16983 20772 16992
rect 20720 16949 20729 16983
rect 20729 16949 20763 16983
rect 20763 16949 20772 16983
rect 20720 16940 20772 16949
rect 22560 16940 22612 16992
rect 28172 17008 28224 17060
rect 29460 17008 29512 17060
rect 23480 16940 23532 16992
rect 24308 16940 24360 16992
rect 24768 16940 24820 16992
rect 24860 16940 24912 16992
rect 26792 16940 26844 16992
rect 27344 16940 27396 16992
rect 27896 16983 27948 16992
rect 27896 16949 27905 16983
rect 27905 16949 27939 16983
rect 27939 16949 27948 16983
rect 27896 16940 27948 16949
rect 27988 16940 28040 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 15660 16736 15712 16788
rect 17684 16779 17736 16788
rect 17684 16745 17693 16779
rect 17693 16745 17727 16779
rect 17727 16745 17736 16779
rect 17684 16736 17736 16745
rect 21548 16779 21600 16788
rect 21548 16745 21557 16779
rect 21557 16745 21591 16779
rect 21591 16745 21600 16779
rect 21548 16736 21600 16745
rect 21640 16736 21692 16788
rect 24768 16736 24820 16788
rect 38292 16779 38344 16788
rect 11704 16668 11756 16720
rect 18236 16668 18288 16720
rect 19340 16668 19392 16720
rect 17776 16600 17828 16652
rect 17224 16464 17276 16516
rect 22284 16668 22336 16720
rect 24124 16668 24176 16720
rect 20996 16600 21048 16652
rect 23572 16643 23624 16652
rect 19984 16507 20036 16516
rect 19984 16473 19993 16507
rect 19993 16473 20027 16507
rect 20027 16473 20036 16507
rect 19984 16464 20036 16473
rect 18788 16439 18840 16448
rect 18788 16405 18797 16439
rect 18797 16405 18831 16439
rect 18831 16405 18840 16439
rect 18788 16396 18840 16405
rect 22192 16464 22244 16516
rect 23572 16609 23581 16643
rect 23581 16609 23615 16643
rect 23615 16609 23624 16643
rect 23572 16600 23624 16609
rect 23756 16600 23808 16652
rect 25964 16600 26016 16652
rect 38292 16745 38301 16779
rect 38301 16745 38335 16779
rect 38335 16745 38344 16779
rect 38292 16736 38344 16745
rect 28908 16668 28960 16720
rect 23664 16532 23716 16584
rect 27988 16575 28040 16584
rect 27988 16541 27997 16575
rect 27997 16541 28031 16575
rect 28031 16541 28040 16575
rect 27988 16532 28040 16541
rect 20812 16396 20864 16448
rect 22928 16396 22980 16448
rect 23756 16396 23808 16448
rect 24400 16396 24452 16448
rect 24860 16464 24912 16516
rect 25780 16507 25832 16516
rect 25780 16473 25789 16507
rect 25789 16473 25823 16507
rect 25823 16473 25832 16507
rect 25780 16464 25832 16473
rect 26700 16507 26752 16516
rect 26700 16473 26709 16507
rect 26709 16473 26743 16507
rect 26743 16473 26752 16507
rect 26700 16464 26752 16473
rect 37924 16464 37976 16516
rect 27252 16396 27304 16448
rect 29184 16396 29236 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 18144 16192 18196 16244
rect 18052 16124 18104 16176
rect 20628 16192 20680 16244
rect 24400 16192 24452 16244
rect 24768 16192 24820 16244
rect 20168 16124 20220 16176
rect 23296 16124 23348 16176
rect 23848 16167 23900 16176
rect 23848 16133 23857 16167
rect 23857 16133 23891 16167
rect 23891 16133 23900 16167
rect 23848 16124 23900 16133
rect 14740 16056 14792 16108
rect 19340 16056 19392 16108
rect 19800 16056 19852 16108
rect 19984 16056 20036 16108
rect 21640 16056 21692 16108
rect 16948 16031 17000 16040
rect 16948 15997 16957 16031
rect 16957 15997 16991 16031
rect 16991 15997 17000 16031
rect 16948 15988 17000 15997
rect 18696 15988 18748 16040
rect 22560 16031 22612 16040
rect 22560 15997 22569 16031
rect 22569 15997 22603 16031
rect 22603 15997 22612 16031
rect 22560 15988 22612 15997
rect 24032 16031 24084 16040
rect 24032 15997 24041 16031
rect 24041 15997 24075 16031
rect 24075 15997 24084 16031
rect 26240 16192 26292 16244
rect 26700 16192 26752 16244
rect 28448 16192 28500 16244
rect 25412 16167 25464 16176
rect 25412 16133 25421 16167
rect 25421 16133 25455 16167
rect 25455 16133 25464 16167
rect 25412 16124 25464 16133
rect 27344 16167 27396 16176
rect 27344 16133 27353 16167
rect 27353 16133 27387 16167
rect 27387 16133 27396 16167
rect 27344 16124 27396 16133
rect 29184 16099 29236 16108
rect 29184 16065 29193 16099
rect 29193 16065 29227 16099
rect 29227 16065 29236 16099
rect 29184 16056 29236 16065
rect 30748 16056 30800 16108
rect 38016 16099 38068 16108
rect 38016 16065 38025 16099
rect 38025 16065 38059 16099
rect 38059 16065 38068 16099
rect 38016 16056 38068 16065
rect 24032 15988 24084 15997
rect 26792 15988 26844 16040
rect 27436 15988 27488 16040
rect 27528 16031 27580 16040
rect 27528 15997 27537 16031
rect 27537 15997 27571 16031
rect 27571 15997 27580 16031
rect 27528 15988 27580 15997
rect 18972 15920 19024 15972
rect 20812 15920 20864 15972
rect 21088 15920 21140 15972
rect 25688 15920 25740 15972
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 2412 15895 2464 15904
rect 2412 15861 2421 15895
rect 2421 15861 2455 15895
rect 2455 15861 2464 15895
rect 2412 15852 2464 15861
rect 16028 15852 16080 15904
rect 17776 15852 17828 15904
rect 20536 15852 20588 15904
rect 20904 15895 20956 15904
rect 20904 15861 20913 15895
rect 20913 15861 20947 15895
rect 20947 15861 20956 15895
rect 20904 15852 20956 15861
rect 25964 15852 26016 15904
rect 28172 15852 28224 15904
rect 28724 15920 28776 15972
rect 28816 15852 28868 15904
rect 29368 15852 29420 15904
rect 38200 15895 38252 15904
rect 38200 15861 38209 15895
rect 38209 15861 38243 15895
rect 38243 15861 38252 15895
rect 38200 15852 38252 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 23848 15648 23900 15700
rect 25412 15648 25464 15700
rect 28816 15648 28868 15700
rect 33600 15691 33652 15700
rect 33600 15657 33609 15691
rect 33609 15657 33643 15691
rect 33643 15657 33652 15691
rect 33600 15648 33652 15657
rect 38016 15691 38068 15700
rect 38016 15657 38025 15691
rect 38025 15657 38059 15691
rect 38059 15657 38068 15691
rect 38016 15648 38068 15657
rect 2412 15580 2464 15632
rect 20904 15580 20956 15632
rect 21456 15580 21508 15632
rect 21916 15580 21968 15632
rect 23112 15623 23164 15632
rect 23112 15589 23121 15623
rect 23121 15589 23155 15623
rect 23155 15589 23164 15623
rect 23112 15580 23164 15589
rect 17224 15555 17276 15564
rect 17224 15521 17233 15555
rect 17233 15521 17267 15555
rect 17267 15521 17276 15555
rect 17224 15512 17276 15521
rect 18696 15555 18748 15564
rect 18696 15521 18705 15555
rect 18705 15521 18739 15555
rect 18739 15521 18748 15555
rect 18696 15512 18748 15521
rect 19524 15555 19576 15564
rect 19524 15521 19533 15555
rect 19533 15521 19567 15555
rect 19567 15521 19576 15555
rect 19524 15512 19576 15521
rect 19800 15512 19852 15564
rect 20628 15487 20680 15496
rect 20628 15453 20637 15487
rect 20637 15453 20671 15487
rect 20671 15453 20680 15487
rect 20628 15444 20680 15453
rect 21640 15512 21692 15564
rect 28540 15580 28592 15632
rect 26424 15512 26476 15564
rect 27896 15512 27948 15564
rect 22192 15487 22244 15496
rect 22192 15453 22201 15487
rect 22201 15453 22235 15487
rect 22235 15453 22244 15487
rect 22192 15444 22244 15453
rect 23296 15487 23348 15496
rect 23296 15453 23305 15487
rect 23305 15453 23339 15487
rect 23339 15453 23348 15487
rect 23296 15444 23348 15453
rect 23664 15444 23716 15496
rect 28264 15444 28316 15496
rect 31668 15580 31720 15632
rect 29092 15512 29144 15564
rect 1952 15308 2004 15360
rect 16212 15419 16264 15428
rect 16212 15385 16221 15419
rect 16221 15385 16255 15419
rect 16255 15385 16264 15419
rect 16212 15376 16264 15385
rect 17408 15419 17460 15428
rect 17408 15385 17417 15419
rect 17417 15385 17451 15419
rect 17451 15385 17460 15419
rect 17408 15376 17460 15385
rect 17776 15376 17828 15428
rect 18604 15419 18656 15428
rect 18604 15385 18613 15419
rect 18613 15385 18647 15419
rect 18647 15385 18656 15419
rect 18604 15376 18656 15385
rect 18880 15376 18932 15428
rect 19524 15376 19576 15428
rect 18788 15308 18840 15360
rect 19708 15376 19760 15428
rect 25228 15419 25280 15428
rect 25228 15385 25237 15419
rect 25237 15385 25271 15419
rect 25271 15385 25280 15419
rect 25228 15376 25280 15385
rect 25412 15376 25464 15428
rect 25872 15419 25924 15428
rect 25872 15385 25881 15419
rect 25881 15385 25915 15419
rect 25915 15385 25924 15419
rect 25872 15376 25924 15385
rect 27528 15419 27580 15428
rect 27528 15385 27537 15419
rect 27537 15385 27571 15419
rect 27571 15385 27580 15419
rect 27528 15376 27580 15385
rect 29828 15444 29880 15496
rect 29920 15487 29972 15496
rect 29920 15453 29929 15487
rect 29929 15453 29963 15487
rect 29963 15453 29972 15487
rect 29920 15444 29972 15453
rect 33508 15487 33560 15496
rect 33508 15453 33517 15487
rect 33517 15453 33551 15487
rect 33551 15453 33560 15487
rect 33508 15444 33560 15453
rect 37832 15487 37884 15496
rect 37832 15453 37841 15487
rect 37841 15453 37875 15487
rect 37875 15453 37884 15487
rect 37832 15444 37884 15453
rect 28540 15376 28592 15428
rect 37740 15376 37792 15428
rect 21088 15308 21140 15360
rect 21272 15351 21324 15360
rect 21272 15317 21281 15351
rect 21281 15317 21315 15351
rect 21315 15317 21324 15351
rect 21272 15308 21324 15317
rect 21732 15308 21784 15360
rect 22376 15308 22428 15360
rect 26976 15351 27028 15360
rect 26976 15317 26985 15351
rect 26985 15317 27019 15351
rect 27019 15317 27028 15351
rect 26976 15308 27028 15317
rect 27252 15308 27304 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 16028 15104 16080 15156
rect 16212 15036 16264 15088
rect 14740 15011 14792 15020
rect 14740 14977 14749 15011
rect 14749 14977 14783 15011
rect 14783 14977 14792 15011
rect 14740 14968 14792 14977
rect 18604 15104 18656 15156
rect 17960 15036 18012 15088
rect 19156 15036 19208 15088
rect 20076 15104 20128 15156
rect 22192 15104 22244 15156
rect 22652 15104 22704 15156
rect 20352 15079 20404 15088
rect 16580 14900 16632 14952
rect 15752 14832 15804 14884
rect 16764 14832 16816 14884
rect 19064 14968 19116 15020
rect 20352 15045 20361 15079
rect 20361 15045 20395 15079
rect 20395 15045 20404 15079
rect 20352 15036 20404 15045
rect 20536 15036 20588 15088
rect 20720 15036 20772 15088
rect 23480 15079 23532 15088
rect 23480 15045 23489 15079
rect 23489 15045 23523 15079
rect 23523 15045 23532 15079
rect 28172 15104 28224 15156
rect 23480 15036 23532 15045
rect 24952 15036 25004 15088
rect 25596 15036 25648 15088
rect 29460 15104 29512 15156
rect 31760 15036 31812 15088
rect 16948 14900 17000 14952
rect 17408 14900 17460 14952
rect 18052 14900 18104 14952
rect 18144 14900 18196 14952
rect 20996 14900 21048 14952
rect 22100 14968 22152 15020
rect 24860 14968 24912 15020
rect 25688 15011 25740 15020
rect 17592 14832 17644 14884
rect 21180 14832 21232 14884
rect 21732 14832 21784 14884
rect 22928 14875 22980 14884
rect 22928 14841 22937 14875
rect 22937 14841 22971 14875
rect 22971 14841 22980 14875
rect 22928 14832 22980 14841
rect 24124 14875 24176 14884
rect 24124 14841 24133 14875
rect 24133 14841 24167 14875
rect 24167 14841 24176 14875
rect 24124 14832 24176 14841
rect 25044 14900 25096 14952
rect 25688 14977 25697 15011
rect 25697 14977 25731 15011
rect 25731 14977 25740 15011
rect 25688 14968 25740 14977
rect 26700 14968 26752 15020
rect 28264 14968 28316 15020
rect 28356 14968 28408 15020
rect 28724 15011 28776 15020
rect 28724 14977 28733 15011
rect 28733 14977 28767 15011
rect 28767 14977 28776 15011
rect 28724 14968 28776 14977
rect 28816 14968 28868 15020
rect 31392 15011 31444 15020
rect 26056 14900 26108 14952
rect 27252 14900 27304 14952
rect 26884 14832 26936 14884
rect 19248 14764 19300 14816
rect 23572 14764 23624 14816
rect 23756 14764 23808 14816
rect 26424 14764 26476 14816
rect 28356 14764 28408 14816
rect 28816 14832 28868 14884
rect 29552 14832 29604 14884
rect 30196 14900 30248 14952
rect 31392 14977 31401 15011
rect 31401 14977 31435 15011
rect 31435 14977 31444 15011
rect 31392 14968 31444 14977
rect 31300 14900 31352 14952
rect 29644 14807 29696 14816
rect 29644 14773 29653 14807
rect 29653 14773 29687 14807
rect 29687 14773 29696 14807
rect 29644 14764 29696 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 4068 14560 4120 14612
rect 14004 14560 14056 14612
rect 17500 14560 17552 14612
rect 22100 14560 22152 14612
rect 23296 14560 23348 14612
rect 23664 14560 23716 14612
rect 25688 14560 25740 14612
rect 28816 14560 28868 14612
rect 28908 14560 28960 14612
rect 31760 14603 31812 14612
rect 31760 14569 31769 14603
rect 31769 14569 31803 14603
rect 31803 14569 31812 14603
rect 31760 14560 31812 14569
rect 32312 14603 32364 14612
rect 32312 14569 32321 14603
rect 32321 14569 32355 14603
rect 32355 14569 32364 14603
rect 32312 14560 32364 14569
rect 38108 14560 38160 14612
rect 16120 14492 16172 14544
rect 17224 14492 17276 14544
rect 20628 14492 20680 14544
rect 23112 14535 23164 14544
rect 23112 14501 23121 14535
rect 23121 14501 23155 14535
rect 23155 14501 23164 14535
rect 23112 14492 23164 14501
rect 23940 14492 23992 14544
rect 26792 14492 26844 14544
rect 26976 14492 27028 14544
rect 1584 14399 1636 14408
rect 1584 14365 1593 14399
rect 1593 14365 1627 14399
rect 1627 14365 1636 14399
rect 1584 14356 1636 14365
rect 5540 14356 5592 14408
rect 14096 14356 14148 14408
rect 13728 14220 13780 14272
rect 15752 14331 15804 14340
rect 15752 14297 15761 14331
rect 15761 14297 15795 14331
rect 15795 14297 15804 14331
rect 15752 14288 15804 14297
rect 16120 14288 16172 14340
rect 17040 14356 17092 14408
rect 17408 14356 17460 14408
rect 17592 14424 17644 14476
rect 19984 14424 20036 14476
rect 23572 14467 23624 14476
rect 20076 14356 20128 14408
rect 18052 14288 18104 14340
rect 18236 14331 18288 14340
rect 18236 14297 18245 14331
rect 18245 14297 18279 14331
rect 18279 14297 18288 14331
rect 18236 14288 18288 14297
rect 18880 14331 18932 14340
rect 17408 14220 17460 14272
rect 17592 14263 17644 14272
rect 17592 14229 17601 14263
rect 17601 14229 17635 14263
rect 17635 14229 17644 14263
rect 17592 14220 17644 14229
rect 18880 14297 18889 14331
rect 18889 14297 18923 14331
rect 18923 14297 18932 14331
rect 18880 14288 18932 14297
rect 23572 14433 23581 14467
rect 23581 14433 23615 14467
rect 23615 14433 23624 14467
rect 23572 14424 23624 14433
rect 22008 14356 22060 14408
rect 22100 14399 22152 14408
rect 22100 14365 22109 14399
rect 22109 14365 22143 14399
rect 22143 14365 22152 14399
rect 24308 14424 24360 14476
rect 25412 14424 25464 14476
rect 25964 14424 26016 14476
rect 26240 14424 26292 14476
rect 22100 14356 22152 14365
rect 23756 14399 23808 14408
rect 23756 14365 23765 14399
rect 23765 14365 23799 14399
rect 23799 14365 23808 14399
rect 24584 14399 24636 14408
rect 23756 14356 23808 14365
rect 24584 14365 24593 14399
rect 24593 14365 24627 14399
rect 24627 14365 24636 14399
rect 24584 14356 24636 14365
rect 25504 14356 25556 14408
rect 29368 14492 29420 14544
rect 29460 14492 29512 14544
rect 28908 14424 28960 14476
rect 28448 14356 28500 14408
rect 29184 14399 29236 14408
rect 29184 14365 29193 14399
rect 29193 14365 29227 14399
rect 29227 14365 29236 14399
rect 29184 14356 29236 14365
rect 29368 14356 29420 14408
rect 20996 14331 21048 14340
rect 20996 14297 21005 14331
rect 21005 14297 21039 14331
rect 21039 14297 21048 14331
rect 20996 14288 21048 14297
rect 21088 14331 21140 14340
rect 21088 14297 21097 14331
rect 21097 14297 21131 14331
rect 21131 14297 21140 14331
rect 21088 14288 21140 14297
rect 20076 14220 20128 14272
rect 21732 14288 21784 14340
rect 22100 14220 22152 14272
rect 23204 14220 23256 14272
rect 25596 14220 25648 14272
rect 27252 14288 27304 14340
rect 27436 14331 27488 14340
rect 27436 14297 27445 14331
rect 27445 14297 27479 14331
rect 27479 14297 27488 14331
rect 27436 14288 27488 14297
rect 30104 14356 30156 14408
rect 32036 14356 32088 14408
rect 31576 14288 31628 14340
rect 27620 14220 27672 14272
rect 29000 14220 29052 14272
rect 29552 14220 29604 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 14004 14059 14056 14068
rect 14004 14025 14013 14059
rect 14013 14025 14047 14059
rect 14047 14025 14056 14059
rect 14004 14016 14056 14025
rect 16028 14016 16080 14068
rect 16212 14059 16264 14068
rect 16212 14025 16221 14059
rect 16221 14025 16255 14059
rect 16255 14025 16264 14059
rect 16212 14016 16264 14025
rect 16304 14016 16356 14068
rect 19984 14016 20036 14068
rect 20076 14016 20128 14068
rect 16396 13948 16448 14000
rect 18972 13948 19024 14000
rect 20812 13948 20864 14000
rect 23480 14016 23532 14068
rect 23848 13991 23900 14000
rect 23848 13957 23857 13991
rect 23857 13957 23891 13991
rect 23891 13957 23900 13991
rect 23848 13948 23900 13957
rect 25228 14016 25280 14068
rect 26884 14016 26936 14068
rect 26976 14016 27028 14068
rect 28264 14016 28316 14068
rect 28172 13948 28224 14000
rect 37372 14016 37424 14068
rect 28540 13948 28592 14000
rect 28724 13948 28776 14000
rect 29460 13948 29512 14000
rect 31208 13991 31260 14000
rect 31208 13957 31217 13991
rect 31217 13957 31251 13991
rect 31251 13957 31260 13991
rect 31208 13948 31260 13957
rect 13728 13880 13780 13932
rect 16580 13880 16632 13932
rect 17132 13880 17184 13932
rect 17500 13923 17552 13932
rect 17500 13889 17509 13923
rect 17509 13889 17543 13923
rect 17543 13889 17552 13923
rect 17500 13880 17552 13889
rect 19064 13880 19116 13932
rect 20628 13880 20680 13932
rect 21640 13880 21692 13932
rect 23296 13880 23348 13932
rect 25320 13880 25372 13932
rect 16304 13812 16356 13864
rect 16948 13855 17000 13864
rect 16948 13821 16957 13855
rect 16957 13821 16991 13855
rect 16991 13821 17000 13855
rect 16948 13812 17000 13821
rect 17408 13812 17460 13864
rect 19340 13812 19392 13864
rect 10876 13744 10928 13796
rect 17960 13744 18012 13796
rect 20904 13744 20956 13796
rect 15568 13719 15620 13728
rect 15568 13685 15577 13719
rect 15577 13685 15611 13719
rect 15611 13685 15620 13719
rect 15568 13676 15620 13685
rect 15752 13676 15804 13728
rect 19432 13676 19484 13728
rect 19524 13676 19576 13728
rect 23480 13812 23532 13864
rect 23756 13812 23808 13864
rect 23388 13744 23440 13796
rect 25136 13855 25188 13864
rect 25136 13821 25145 13855
rect 25145 13821 25179 13855
rect 25179 13821 25188 13855
rect 25136 13812 25188 13821
rect 25412 13812 25464 13864
rect 25688 13855 25740 13864
rect 25688 13821 25697 13855
rect 25697 13821 25731 13855
rect 25731 13821 25740 13855
rect 25688 13812 25740 13821
rect 26056 13812 26108 13864
rect 26608 13812 26660 13864
rect 27160 13812 27212 13864
rect 27620 13855 27672 13864
rect 27620 13821 27629 13855
rect 27629 13821 27663 13855
rect 27663 13821 27672 13855
rect 27620 13812 27672 13821
rect 27988 13880 28040 13932
rect 29184 13812 29236 13864
rect 22744 13719 22796 13728
rect 22744 13685 22753 13719
rect 22753 13685 22787 13719
rect 22787 13685 22796 13719
rect 22744 13676 22796 13685
rect 24860 13676 24912 13728
rect 28172 13744 28224 13796
rect 28908 13787 28960 13796
rect 28908 13753 28917 13787
rect 28917 13753 28951 13787
rect 28951 13753 28960 13787
rect 28908 13744 28960 13753
rect 29000 13744 29052 13796
rect 29828 13880 29880 13932
rect 32588 13880 32640 13932
rect 38292 13923 38344 13932
rect 38292 13889 38301 13923
rect 38301 13889 38335 13923
rect 38335 13889 38344 13923
rect 38292 13880 38344 13889
rect 29920 13812 29972 13864
rect 31116 13855 31168 13864
rect 31116 13821 31125 13855
rect 31125 13821 31159 13855
rect 31159 13821 31168 13855
rect 31116 13812 31168 13821
rect 31300 13744 31352 13796
rect 31760 13744 31812 13796
rect 35532 13744 35584 13796
rect 27252 13676 27304 13728
rect 29736 13676 29788 13728
rect 30196 13676 30248 13728
rect 30472 13676 30524 13728
rect 33508 13676 33560 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 13728 13515 13780 13524
rect 13728 13481 13737 13515
rect 13737 13481 13771 13515
rect 13771 13481 13780 13515
rect 13728 13472 13780 13481
rect 15660 13472 15712 13524
rect 18512 13404 18564 13456
rect 2320 13336 2372 13388
rect 10876 13336 10928 13388
rect 15752 13336 15804 13388
rect 17500 13336 17552 13388
rect 18236 13336 18288 13388
rect 21456 13472 21508 13524
rect 24124 13472 24176 13524
rect 18788 13404 18840 13456
rect 22928 13404 22980 13456
rect 23020 13404 23072 13456
rect 19524 13379 19576 13388
rect 19524 13345 19533 13379
rect 19533 13345 19567 13379
rect 19567 13345 19576 13379
rect 19524 13336 19576 13345
rect 20812 13379 20864 13388
rect 20812 13345 20821 13379
rect 20821 13345 20855 13379
rect 20855 13345 20864 13379
rect 20812 13336 20864 13345
rect 21180 13379 21232 13388
rect 21180 13345 21189 13379
rect 21189 13345 21223 13379
rect 21223 13345 21232 13379
rect 21180 13336 21232 13345
rect 21916 13336 21968 13388
rect 23112 13336 23164 13388
rect 23296 13379 23348 13388
rect 23296 13345 23305 13379
rect 23305 13345 23339 13379
rect 23339 13345 23348 13379
rect 23296 13336 23348 13345
rect 13360 13268 13412 13320
rect 13820 13200 13872 13252
rect 17684 13268 17736 13320
rect 27160 13472 27212 13524
rect 28908 13472 28960 13524
rect 30472 13472 30524 13524
rect 30564 13472 30616 13524
rect 31668 13515 31720 13524
rect 31668 13481 31677 13515
rect 31677 13481 31711 13515
rect 31711 13481 31720 13515
rect 31668 13472 31720 13481
rect 25412 13404 25464 13456
rect 25780 13336 25832 13388
rect 27252 13336 27304 13388
rect 28172 13404 28224 13456
rect 29736 13404 29788 13456
rect 29828 13404 29880 13456
rect 31760 13404 31812 13456
rect 27620 13336 27672 13388
rect 29000 13336 29052 13388
rect 17316 13243 17368 13252
rect 17316 13209 17325 13243
rect 17325 13209 17359 13243
rect 17359 13209 17368 13243
rect 17316 13200 17368 13209
rect 18052 13243 18104 13252
rect 18052 13209 18061 13243
rect 18061 13209 18095 13243
rect 18095 13209 18104 13243
rect 18052 13200 18104 13209
rect 18328 13200 18380 13252
rect 18788 13200 18840 13252
rect 20904 13243 20956 13252
rect 15844 13132 15896 13184
rect 17224 13175 17276 13184
rect 17224 13141 17233 13175
rect 17233 13141 17267 13175
rect 17267 13141 17276 13175
rect 17224 13132 17276 13141
rect 19248 13132 19300 13184
rect 20904 13209 20913 13243
rect 20913 13209 20947 13243
rect 20947 13209 20956 13243
rect 20904 13200 20956 13209
rect 23204 13243 23256 13252
rect 23204 13209 23213 13243
rect 23213 13209 23247 13243
rect 23247 13209 23256 13243
rect 23204 13200 23256 13209
rect 25688 13243 25740 13252
rect 25688 13209 25697 13243
rect 25697 13209 25731 13243
rect 25731 13209 25740 13243
rect 25688 13200 25740 13209
rect 25964 13200 26016 13252
rect 21180 13132 21232 13184
rect 24768 13132 24820 13184
rect 25872 13132 25924 13184
rect 27528 13200 27580 13252
rect 30472 13311 30524 13320
rect 30472 13277 30481 13311
rect 30481 13277 30515 13311
rect 30515 13277 30524 13311
rect 30472 13268 30524 13277
rect 31024 13268 31076 13320
rect 32128 13268 32180 13320
rect 32864 13311 32916 13320
rect 29184 13243 29236 13252
rect 29184 13209 29193 13243
rect 29193 13209 29227 13243
rect 29227 13209 29236 13243
rect 29184 13200 29236 13209
rect 29644 13200 29696 13252
rect 30288 13200 30340 13252
rect 31392 13132 31444 13184
rect 32864 13277 32873 13311
rect 32873 13277 32907 13311
rect 32907 13277 32916 13311
rect 32864 13268 32916 13277
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 13360 12971 13412 12980
rect 13360 12937 13369 12971
rect 13369 12937 13403 12971
rect 13403 12937 13412 12971
rect 13360 12928 13412 12937
rect 14464 12971 14516 12980
rect 14464 12937 14473 12971
rect 14473 12937 14507 12971
rect 14507 12937 14516 12971
rect 14464 12928 14516 12937
rect 17316 12928 17368 12980
rect 15660 12903 15712 12912
rect 15660 12869 15669 12903
rect 15669 12869 15703 12903
rect 15703 12869 15712 12903
rect 15660 12860 15712 12869
rect 15844 12860 15896 12912
rect 16028 12860 16080 12912
rect 17868 12928 17920 12980
rect 4068 12792 4120 12844
rect 14924 12835 14976 12844
rect 14924 12801 14933 12835
rect 14933 12801 14967 12835
rect 14967 12801 14976 12835
rect 14924 12792 14976 12801
rect 17592 12860 17644 12912
rect 17040 12724 17092 12776
rect 17316 12724 17368 12776
rect 17868 12767 17920 12776
rect 17868 12733 17877 12767
rect 17877 12733 17911 12767
rect 17911 12733 17920 12767
rect 17868 12724 17920 12733
rect 19340 12860 19392 12912
rect 22744 12928 22796 12980
rect 23204 12928 23256 12980
rect 21456 12903 21508 12912
rect 21456 12869 21465 12903
rect 21465 12869 21499 12903
rect 21499 12869 21508 12903
rect 21456 12860 21508 12869
rect 19064 12767 19116 12776
rect 15752 12656 15804 12708
rect 19064 12733 19073 12767
rect 19073 12733 19107 12767
rect 19107 12733 19116 12767
rect 19064 12724 19116 12733
rect 20168 12724 20220 12776
rect 20536 12724 20588 12776
rect 18880 12656 18932 12708
rect 1676 12631 1728 12640
rect 1676 12597 1685 12631
rect 1685 12597 1719 12631
rect 1719 12597 1728 12631
rect 1676 12588 1728 12597
rect 16488 12588 16540 12640
rect 20076 12588 20128 12640
rect 20260 12656 20312 12708
rect 23480 12860 23532 12912
rect 25320 12860 25372 12912
rect 25780 12860 25832 12912
rect 30288 12928 30340 12980
rect 26976 12860 27028 12912
rect 29828 12860 29880 12912
rect 32956 12903 33008 12912
rect 32956 12869 32965 12903
rect 32965 12869 32999 12903
rect 32999 12869 33008 12903
rect 32956 12860 33008 12869
rect 23020 12767 23072 12776
rect 23020 12733 23029 12767
rect 23029 12733 23063 12767
rect 23063 12733 23072 12767
rect 23020 12724 23072 12733
rect 23388 12724 23440 12776
rect 24768 12724 24820 12776
rect 28908 12792 28960 12844
rect 29000 12835 29052 12844
rect 29000 12801 29009 12835
rect 29009 12801 29043 12835
rect 29043 12801 29052 12835
rect 29000 12792 29052 12801
rect 29644 12833 29696 12844
rect 29644 12799 29653 12833
rect 29653 12799 29687 12833
rect 29687 12799 29696 12833
rect 29644 12792 29696 12799
rect 31576 12835 31628 12844
rect 25872 12724 25924 12776
rect 26056 12724 26108 12776
rect 29184 12724 29236 12776
rect 30656 12724 30708 12776
rect 31576 12801 31585 12835
rect 31585 12801 31619 12835
rect 31619 12801 31628 12835
rect 31576 12792 31628 12801
rect 33600 12792 33652 12844
rect 31852 12724 31904 12776
rect 27896 12656 27948 12708
rect 28448 12656 28500 12708
rect 25596 12588 25648 12640
rect 26056 12588 26108 12640
rect 26332 12588 26384 12640
rect 37648 12588 37700 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 13728 12384 13780 12436
rect 14280 12384 14332 12436
rect 17868 12316 17920 12368
rect 18144 12384 18196 12436
rect 19156 12384 19208 12436
rect 1860 12248 1912 12300
rect 8300 12248 8352 12300
rect 14464 12223 14516 12232
rect 14464 12189 14473 12223
rect 14473 12189 14507 12223
rect 14507 12189 14516 12223
rect 14464 12180 14516 12189
rect 15844 12180 15896 12232
rect 16856 12248 16908 12300
rect 17592 12248 17644 12300
rect 19340 12316 19392 12368
rect 18236 12248 18288 12300
rect 24124 12384 24176 12436
rect 24492 12384 24544 12436
rect 26332 12384 26384 12436
rect 26424 12384 26476 12436
rect 28448 12384 28500 12436
rect 28540 12384 28592 12436
rect 31760 12427 31812 12436
rect 31760 12393 31769 12427
rect 31769 12393 31803 12427
rect 31803 12393 31812 12427
rect 31760 12384 31812 12393
rect 21916 12316 21968 12368
rect 16028 12180 16080 12232
rect 20720 12248 20772 12300
rect 22928 12316 22980 12368
rect 27436 12316 27488 12368
rect 23112 12291 23164 12300
rect 23112 12257 23121 12291
rect 23121 12257 23155 12291
rect 23155 12257 23164 12291
rect 23112 12248 23164 12257
rect 23572 12248 23624 12300
rect 24584 12248 24636 12300
rect 25136 12248 25188 12300
rect 25872 12248 25924 12300
rect 26148 12291 26200 12300
rect 26148 12257 26157 12291
rect 26157 12257 26191 12291
rect 26191 12257 26200 12291
rect 26148 12248 26200 12257
rect 29000 12248 29052 12300
rect 31576 12316 31628 12368
rect 32404 12291 32456 12300
rect 32404 12257 32413 12291
rect 32413 12257 32447 12291
rect 32447 12257 32456 12291
rect 32404 12248 32456 12257
rect 29920 12223 29972 12232
rect 29920 12189 29929 12223
rect 29929 12189 29963 12223
rect 29963 12189 29972 12223
rect 29920 12180 29972 12189
rect 30380 12223 30432 12232
rect 30380 12189 30389 12223
rect 30389 12189 30423 12223
rect 30423 12189 30432 12223
rect 30380 12180 30432 12189
rect 16304 12112 16356 12164
rect 16948 12155 17000 12164
rect 16948 12121 16957 12155
rect 16957 12121 16991 12155
rect 16991 12121 17000 12155
rect 16948 12112 17000 12121
rect 18512 12112 18564 12164
rect 18880 12112 18932 12164
rect 21180 12112 21232 12164
rect 23756 12112 23808 12164
rect 24584 12155 24636 12164
rect 24584 12121 24593 12155
rect 24593 12121 24627 12155
rect 24627 12121 24636 12155
rect 24584 12112 24636 12121
rect 26424 12155 26476 12164
rect 14924 12044 14976 12096
rect 15200 12087 15252 12096
rect 15200 12053 15209 12087
rect 15209 12053 15243 12087
rect 15243 12053 15252 12087
rect 15200 12044 15252 12053
rect 19984 12044 20036 12096
rect 20812 12044 20864 12096
rect 23572 12044 23624 12096
rect 26424 12121 26433 12155
rect 26433 12121 26467 12155
rect 26467 12121 26476 12155
rect 26424 12112 26476 12121
rect 27528 12112 27580 12164
rect 28356 12112 28408 12164
rect 28448 12155 28500 12164
rect 28448 12121 28457 12155
rect 28457 12121 28491 12155
rect 28491 12121 28500 12155
rect 28448 12112 28500 12121
rect 29000 12155 29052 12164
rect 29000 12121 29009 12155
rect 29009 12121 29043 12155
rect 29043 12121 29052 12155
rect 30472 12155 30524 12164
rect 29000 12112 29052 12121
rect 30472 12121 30481 12155
rect 30481 12121 30515 12155
rect 30515 12121 30524 12155
rect 30472 12112 30524 12121
rect 29092 12044 29144 12096
rect 30104 12044 30156 12096
rect 31668 12223 31720 12232
rect 31668 12189 31677 12223
rect 31677 12189 31711 12223
rect 31711 12189 31720 12223
rect 31668 12180 31720 12189
rect 34428 12180 34480 12232
rect 37556 12112 37608 12164
rect 37832 12044 37884 12096
rect 37924 12087 37976 12096
rect 37924 12053 37933 12087
rect 37933 12053 37967 12087
rect 37967 12053 37976 12087
rect 37924 12044 37976 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 6552 11883 6604 11892
rect 6552 11849 6561 11883
rect 6561 11849 6595 11883
rect 6595 11849 6604 11883
rect 6552 11840 6604 11849
rect 15200 11840 15252 11892
rect 15752 11772 15804 11824
rect 17684 11815 17736 11824
rect 14280 11747 14332 11756
rect 14280 11713 14289 11747
rect 14289 11713 14323 11747
rect 14323 11713 14332 11747
rect 14280 11704 14332 11713
rect 15568 11704 15620 11756
rect 16396 11636 16448 11688
rect 17684 11781 17693 11815
rect 17693 11781 17727 11815
rect 17727 11781 17736 11815
rect 17684 11772 17736 11781
rect 17960 11772 18012 11824
rect 20260 11840 20312 11892
rect 22008 11840 22060 11892
rect 20812 11772 20864 11824
rect 20996 11815 21048 11824
rect 20996 11781 21005 11815
rect 21005 11781 21039 11815
rect 21039 11781 21048 11815
rect 20996 11772 21048 11781
rect 22100 11772 22152 11824
rect 19800 11747 19852 11756
rect 19800 11713 19809 11747
rect 19809 11713 19843 11747
rect 19843 11713 19852 11747
rect 19800 11704 19852 11713
rect 23296 11840 23348 11892
rect 24492 11840 24544 11892
rect 23940 11772 23992 11824
rect 24308 11772 24360 11824
rect 24860 11815 24912 11824
rect 24860 11781 24869 11815
rect 24869 11781 24903 11815
rect 24903 11781 24912 11815
rect 24860 11772 24912 11781
rect 25136 11772 25188 11824
rect 26240 11772 26292 11824
rect 28724 11840 28776 11892
rect 28264 11704 28316 11756
rect 29092 11704 29144 11756
rect 30840 11840 30892 11892
rect 29736 11772 29788 11824
rect 29828 11747 29880 11756
rect 29828 11713 29837 11747
rect 29837 11713 29871 11747
rect 29871 11713 29880 11747
rect 29828 11704 29880 11713
rect 30288 11704 30340 11756
rect 31208 11840 31260 11892
rect 15660 11611 15712 11620
rect 15660 11577 15669 11611
rect 15669 11577 15703 11611
rect 15703 11577 15712 11611
rect 15660 11568 15712 11577
rect 16028 11568 16080 11620
rect 17960 11636 18012 11688
rect 18604 11636 18656 11688
rect 21824 11636 21876 11688
rect 27436 11636 27488 11688
rect 27528 11636 27580 11688
rect 31208 11704 31260 11756
rect 33416 11704 33468 11756
rect 38200 11747 38252 11756
rect 38200 11713 38209 11747
rect 38209 11713 38243 11747
rect 38243 11713 38252 11747
rect 38200 11704 38252 11713
rect 31852 11636 31904 11688
rect 38384 11636 38436 11688
rect 18788 11568 18840 11620
rect 5724 11543 5776 11552
rect 5724 11509 5733 11543
rect 5733 11509 5767 11543
rect 5767 11509 5776 11543
rect 5724 11500 5776 11509
rect 17040 11500 17092 11552
rect 17408 11500 17460 11552
rect 21456 11568 21508 11620
rect 20076 11500 20128 11552
rect 21916 11500 21968 11552
rect 22008 11500 22060 11552
rect 28172 11568 28224 11620
rect 28540 11568 28592 11620
rect 31116 11568 31168 11620
rect 38016 11611 38068 11620
rect 38016 11577 38025 11611
rect 38025 11577 38059 11611
rect 38059 11577 38068 11611
rect 38016 11568 38068 11577
rect 29092 11500 29144 11552
rect 31208 11500 31260 11552
rect 37372 11500 37424 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 15476 11296 15528 11348
rect 15660 11296 15712 11348
rect 16396 11203 16448 11212
rect 16396 11169 16405 11203
rect 16405 11169 16439 11203
rect 16439 11169 16448 11203
rect 16396 11160 16448 11169
rect 17408 11160 17460 11212
rect 5540 11092 5592 11144
rect 6368 11092 6420 11144
rect 13360 11092 13412 11144
rect 13544 11135 13596 11144
rect 13544 11101 13553 11135
rect 13553 11101 13587 11135
rect 13587 11101 13596 11135
rect 13544 11092 13596 11101
rect 14280 11135 14332 11144
rect 14280 11101 14289 11135
rect 14289 11101 14323 11135
rect 14323 11101 14332 11135
rect 14280 11092 14332 11101
rect 20812 11228 20864 11280
rect 20996 11296 21048 11348
rect 22836 11228 22888 11280
rect 18328 11160 18380 11212
rect 18604 11203 18656 11212
rect 18604 11169 18613 11203
rect 18613 11169 18647 11203
rect 18647 11169 18656 11203
rect 18604 11160 18656 11169
rect 20168 11160 20220 11212
rect 18052 11092 18104 11144
rect 15016 11067 15068 11076
rect 15016 11033 15025 11067
rect 15025 11033 15059 11067
rect 15059 11033 15068 11067
rect 15016 11024 15068 11033
rect 15108 11067 15160 11076
rect 15108 11033 15117 11067
rect 15117 11033 15151 11067
rect 15151 11033 15160 11067
rect 15108 11024 15160 11033
rect 16488 11067 16540 11076
rect 16488 11033 16497 11067
rect 16497 11033 16531 11067
rect 16531 11033 16540 11067
rect 16488 11024 16540 11033
rect 14280 10956 14332 11008
rect 15200 10956 15252 11008
rect 15476 10956 15528 11008
rect 17960 11024 18012 11076
rect 18328 11067 18380 11076
rect 18328 11033 18337 11067
rect 18337 11033 18371 11067
rect 18371 11033 18380 11067
rect 18328 11024 18380 11033
rect 19064 11024 19116 11076
rect 16764 10956 16816 11008
rect 17868 10956 17920 11008
rect 20076 11067 20128 11076
rect 20076 11033 20085 11067
rect 20085 11033 20119 11067
rect 20119 11033 20128 11067
rect 22008 11160 22060 11212
rect 23480 11228 23532 11280
rect 23848 11296 23900 11348
rect 27068 11339 27120 11348
rect 27068 11305 27077 11339
rect 27077 11305 27111 11339
rect 27111 11305 27120 11339
rect 27068 11296 27120 11305
rect 27252 11296 27304 11348
rect 29092 11296 29144 11348
rect 30472 11339 30524 11348
rect 30472 11305 30481 11339
rect 30481 11305 30515 11339
rect 30515 11305 30524 11339
rect 30472 11296 30524 11305
rect 31852 11296 31904 11348
rect 24584 11228 24636 11280
rect 27712 11271 27764 11280
rect 27712 11237 27721 11271
rect 27721 11237 27755 11271
rect 27755 11237 27764 11271
rect 27712 11228 27764 11237
rect 21456 11135 21508 11144
rect 21456 11101 21465 11135
rect 21465 11101 21499 11135
rect 21499 11101 21508 11135
rect 21456 11092 21508 11101
rect 23756 11092 23808 11144
rect 20076 11024 20128 11033
rect 21640 11024 21692 11076
rect 22652 11067 22704 11076
rect 22652 11033 22661 11067
rect 22661 11033 22695 11067
rect 22695 11033 22704 11067
rect 22652 11024 22704 11033
rect 23204 11067 23256 11076
rect 23204 11033 23213 11067
rect 23213 11033 23247 11067
rect 23247 11033 23256 11067
rect 23204 11024 23256 11033
rect 24952 11160 25004 11212
rect 25228 11203 25280 11212
rect 25228 11169 25237 11203
rect 25237 11169 25271 11203
rect 25271 11169 25280 11203
rect 25228 11160 25280 11169
rect 26148 11203 26200 11212
rect 26148 11169 26157 11203
rect 26157 11169 26191 11203
rect 26191 11169 26200 11203
rect 26148 11160 26200 11169
rect 26240 11160 26292 11212
rect 29920 11228 29972 11280
rect 34796 11296 34848 11348
rect 28356 11160 28408 11212
rect 29736 11160 29788 11212
rect 30472 11160 30524 11212
rect 31668 11160 31720 11212
rect 24584 11067 24636 11076
rect 24584 11033 24593 11067
rect 24593 11033 24627 11067
rect 24627 11033 24636 11067
rect 25136 11067 25188 11076
rect 24584 11024 24636 11033
rect 25136 11033 25145 11067
rect 25145 11033 25179 11067
rect 25179 11033 25188 11067
rect 25136 11024 25188 11033
rect 25228 11024 25280 11076
rect 20720 10956 20772 11008
rect 21732 10956 21784 11008
rect 28724 11092 28776 11144
rect 29092 11135 29144 11144
rect 29092 11101 29101 11135
rect 29101 11101 29135 11135
rect 29135 11101 29144 11135
rect 29092 11092 29144 11101
rect 29184 11092 29236 11144
rect 29920 11135 29972 11144
rect 29920 11101 29929 11135
rect 29929 11101 29963 11135
rect 29963 11101 29972 11135
rect 29920 11092 29972 11101
rect 30564 11135 30616 11144
rect 30564 11101 30573 11135
rect 30573 11101 30607 11135
rect 30607 11101 30616 11135
rect 30564 11092 30616 11101
rect 27804 11024 27856 11076
rect 30288 11024 30340 11076
rect 26792 10956 26844 11008
rect 29184 10956 29236 11008
rect 29644 10956 29696 11008
rect 33876 11024 33928 11076
rect 34520 11024 34572 11076
rect 35808 11024 35860 11076
rect 36084 11067 36136 11076
rect 36084 11033 36093 11067
rect 36093 11033 36127 11067
rect 36127 11033 36136 11067
rect 36084 11024 36136 11033
rect 36820 11024 36872 11076
rect 36912 11024 36964 11076
rect 38108 11024 38160 11076
rect 30932 10956 30984 11008
rect 32864 10956 32916 11008
rect 35716 10956 35768 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 5724 10616 5776 10668
rect 21548 10752 21600 10804
rect 28172 10752 28224 10804
rect 29828 10752 29880 10804
rect 30104 10752 30156 10804
rect 14648 10684 14700 10736
rect 18512 10727 18564 10736
rect 18512 10693 18521 10727
rect 18521 10693 18555 10727
rect 18555 10693 18564 10727
rect 18512 10684 18564 10693
rect 19064 10727 19116 10736
rect 19064 10693 19073 10727
rect 19073 10693 19107 10727
rect 19107 10693 19116 10727
rect 19064 10684 19116 10693
rect 19340 10684 19392 10736
rect 20076 10684 20128 10736
rect 16120 10659 16172 10668
rect 16120 10625 16129 10659
rect 16129 10625 16163 10659
rect 16163 10625 16172 10659
rect 16120 10616 16172 10625
rect 17040 10616 17092 10668
rect 20260 10659 20312 10668
rect 20260 10625 20269 10659
rect 20269 10625 20303 10659
rect 20303 10625 20312 10659
rect 20260 10616 20312 10625
rect 15016 10591 15068 10600
rect 15016 10557 15025 10591
rect 15025 10557 15059 10591
rect 15059 10557 15068 10591
rect 15016 10548 15068 10557
rect 17224 10591 17276 10600
rect 17224 10557 17233 10591
rect 17233 10557 17267 10591
rect 17267 10557 17276 10591
rect 17224 10548 17276 10557
rect 15108 10480 15160 10532
rect 15844 10480 15896 10532
rect 18236 10548 18288 10600
rect 18420 10591 18472 10600
rect 18420 10557 18429 10591
rect 18429 10557 18463 10591
rect 18463 10557 18472 10591
rect 19616 10591 19668 10600
rect 18420 10548 18472 10557
rect 19616 10557 19625 10591
rect 19625 10557 19659 10591
rect 19659 10557 19668 10591
rect 19616 10548 19668 10557
rect 20812 10591 20864 10600
rect 20812 10557 20821 10591
rect 20821 10557 20855 10591
rect 20855 10557 20864 10591
rect 20812 10548 20864 10557
rect 17776 10523 17828 10532
rect 17776 10489 17785 10523
rect 17785 10489 17819 10523
rect 17819 10489 17828 10523
rect 17776 10480 17828 10489
rect 18144 10480 18196 10532
rect 22560 10684 22612 10736
rect 22836 10684 22888 10736
rect 23664 10684 23716 10736
rect 25044 10684 25096 10736
rect 25412 10727 25464 10736
rect 25412 10693 25421 10727
rect 25421 10693 25455 10727
rect 25455 10693 25464 10727
rect 25412 10684 25464 10693
rect 27804 10684 27856 10736
rect 29736 10684 29788 10736
rect 22008 10659 22060 10668
rect 22008 10625 22017 10659
rect 22017 10625 22051 10659
rect 22051 10625 22060 10659
rect 22008 10616 22060 10625
rect 21548 10548 21600 10600
rect 22652 10548 22704 10600
rect 24124 10480 24176 10532
rect 1676 10455 1728 10464
rect 1676 10421 1685 10455
rect 1685 10421 1719 10455
rect 1719 10421 1728 10455
rect 1676 10412 1728 10421
rect 13360 10412 13412 10464
rect 13820 10455 13872 10464
rect 13820 10421 13829 10455
rect 13829 10421 13863 10455
rect 13863 10421 13872 10455
rect 13820 10412 13872 10421
rect 16120 10412 16172 10464
rect 20076 10412 20128 10464
rect 20260 10412 20312 10464
rect 22100 10412 22152 10464
rect 22284 10455 22336 10464
rect 22284 10421 22314 10455
rect 22314 10421 22336 10455
rect 22284 10412 22336 10421
rect 22652 10412 22704 10464
rect 27160 10548 27212 10600
rect 26424 10480 26476 10532
rect 30656 10616 30708 10668
rect 33692 10616 33744 10668
rect 34428 10616 34480 10668
rect 34704 10548 34756 10600
rect 38292 10591 38344 10600
rect 38292 10557 38301 10591
rect 38301 10557 38335 10591
rect 38335 10557 38344 10591
rect 38292 10548 38344 10557
rect 29920 10480 29972 10532
rect 35624 10480 35676 10532
rect 30104 10412 30156 10464
rect 30288 10412 30340 10464
rect 30564 10412 30616 10464
rect 32404 10455 32456 10464
rect 32404 10421 32413 10455
rect 32413 10421 32447 10455
rect 32447 10421 32456 10455
rect 32404 10412 32456 10421
rect 33876 10455 33928 10464
rect 33876 10421 33885 10455
rect 33885 10421 33919 10455
rect 33919 10421 33928 10455
rect 33876 10412 33928 10421
rect 35716 10412 35768 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 14648 10251 14700 10260
rect 14648 10217 14657 10251
rect 14657 10217 14691 10251
rect 14691 10217 14700 10251
rect 14648 10208 14700 10217
rect 14740 10208 14792 10260
rect 18420 10208 18472 10260
rect 18788 10251 18840 10260
rect 18788 10217 18797 10251
rect 18797 10217 18831 10251
rect 18831 10217 18840 10251
rect 18788 10208 18840 10217
rect 19616 10208 19668 10260
rect 21824 10208 21876 10260
rect 22192 10208 22244 10260
rect 22744 10208 22796 10260
rect 23112 10208 23164 10260
rect 14096 10140 14148 10192
rect 15660 10072 15712 10124
rect 15844 10115 15896 10124
rect 15844 10081 15853 10115
rect 15853 10081 15887 10115
rect 15887 10081 15896 10115
rect 15844 10072 15896 10081
rect 18880 10140 18932 10192
rect 20536 10140 20588 10192
rect 21916 10140 21968 10192
rect 22560 10140 22612 10192
rect 24308 10140 24360 10192
rect 24860 10208 24912 10260
rect 26148 10208 26200 10260
rect 29644 10208 29696 10260
rect 30196 10208 30248 10260
rect 36912 10208 36964 10260
rect 37648 10251 37700 10260
rect 37648 10217 37657 10251
rect 37657 10217 37691 10251
rect 37691 10217 37700 10251
rect 37648 10208 37700 10217
rect 38292 10251 38344 10260
rect 38292 10217 38301 10251
rect 38301 10217 38335 10251
rect 38335 10217 38344 10251
rect 38292 10208 38344 10217
rect 17408 10072 17460 10124
rect 20812 10115 20864 10124
rect 12900 9868 12952 9920
rect 16580 10047 16632 10056
rect 16580 10013 16589 10047
rect 16589 10013 16623 10047
rect 16623 10013 16632 10047
rect 16580 10004 16632 10013
rect 20812 10081 20821 10115
rect 20821 10081 20855 10115
rect 20855 10081 20864 10115
rect 20812 10072 20864 10081
rect 21824 10072 21876 10124
rect 22192 10072 22244 10124
rect 25228 10072 25280 10124
rect 26884 10140 26936 10192
rect 29000 10140 29052 10192
rect 29460 10140 29512 10192
rect 30656 10140 30708 10192
rect 20076 10004 20128 10056
rect 15660 9936 15712 9988
rect 17776 9979 17828 9988
rect 15108 9868 15160 9920
rect 17776 9945 17785 9979
rect 17785 9945 17819 9979
rect 17819 9945 17828 9979
rect 17776 9936 17828 9945
rect 21916 10004 21968 10056
rect 24032 10004 24084 10056
rect 25044 10004 25096 10056
rect 34060 10072 34112 10124
rect 27804 10047 27856 10056
rect 20720 9936 20772 9988
rect 16488 9868 16540 9920
rect 16580 9868 16632 9920
rect 17316 9868 17368 9920
rect 22192 9868 22244 9920
rect 24676 9868 24728 9920
rect 27804 10013 27813 10047
rect 27813 10013 27847 10047
rect 27847 10013 27856 10047
rect 27804 10004 27856 10013
rect 29644 10004 29696 10056
rect 32312 10004 32364 10056
rect 32404 10004 32456 10056
rect 28908 9936 28960 9988
rect 29092 9979 29144 9988
rect 29092 9945 29101 9979
rect 29101 9945 29135 9979
rect 29135 9945 29144 9979
rect 30288 9979 30340 9988
rect 29092 9936 29144 9945
rect 30288 9945 30297 9979
rect 30297 9945 30331 9979
rect 30331 9945 30340 9979
rect 30288 9936 30340 9945
rect 35716 9936 35768 9988
rect 27252 9868 27304 9920
rect 30656 9868 30708 9920
rect 34980 9911 35032 9920
rect 34980 9877 34989 9911
rect 34989 9877 35023 9911
rect 35023 9877 35032 9911
rect 34980 9868 35032 9877
rect 35440 9911 35492 9920
rect 35440 9877 35449 9911
rect 35449 9877 35483 9911
rect 35483 9877 35492 9911
rect 35440 9868 35492 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4068 9596 4120 9648
rect 10968 9596 11020 9648
rect 13084 9596 13136 9648
rect 13452 9596 13504 9648
rect 14188 9528 14240 9580
rect 16120 9664 16172 9716
rect 16580 9596 16632 9648
rect 17040 9639 17092 9648
rect 17040 9605 17049 9639
rect 17049 9605 17083 9639
rect 17083 9605 17092 9639
rect 17040 9596 17092 9605
rect 17592 9664 17644 9716
rect 21548 9664 21600 9716
rect 24952 9664 25004 9716
rect 17960 9596 18012 9648
rect 18052 9596 18104 9648
rect 19984 9639 20036 9648
rect 19984 9605 19993 9639
rect 19993 9605 20027 9639
rect 20027 9605 20036 9639
rect 19984 9596 20036 9605
rect 20444 9596 20496 9648
rect 21916 9596 21968 9648
rect 23848 9596 23900 9648
rect 24216 9596 24268 9648
rect 14924 9571 14976 9580
rect 14924 9537 14933 9571
rect 14933 9537 14967 9571
rect 14967 9537 14976 9571
rect 14924 9528 14976 9537
rect 16304 9571 16356 9580
rect 16304 9537 16313 9571
rect 16313 9537 16347 9571
rect 16347 9537 16356 9571
rect 16304 9528 16356 9537
rect 24124 9528 24176 9580
rect 25044 9596 25096 9648
rect 27436 9596 27488 9648
rect 15476 9460 15528 9512
rect 17132 9460 17184 9512
rect 17408 9460 17460 9512
rect 17592 9503 17644 9512
rect 17592 9469 17601 9503
rect 17601 9469 17635 9503
rect 17635 9469 17644 9503
rect 17592 9460 17644 9469
rect 19156 9503 19208 9512
rect 16672 9392 16724 9444
rect 16764 9392 16816 9444
rect 18052 9392 18104 9444
rect 19156 9469 19165 9503
rect 19165 9469 19199 9503
rect 19199 9469 19208 9503
rect 19156 9460 19208 9469
rect 20720 9460 20772 9512
rect 20996 9460 21048 9512
rect 22008 9503 22060 9512
rect 22008 9469 22017 9503
rect 22017 9469 22051 9503
rect 22051 9469 22060 9503
rect 22008 9460 22060 9469
rect 22284 9460 22336 9512
rect 28724 9664 28776 9716
rect 30564 9664 30616 9716
rect 32496 9664 32548 9716
rect 37280 9664 37332 9716
rect 32956 9596 33008 9648
rect 36268 9639 36320 9648
rect 36268 9605 36277 9639
rect 36277 9605 36311 9639
rect 36311 9605 36320 9639
rect 36268 9596 36320 9605
rect 36912 9596 36964 9648
rect 24308 9460 24360 9512
rect 25320 9460 25372 9512
rect 26516 9503 26568 9512
rect 26516 9469 26525 9503
rect 26525 9469 26559 9503
rect 26559 9469 26568 9503
rect 26516 9460 26568 9469
rect 19248 9392 19300 9444
rect 17868 9324 17920 9376
rect 19708 9324 19760 9376
rect 22100 9324 22152 9376
rect 24032 9324 24084 9376
rect 25228 9324 25280 9376
rect 32772 9392 32824 9444
rect 37280 9460 37332 9512
rect 37924 9460 37976 9512
rect 34980 9392 35032 9444
rect 35348 9392 35400 9444
rect 29736 9324 29788 9376
rect 30196 9367 30248 9376
rect 30196 9333 30205 9367
rect 30205 9333 30239 9367
rect 30239 9333 30248 9367
rect 30196 9324 30248 9333
rect 30288 9324 30340 9376
rect 30840 9324 30892 9376
rect 31116 9324 31168 9376
rect 32864 9367 32916 9376
rect 32864 9333 32873 9367
rect 32873 9333 32907 9367
rect 32907 9333 32916 9367
rect 32864 9324 32916 9333
rect 35716 9367 35768 9376
rect 35716 9333 35725 9367
rect 35725 9333 35759 9367
rect 35759 9333 35768 9367
rect 35716 9324 35768 9333
rect 37648 9324 37700 9376
rect 38200 9367 38252 9376
rect 38200 9333 38209 9367
rect 38209 9333 38243 9367
rect 38243 9333 38252 9367
rect 38200 9324 38252 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 17040 9120 17092 9172
rect 17132 9120 17184 9172
rect 1860 9095 1912 9104
rect 1860 9061 1869 9095
rect 1869 9061 1903 9095
rect 1903 9061 1912 9095
rect 1860 9052 1912 9061
rect 13544 8916 13596 8968
rect 14280 8959 14332 8968
rect 14280 8925 14289 8959
rect 14289 8925 14323 8959
rect 14323 8925 14332 8959
rect 14280 8916 14332 8925
rect 14924 8959 14976 8968
rect 14924 8925 14933 8959
rect 14933 8925 14967 8959
rect 14967 8925 14976 8959
rect 16856 9052 16908 9104
rect 18512 9052 18564 9104
rect 18604 9052 18656 9104
rect 20536 9052 20588 9104
rect 23664 9120 23716 9172
rect 24676 9163 24728 9172
rect 24676 9129 24685 9163
rect 24685 9129 24719 9163
rect 24719 9129 24728 9163
rect 24676 9120 24728 9129
rect 24768 9120 24820 9172
rect 26148 9163 26200 9172
rect 26148 9129 26172 9163
rect 26172 9129 26200 9163
rect 26148 9120 26200 9129
rect 26792 9120 26844 9172
rect 24216 9052 24268 9104
rect 27252 9052 27304 9104
rect 30288 9052 30340 9104
rect 15936 8984 15988 9036
rect 17500 8984 17552 9036
rect 21732 8984 21784 9036
rect 22192 8984 22244 9036
rect 14924 8916 14976 8925
rect 16672 8916 16724 8968
rect 17776 8916 17828 8968
rect 20904 8959 20956 8968
rect 20904 8925 20913 8959
rect 20913 8925 20947 8959
rect 20947 8925 20956 8959
rect 20904 8916 20956 8925
rect 23112 8984 23164 9036
rect 23664 8984 23716 9036
rect 23388 8959 23440 8968
rect 23388 8925 23397 8959
rect 23397 8925 23431 8959
rect 23431 8925 23440 8959
rect 23388 8916 23440 8925
rect 24768 8959 24820 8968
rect 24768 8925 24777 8959
rect 24777 8925 24811 8959
rect 24811 8925 24820 8959
rect 24768 8916 24820 8925
rect 25044 8984 25096 9036
rect 25320 8916 25372 8968
rect 25688 8916 25740 8968
rect 26240 8984 26292 9036
rect 29460 8984 29512 9036
rect 36268 9120 36320 9172
rect 31024 8984 31076 9036
rect 27988 8916 28040 8968
rect 32864 8916 32916 8968
rect 1676 8891 1728 8900
rect 1676 8857 1685 8891
rect 1685 8857 1719 8891
rect 1719 8857 1728 8891
rect 1676 8848 1728 8857
rect 14372 8823 14424 8832
rect 14372 8789 14381 8823
rect 14381 8789 14415 8823
rect 14415 8789 14424 8823
rect 14372 8780 14424 8789
rect 15108 8780 15160 8832
rect 15936 8848 15988 8900
rect 17224 8848 17276 8900
rect 15844 8780 15896 8832
rect 18512 8848 18564 8900
rect 18696 8891 18748 8900
rect 18696 8857 18705 8891
rect 18705 8857 18739 8891
rect 18739 8857 18748 8891
rect 18696 8848 18748 8857
rect 18788 8891 18840 8900
rect 18788 8857 18797 8891
rect 18797 8857 18831 8891
rect 18831 8857 18840 8891
rect 18788 8848 18840 8857
rect 19156 8848 19208 8900
rect 19708 8848 19760 8900
rect 23940 8848 23992 8900
rect 24400 8848 24452 8900
rect 26424 8848 26476 8900
rect 27528 8848 27580 8900
rect 31024 8848 31076 8900
rect 31944 8848 31996 8900
rect 23664 8780 23716 8832
rect 23756 8780 23808 8832
rect 26516 8780 26568 8832
rect 27160 8780 27212 8832
rect 29092 8780 29144 8832
rect 29828 8780 29880 8832
rect 34796 8848 34848 8900
rect 35348 8848 35400 8900
rect 32864 8823 32916 8832
rect 32864 8789 32873 8823
rect 32873 8789 32907 8823
rect 32907 8789 32916 8823
rect 32864 8780 32916 8789
rect 34428 8780 34480 8832
rect 35716 8780 35768 8832
rect 37280 8780 37332 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 1676 8619 1728 8628
rect 1676 8585 1685 8619
rect 1685 8585 1719 8619
rect 1719 8585 1728 8619
rect 1676 8576 1728 8585
rect 14096 8551 14148 8560
rect 14096 8517 14105 8551
rect 14105 8517 14139 8551
rect 14139 8517 14148 8551
rect 14096 8508 14148 8517
rect 14372 8576 14424 8628
rect 14556 8508 14608 8560
rect 15752 8508 15804 8560
rect 16580 8508 16632 8560
rect 2504 8440 2556 8492
rect 14556 8372 14608 8424
rect 15844 8372 15896 8424
rect 17408 8576 17460 8628
rect 18604 8576 18656 8628
rect 18696 8576 18748 8628
rect 19432 8576 19484 8628
rect 19892 8576 19944 8628
rect 22008 8576 22060 8628
rect 17040 8551 17092 8560
rect 17040 8517 17049 8551
rect 17049 8517 17083 8551
rect 17083 8517 17092 8551
rect 17040 8508 17092 8517
rect 17592 8508 17644 8560
rect 18512 8508 18564 8560
rect 20904 8508 20956 8560
rect 19248 8440 19300 8492
rect 31208 8576 31260 8628
rect 32772 8576 32824 8628
rect 25688 8508 25740 8560
rect 27528 8508 27580 8560
rect 29828 8508 29880 8560
rect 30104 8508 30156 8560
rect 30840 8508 30892 8560
rect 31944 8508 31996 8560
rect 32220 8508 32272 8560
rect 24860 8440 24912 8492
rect 14096 8304 14148 8356
rect 17500 8347 17552 8356
rect 17500 8313 17509 8347
rect 17509 8313 17543 8347
rect 17543 8313 17552 8347
rect 17500 8304 17552 8313
rect 20720 8372 20772 8424
rect 21180 8415 21232 8424
rect 21180 8381 21189 8415
rect 21189 8381 21223 8415
rect 21223 8381 21232 8415
rect 21180 8372 21232 8381
rect 21456 8415 21508 8424
rect 21456 8381 21465 8415
rect 21465 8381 21499 8415
rect 21499 8381 21508 8415
rect 21456 8372 21508 8381
rect 22008 8372 22060 8424
rect 24032 8372 24084 8424
rect 25228 8372 25280 8424
rect 25320 8372 25372 8424
rect 26240 8415 26292 8424
rect 26240 8381 26249 8415
rect 26249 8381 26283 8415
rect 26283 8381 26292 8415
rect 26240 8372 26292 8381
rect 27160 8415 27212 8424
rect 27160 8381 27169 8415
rect 27169 8381 27203 8415
rect 27203 8381 27212 8415
rect 27160 8372 27212 8381
rect 15200 8236 15252 8288
rect 16396 8236 16448 8288
rect 16672 8236 16724 8288
rect 18604 8304 18656 8356
rect 20168 8304 20220 8356
rect 21824 8304 21876 8356
rect 22100 8304 22152 8356
rect 26424 8304 26476 8356
rect 27068 8304 27120 8356
rect 27528 8372 27580 8424
rect 29276 8372 29328 8424
rect 32864 8440 32916 8492
rect 35716 8483 35768 8492
rect 35716 8449 35725 8483
rect 35725 8449 35759 8483
rect 35759 8449 35768 8483
rect 35716 8440 35768 8449
rect 38292 8483 38344 8492
rect 38292 8449 38301 8483
rect 38301 8449 38335 8483
rect 38335 8449 38344 8483
rect 38292 8440 38344 8449
rect 30656 8372 30708 8424
rect 31024 8372 31076 8424
rect 18880 8236 18932 8288
rect 30104 8304 30156 8356
rect 29920 8236 29972 8288
rect 35348 8304 35400 8356
rect 32864 8236 32916 8288
rect 34612 8236 34664 8288
rect 37280 8236 37332 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 17040 8032 17092 8084
rect 17592 8032 17644 8084
rect 18328 8032 18380 8084
rect 19340 8032 19392 8084
rect 21640 8032 21692 8084
rect 16672 7964 16724 8016
rect 17224 7964 17276 8016
rect 14648 7939 14700 7948
rect 14648 7905 14657 7939
rect 14657 7905 14691 7939
rect 14691 7905 14700 7939
rect 14648 7896 14700 7905
rect 15016 7896 15068 7948
rect 17960 7964 18012 8016
rect 18696 7964 18748 8016
rect 20812 7964 20864 8016
rect 16948 7871 17000 7880
rect 16948 7837 16957 7871
rect 16957 7837 16991 7871
rect 16991 7837 17000 7871
rect 16948 7828 17000 7837
rect 21364 7896 21416 7948
rect 28632 7964 28684 8016
rect 29736 8007 29788 8016
rect 29736 7973 29745 8007
rect 29745 7973 29779 8007
rect 29779 7973 29788 8007
rect 29736 7964 29788 7973
rect 30564 7964 30616 8016
rect 18696 7871 18748 7880
rect 18144 7760 18196 7812
rect 18696 7837 18705 7871
rect 18705 7837 18739 7871
rect 18739 7837 18748 7871
rect 18696 7828 18748 7837
rect 19340 7828 19392 7880
rect 19984 7828 20036 7880
rect 20628 7828 20680 7880
rect 24584 7871 24636 7880
rect 24584 7837 24593 7871
rect 24593 7837 24627 7871
rect 24627 7837 24636 7871
rect 24584 7828 24636 7837
rect 30380 7896 30432 7948
rect 31668 8032 31720 8084
rect 34612 8032 34664 8084
rect 36268 8032 36320 8084
rect 37188 8032 37240 8084
rect 27160 7871 27212 7880
rect 27160 7837 27169 7871
rect 27169 7837 27203 7871
rect 27203 7837 27212 7871
rect 27160 7828 27212 7837
rect 30288 7828 30340 7880
rect 20812 7760 20864 7812
rect 20904 7760 20956 7812
rect 22468 7760 22520 7812
rect 23112 7760 23164 7812
rect 23572 7760 23624 7812
rect 24768 7760 24820 7812
rect 35624 7828 35676 7880
rect 15476 7692 15528 7744
rect 18052 7692 18104 7744
rect 20260 7692 20312 7744
rect 23204 7692 23256 7744
rect 23388 7692 23440 7744
rect 24308 7692 24360 7744
rect 27252 7692 27304 7744
rect 27620 7692 27672 7744
rect 29000 7692 29052 7744
rect 30380 7692 30432 7744
rect 33048 7760 33100 7812
rect 33784 7692 33836 7744
rect 37280 7692 37332 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 13636 7488 13688 7540
rect 15016 7531 15068 7540
rect 15016 7497 15025 7531
rect 15025 7497 15059 7531
rect 15059 7497 15068 7531
rect 15016 7488 15068 7497
rect 14188 7420 14240 7472
rect 2504 7395 2556 7404
rect 2504 7361 2513 7395
rect 2513 7361 2547 7395
rect 2547 7361 2556 7395
rect 2504 7352 2556 7361
rect 10048 7352 10100 7404
rect 17224 7420 17276 7472
rect 17408 7463 17460 7472
rect 17408 7429 17417 7463
rect 17417 7429 17451 7463
rect 17451 7429 17460 7463
rect 17408 7420 17460 7429
rect 17960 7488 18012 7540
rect 18328 7488 18380 7540
rect 18788 7488 18840 7540
rect 19156 7531 19208 7540
rect 19156 7497 19165 7531
rect 19165 7497 19199 7531
rect 19199 7497 19208 7531
rect 19156 7488 19208 7497
rect 19248 7420 19300 7472
rect 16764 7352 16816 7404
rect 19064 7395 19116 7404
rect 19064 7361 19073 7395
rect 19073 7361 19107 7395
rect 19107 7361 19116 7395
rect 19064 7352 19116 7361
rect 16672 7284 16724 7336
rect 22192 7420 22244 7472
rect 22928 7488 22980 7540
rect 24952 7420 25004 7472
rect 25964 7463 26016 7472
rect 25964 7429 25973 7463
rect 25973 7429 26007 7463
rect 26007 7429 26016 7463
rect 25964 7420 26016 7429
rect 27068 7488 27120 7540
rect 27344 7420 27396 7472
rect 29552 7488 29604 7540
rect 29828 7488 29880 7540
rect 31116 7488 31168 7540
rect 31668 7488 31720 7540
rect 35716 7531 35768 7540
rect 35716 7497 35725 7531
rect 35725 7497 35759 7531
rect 35759 7497 35768 7531
rect 35716 7488 35768 7497
rect 37188 7488 37240 7540
rect 32956 7420 33008 7472
rect 20076 7352 20128 7404
rect 21456 7395 21508 7404
rect 21456 7361 21465 7395
rect 21465 7361 21499 7395
rect 21499 7361 21508 7395
rect 21456 7352 21508 7361
rect 21640 7352 21692 7404
rect 26240 7395 26292 7404
rect 26240 7361 26249 7395
rect 26249 7361 26283 7395
rect 26283 7361 26292 7395
rect 26240 7352 26292 7361
rect 20628 7284 20680 7336
rect 22376 7284 22428 7336
rect 25872 7284 25924 7336
rect 26332 7284 26384 7336
rect 26700 7284 26752 7336
rect 27160 7327 27212 7336
rect 27160 7293 27169 7327
rect 27169 7293 27203 7327
rect 27203 7293 27212 7327
rect 27160 7284 27212 7293
rect 29000 7352 29052 7404
rect 30012 7352 30064 7404
rect 37280 7352 37332 7404
rect 17132 7216 17184 7268
rect 17316 7216 17368 7268
rect 31024 7284 31076 7336
rect 1676 7191 1728 7200
rect 1676 7157 1685 7191
rect 1685 7157 1719 7191
rect 1719 7157 1728 7191
rect 1676 7148 1728 7157
rect 15568 7148 15620 7200
rect 18788 7148 18840 7200
rect 19984 7148 20036 7200
rect 28632 7216 28684 7268
rect 28908 7216 28960 7268
rect 30196 7216 30248 7268
rect 21916 7148 21968 7200
rect 22100 7148 22152 7200
rect 22652 7148 22704 7200
rect 23388 7148 23440 7200
rect 25228 7148 25280 7200
rect 29276 7148 29328 7200
rect 29736 7148 29788 7200
rect 30288 7148 30340 7200
rect 31668 7191 31720 7200
rect 31668 7157 31677 7191
rect 31677 7157 31711 7191
rect 31711 7157 31720 7191
rect 31668 7148 31720 7157
rect 32864 7191 32916 7200
rect 32864 7157 32873 7191
rect 32873 7157 32907 7191
rect 32907 7157 32916 7191
rect 32864 7148 32916 7157
rect 38016 7191 38068 7200
rect 38016 7157 38025 7191
rect 38025 7157 38059 7191
rect 38059 7157 38068 7191
rect 38016 7148 38068 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 15292 6851 15344 6860
rect 15292 6817 15301 6851
rect 15301 6817 15335 6851
rect 15335 6817 15344 6851
rect 15292 6808 15344 6817
rect 15752 6808 15804 6860
rect 6368 6783 6420 6792
rect 6368 6749 6377 6783
rect 6377 6749 6411 6783
rect 6411 6749 6420 6783
rect 17316 6876 17368 6928
rect 18236 6876 18288 6928
rect 16580 6851 16632 6860
rect 16580 6817 16589 6851
rect 16589 6817 16623 6851
rect 16623 6817 16632 6851
rect 16580 6808 16632 6817
rect 18420 6851 18472 6860
rect 6368 6740 6420 6749
rect 18144 6740 18196 6792
rect 18420 6817 18429 6851
rect 18429 6817 18463 6851
rect 18463 6817 18472 6851
rect 18420 6808 18472 6817
rect 18788 6944 18840 6996
rect 23296 6944 23348 6996
rect 26056 6944 26108 6996
rect 29000 6944 29052 6996
rect 29552 6944 29604 6996
rect 30748 6944 30800 6996
rect 31760 6944 31812 6996
rect 33692 6944 33744 6996
rect 19156 6876 19208 6928
rect 20076 6876 20128 6928
rect 22376 6876 22428 6928
rect 25136 6876 25188 6928
rect 31208 6876 31260 6928
rect 33324 6876 33376 6928
rect 14648 6715 14700 6724
rect 14648 6681 14657 6715
rect 14657 6681 14691 6715
rect 14691 6681 14700 6715
rect 14648 6672 14700 6681
rect 15844 6672 15896 6724
rect 16488 6672 16540 6724
rect 17776 6715 17828 6724
rect 17776 6681 17785 6715
rect 17785 6681 17819 6715
rect 17819 6681 17828 6715
rect 17776 6672 17828 6681
rect 6552 6647 6604 6656
rect 6552 6613 6561 6647
rect 6561 6613 6595 6647
rect 6595 6613 6604 6647
rect 6552 6604 6604 6613
rect 18788 6740 18840 6792
rect 19432 6808 19484 6860
rect 19248 6740 19300 6792
rect 20260 6808 20312 6860
rect 21732 6808 21784 6860
rect 22560 6808 22612 6860
rect 24400 6808 24452 6860
rect 26148 6808 26200 6860
rect 27344 6808 27396 6860
rect 30564 6808 30616 6860
rect 19708 6740 19760 6792
rect 22468 6740 22520 6792
rect 27160 6740 27212 6792
rect 29000 6783 29052 6792
rect 29000 6749 29009 6783
rect 29009 6749 29043 6783
rect 29043 6749 29052 6783
rect 29736 6783 29788 6792
rect 29000 6740 29052 6749
rect 29736 6749 29745 6783
rect 29745 6749 29779 6783
rect 29779 6749 29788 6783
rect 29736 6740 29788 6749
rect 33048 6740 33100 6792
rect 33508 6783 33560 6792
rect 33508 6749 33517 6783
rect 33517 6749 33551 6783
rect 33551 6749 33560 6783
rect 34060 6783 34112 6792
rect 33508 6740 33560 6749
rect 34060 6749 34069 6783
rect 34069 6749 34103 6783
rect 34103 6749 34112 6783
rect 34060 6740 34112 6749
rect 34888 6740 34940 6792
rect 35532 6740 35584 6792
rect 37280 6740 37332 6792
rect 20720 6604 20772 6656
rect 21916 6604 21968 6656
rect 22192 6672 22244 6724
rect 26240 6715 26292 6724
rect 26240 6681 26249 6715
rect 26249 6681 26283 6715
rect 26283 6681 26292 6715
rect 26240 6672 26292 6681
rect 22376 6604 22428 6656
rect 22744 6604 22796 6656
rect 24308 6604 24360 6656
rect 24860 6604 24912 6656
rect 30288 6672 30340 6724
rect 31668 6672 31720 6724
rect 35348 6672 35400 6724
rect 26424 6604 26476 6656
rect 27988 6604 28040 6656
rect 28816 6604 28868 6656
rect 28908 6604 28960 6656
rect 29552 6604 29604 6656
rect 30932 6604 30984 6656
rect 31024 6604 31076 6656
rect 34520 6604 34572 6656
rect 36636 6604 36688 6656
rect 38016 6604 38068 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 15476 6400 15528 6452
rect 18696 6400 18748 6452
rect 19984 6400 20036 6452
rect 24216 6443 24268 6452
rect 9772 6332 9824 6384
rect 13820 6332 13872 6384
rect 19432 6332 19484 6384
rect 21732 6332 21784 6384
rect 24216 6409 24225 6443
rect 24225 6409 24259 6443
rect 24259 6409 24268 6443
rect 24216 6400 24268 6409
rect 24308 6400 24360 6452
rect 26608 6400 26660 6452
rect 23204 6332 23256 6384
rect 25228 6332 25280 6384
rect 26424 6332 26476 6384
rect 26884 6332 26936 6384
rect 28356 6400 28408 6452
rect 29000 6400 29052 6452
rect 29736 6400 29788 6452
rect 27068 6332 27120 6384
rect 28724 6332 28776 6384
rect 29092 6332 29144 6384
rect 30564 6400 30616 6452
rect 32680 6443 32732 6452
rect 30288 6332 30340 6384
rect 19524 6264 19576 6316
rect 21640 6264 21692 6316
rect 22468 6307 22520 6316
rect 22468 6273 22477 6307
rect 22477 6273 22511 6307
rect 22511 6273 22520 6307
rect 22468 6264 22520 6273
rect 26056 6264 26108 6316
rect 26608 6264 26660 6316
rect 29276 6264 29328 6316
rect 32680 6409 32689 6443
rect 32689 6409 32723 6443
rect 32723 6409 32732 6443
rect 32680 6400 32732 6409
rect 33324 6443 33376 6452
rect 33324 6409 33333 6443
rect 33333 6409 33367 6443
rect 33367 6409 33376 6443
rect 33324 6400 33376 6409
rect 33508 6400 33560 6452
rect 34612 6443 34664 6452
rect 34612 6409 34621 6443
rect 34621 6409 34655 6443
rect 34655 6409 34664 6443
rect 34612 6400 34664 6409
rect 34796 6400 34848 6452
rect 36544 6400 36596 6452
rect 34428 6332 34480 6384
rect 31116 6264 31168 6316
rect 17040 6196 17092 6248
rect 19616 6196 19668 6248
rect 19984 6239 20036 6248
rect 16948 6128 17000 6180
rect 19432 6128 19484 6180
rect 14464 6060 14516 6112
rect 16120 6060 16172 6112
rect 17776 6060 17828 6112
rect 19248 6060 19300 6112
rect 19340 6060 19392 6112
rect 19616 6060 19668 6112
rect 19984 6205 19993 6239
rect 19993 6205 20027 6239
rect 20027 6205 20036 6239
rect 19984 6196 20036 6205
rect 24584 6196 24636 6248
rect 20996 6128 21048 6180
rect 21548 6128 21600 6180
rect 22192 6128 22244 6180
rect 23940 6128 23992 6180
rect 29828 6196 29880 6248
rect 30196 6196 30248 6248
rect 33140 6264 33192 6316
rect 34612 6264 34664 6316
rect 35624 6332 35676 6384
rect 36636 6264 36688 6316
rect 37556 6264 37608 6316
rect 38200 6264 38252 6316
rect 36268 6196 36320 6248
rect 27160 6171 27212 6180
rect 21640 6060 21692 6112
rect 21824 6060 21876 6112
rect 23756 6060 23808 6112
rect 24584 6060 24636 6112
rect 27160 6137 27169 6171
rect 27169 6137 27203 6171
rect 27203 6137 27212 6171
rect 27160 6128 27212 6137
rect 28356 6128 28408 6180
rect 26424 6103 26476 6112
rect 26424 6069 26433 6103
rect 26433 6069 26467 6103
rect 26467 6069 26476 6103
rect 26424 6060 26476 6069
rect 26516 6060 26568 6112
rect 34244 6128 34296 6180
rect 34612 6128 34664 6180
rect 35532 6128 35584 6180
rect 30932 6060 30984 6112
rect 32588 6060 32640 6112
rect 32956 6060 33008 6112
rect 34796 6060 34848 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 14832 5856 14884 5908
rect 17408 5856 17460 5908
rect 19064 5856 19116 5908
rect 19248 5856 19300 5908
rect 20904 5856 20956 5908
rect 21180 5856 21232 5908
rect 21548 5856 21600 5908
rect 22100 5856 22152 5908
rect 23664 5856 23716 5908
rect 23756 5899 23808 5908
rect 23756 5865 23765 5899
rect 23765 5865 23799 5899
rect 23799 5865 23808 5899
rect 23756 5856 23808 5865
rect 25964 5856 26016 5908
rect 26056 5856 26108 5908
rect 17224 5788 17276 5840
rect 14648 5720 14700 5772
rect 16028 5763 16080 5772
rect 16028 5729 16037 5763
rect 16037 5729 16071 5763
rect 16071 5729 16080 5763
rect 16028 5720 16080 5729
rect 16304 5720 16356 5772
rect 23296 5788 23348 5840
rect 24768 5788 24820 5840
rect 19340 5720 19392 5772
rect 13452 5652 13504 5704
rect 14464 5695 14516 5704
rect 14464 5661 14473 5695
rect 14473 5661 14507 5695
rect 14507 5661 14516 5695
rect 14464 5652 14516 5661
rect 15936 5627 15988 5636
rect 15936 5593 15945 5627
rect 15945 5593 15979 5627
rect 15979 5593 15988 5627
rect 15936 5584 15988 5593
rect 20168 5652 20220 5704
rect 20260 5695 20312 5704
rect 20260 5661 20269 5695
rect 20269 5661 20303 5695
rect 20303 5661 20312 5695
rect 20260 5652 20312 5661
rect 20628 5652 20680 5704
rect 21456 5695 21508 5704
rect 21456 5661 21465 5695
rect 21465 5661 21499 5695
rect 21499 5661 21508 5695
rect 21456 5652 21508 5661
rect 26424 5720 26476 5772
rect 27528 5720 27580 5772
rect 19064 5584 19116 5636
rect 20904 5584 20956 5636
rect 2780 5559 2832 5568
rect 2780 5525 2789 5559
rect 2789 5525 2823 5559
rect 2823 5525 2832 5559
rect 2780 5516 2832 5525
rect 13084 5516 13136 5568
rect 16672 5516 16724 5568
rect 18604 5516 18656 5568
rect 19616 5516 19668 5568
rect 19984 5516 20036 5568
rect 26332 5695 26384 5704
rect 26332 5661 26341 5695
rect 26341 5661 26375 5695
rect 26375 5661 26384 5695
rect 26332 5652 26384 5661
rect 27160 5652 27212 5704
rect 29644 5788 29696 5840
rect 30196 5788 30248 5840
rect 31484 5856 31536 5908
rect 33324 5856 33376 5908
rect 28908 5763 28960 5772
rect 28908 5729 28917 5763
rect 28917 5729 28951 5763
rect 28951 5729 28960 5763
rect 28908 5720 28960 5729
rect 30656 5720 30708 5772
rect 31668 5720 31720 5772
rect 32588 5720 32640 5772
rect 32956 5695 33008 5704
rect 26056 5627 26108 5636
rect 21824 5516 21876 5568
rect 23848 5516 23900 5568
rect 24308 5516 24360 5568
rect 24584 5559 24636 5568
rect 24584 5525 24593 5559
rect 24593 5525 24627 5559
rect 24627 5525 24636 5559
rect 24584 5516 24636 5525
rect 26056 5593 26065 5627
rect 26065 5593 26099 5627
rect 26099 5593 26108 5627
rect 26056 5584 26108 5593
rect 29000 5584 29052 5636
rect 32956 5661 32965 5695
rect 32965 5661 32999 5695
rect 32999 5661 33008 5695
rect 32956 5652 33008 5661
rect 33140 5652 33192 5704
rect 34152 5695 34204 5704
rect 34152 5661 34161 5695
rect 34161 5661 34195 5695
rect 34195 5661 34204 5695
rect 34152 5652 34204 5661
rect 35072 5695 35124 5704
rect 35072 5661 35081 5695
rect 35081 5661 35115 5695
rect 35115 5661 35124 5695
rect 35072 5652 35124 5661
rect 35808 5652 35860 5704
rect 36268 5652 36320 5704
rect 37280 5652 37332 5704
rect 38016 5652 38068 5704
rect 29920 5584 29972 5636
rect 32496 5516 32548 5568
rect 37280 5516 37332 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 1860 5219 1912 5228
rect 1860 5185 1869 5219
rect 1869 5185 1903 5219
rect 1903 5185 1912 5219
rect 1860 5176 1912 5185
rect 13544 5312 13596 5364
rect 15016 5355 15068 5364
rect 15016 5321 15025 5355
rect 15025 5321 15059 5355
rect 15059 5321 15068 5355
rect 15016 5312 15068 5321
rect 13084 5287 13136 5296
rect 13084 5253 13093 5287
rect 13093 5253 13127 5287
rect 13127 5253 13136 5287
rect 13084 5244 13136 5253
rect 16580 5312 16632 5364
rect 16764 5312 16816 5364
rect 11888 5219 11940 5228
rect 11888 5185 11897 5219
rect 11897 5185 11931 5219
rect 11931 5185 11940 5219
rect 11888 5176 11940 5185
rect 13452 5176 13504 5228
rect 13912 5176 13964 5228
rect 14464 5176 14516 5228
rect 14924 5219 14976 5228
rect 14924 5185 14933 5219
rect 14933 5185 14967 5219
rect 14967 5185 14976 5219
rect 14924 5176 14976 5185
rect 15844 5219 15896 5228
rect 15844 5185 15853 5219
rect 15853 5185 15887 5219
rect 15887 5185 15896 5219
rect 15844 5176 15896 5185
rect 17040 5219 17092 5228
rect 17040 5185 17049 5219
rect 17049 5185 17083 5219
rect 17083 5185 17092 5219
rect 17040 5176 17092 5185
rect 17408 5244 17460 5296
rect 21456 5312 21508 5364
rect 22468 5312 22520 5364
rect 19892 5176 19944 5228
rect 21456 5219 21508 5228
rect 21456 5185 21465 5219
rect 21465 5185 21499 5219
rect 21499 5185 21508 5219
rect 22192 5244 22244 5296
rect 29644 5312 29696 5364
rect 23112 5287 23164 5296
rect 23112 5253 23121 5287
rect 23121 5253 23155 5287
rect 23155 5253 23164 5287
rect 23112 5244 23164 5253
rect 24032 5244 24084 5296
rect 24400 5287 24452 5296
rect 24400 5253 24409 5287
rect 24409 5253 24443 5287
rect 24443 5253 24452 5287
rect 24400 5244 24452 5253
rect 25780 5244 25832 5296
rect 26516 5244 26568 5296
rect 29920 5312 29972 5364
rect 30288 5312 30340 5364
rect 32036 5244 32088 5296
rect 33784 5287 33836 5296
rect 33784 5253 33793 5287
rect 33793 5253 33827 5287
rect 33827 5253 33836 5287
rect 33784 5244 33836 5253
rect 37924 5244 37976 5296
rect 38108 5244 38160 5296
rect 21456 5176 21508 5185
rect 23204 5176 23256 5228
rect 24124 5219 24176 5228
rect 24124 5185 24133 5219
rect 24133 5185 24167 5219
rect 24167 5185 24176 5219
rect 24124 5176 24176 5185
rect 12440 5083 12492 5092
rect 12440 5049 12449 5083
rect 12449 5049 12483 5083
rect 12483 5049 12492 5083
rect 12440 5040 12492 5049
rect 1676 5015 1728 5024
rect 1676 4981 1685 5015
rect 1685 4981 1719 5015
rect 1719 4981 1728 5015
rect 1676 4972 1728 4981
rect 9772 5015 9824 5024
rect 9772 4981 9781 5015
rect 9781 4981 9815 5015
rect 9815 4981 9824 5015
rect 9772 4972 9824 4981
rect 16764 5108 16816 5160
rect 18328 5108 18380 5160
rect 19248 5108 19300 5160
rect 20812 5108 20864 5160
rect 21640 5108 21692 5160
rect 22192 5108 22244 5160
rect 14648 5040 14700 5092
rect 14372 5015 14424 5024
rect 14372 4981 14381 5015
rect 14381 4981 14415 5015
rect 14415 4981 14424 5015
rect 16856 5015 16908 5024
rect 14372 4972 14424 4981
rect 16856 4981 16865 5015
rect 16865 4981 16899 5015
rect 16899 4981 16908 5015
rect 16856 4972 16908 4981
rect 17776 4972 17828 5024
rect 18144 5015 18196 5024
rect 18144 4981 18153 5015
rect 18153 4981 18187 5015
rect 18187 4981 18196 5015
rect 18144 4972 18196 4981
rect 19248 5015 19300 5024
rect 19248 4981 19257 5015
rect 19257 4981 19291 5015
rect 19291 4981 19300 5015
rect 19248 4972 19300 4981
rect 19708 5015 19760 5024
rect 19708 4981 19717 5015
rect 19717 4981 19751 5015
rect 19751 4981 19760 5015
rect 19708 4972 19760 4981
rect 19892 5040 19944 5092
rect 20076 5040 20128 5092
rect 24952 5108 25004 5160
rect 25136 5108 25188 5160
rect 22192 4972 22244 5024
rect 22560 5040 22612 5092
rect 24032 5040 24084 5092
rect 22468 4972 22520 5024
rect 23020 4972 23072 5024
rect 26884 5176 26936 5228
rect 27988 5108 28040 5160
rect 30288 5176 30340 5228
rect 31300 5176 31352 5228
rect 34152 5176 34204 5228
rect 34336 5176 34388 5228
rect 34520 5176 34572 5228
rect 34796 5176 34848 5228
rect 35072 5176 35124 5228
rect 36268 5176 36320 5228
rect 29460 5108 29512 5160
rect 33692 5108 33744 5160
rect 34060 5151 34112 5160
rect 34060 5117 34069 5151
rect 34069 5117 34103 5151
rect 34103 5117 34112 5151
rect 34060 5108 34112 5117
rect 34428 5108 34480 5160
rect 34336 5040 34388 5092
rect 31576 4972 31628 5024
rect 32312 5015 32364 5024
rect 32312 4981 32321 5015
rect 32321 4981 32355 5015
rect 32355 4981 32364 5015
rect 32312 4972 32364 4981
rect 35900 5015 35952 5024
rect 35900 4981 35909 5015
rect 35909 4981 35943 5015
rect 35943 4981 35952 5015
rect 35900 4972 35952 4981
rect 36544 5015 36596 5024
rect 36544 4981 36553 5015
rect 36553 4981 36587 5015
rect 36587 4981 36596 5015
rect 36544 4972 36596 4981
rect 37556 5015 37608 5024
rect 37556 4981 37565 5015
rect 37565 4981 37599 5015
rect 37599 4981 37608 5015
rect 37556 4972 37608 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 12348 4811 12400 4820
rect 12348 4777 12357 4811
rect 12357 4777 12391 4811
rect 12391 4777 12400 4811
rect 12348 4768 12400 4777
rect 13820 4768 13872 4820
rect 14648 4811 14700 4820
rect 14648 4777 14657 4811
rect 14657 4777 14691 4811
rect 14691 4777 14700 4811
rect 14648 4768 14700 4777
rect 15936 4768 15988 4820
rect 16028 4768 16080 4820
rect 22836 4768 22888 4820
rect 23020 4768 23072 4820
rect 24124 4768 24176 4820
rect 24216 4768 24268 4820
rect 19340 4700 19392 4752
rect 19708 4700 19760 4752
rect 20352 4700 20404 4752
rect 22376 4743 22428 4752
rect 22376 4709 22385 4743
rect 22385 4709 22419 4743
rect 22419 4709 22428 4743
rect 22376 4700 22428 4709
rect 24676 4700 24728 4752
rect 24860 4768 24912 4820
rect 26424 4768 26476 4820
rect 26700 4768 26752 4820
rect 31300 4768 31352 4820
rect 31392 4768 31444 4820
rect 32220 4811 32272 4820
rect 32220 4777 32250 4811
rect 32250 4777 32272 4811
rect 32220 4768 32272 4777
rect 11796 4607 11848 4616
rect 11796 4573 11805 4607
rect 11805 4573 11839 4607
rect 11839 4573 11848 4607
rect 11796 4564 11848 4573
rect 13452 4564 13504 4616
rect 13912 4564 13964 4616
rect 14924 4564 14976 4616
rect 15292 4564 15344 4616
rect 20260 4632 20312 4684
rect 15844 4607 15896 4616
rect 15844 4573 15853 4607
rect 15853 4573 15887 4607
rect 15887 4573 15896 4607
rect 15844 4564 15896 4573
rect 16028 4496 16080 4548
rect 15936 4471 15988 4480
rect 15936 4437 15945 4471
rect 15945 4437 15979 4471
rect 15979 4437 15988 4471
rect 15936 4428 15988 4437
rect 16120 4428 16172 4480
rect 16672 4564 16724 4616
rect 17592 4564 17644 4616
rect 17224 4539 17276 4548
rect 17224 4505 17233 4539
rect 17233 4505 17267 4539
rect 17267 4505 17276 4539
rect 17224 4496 17276 4505
rect 19432 4564 19484 4616
rect 21456 4632 21508 4684
rect 23756 4632 23808 4684
rect 24492 4632 24544 4684
rect 24860 4632 24912 4684
rect 28264 4675 28316 4684
rect 28264 4641 28273 4675
rect 28273 4641 28307 4675
rect 28307 4641 28316 4675
rect 28264 4632 28316 4641
rect 29000 4632 29052 4684
rect 31300 4632 31352 4684
rect 33508 4700 33560 4752
rect 18604 4428 18656 4480
rect 19248 4428 19300 4480
rect 23020 4564 23072 4616
rect 26332 4607 26384 4616
rect 26332 4573 26341 4607
rect 26341 4573 26375 4607
rect 26375 4573 26384 4607
rect 26332 4564 26384 4573
rect 20260 4496 20312 4548
rect 20904 4539 20956 4548
rect 20904 4505 20913 4539
rect 20913 4505 20947 4539
rect 20947 4505 20956 4539
rect 20904 4496 20956 4505
rect 21640 4496 21692 4548
rect 20168 4428 20220 4480
rect 22836 4496 22888 4548
rect 23756 4428 23808 4480
rect 24676 4428 24728 4480
rect 28908 4496 28960 4548
rect 29000 4471 29052 4480
rect 29000 4437 29009 4471
rect 29009 4437 29043 4471
rect 29043 4437 29052 4471
rect 29000 4428 29052 4437
rect 29184 4496 29236 4548
rect 31668 4564 31720 4616
rect 35900 4632 35952 4684
rect 34152 4564 34204 4616
rect 34612 4564 34664 4616
rect 35808 4564 35860 4616
rect 36360 4607 36412 4616
rect 36360 4573 36369 4607
rect 36369 4573 36403 4607
rect 36403 4573 36412 4607
rect 36360 4564 36412 4573
rect 37648 4607 37700 4616
rect 37648 4573 37657 4607
rect 37657 4573 37691 4607
rect 37691 4573 37700 4607
rect 37648 4564 37700 4573
rect 38016 4564 38068 4616
rect 32496 4496 32548 4548
rect 33784 4428 33836 4480
rect 34980 4471 35032 4480
rect 34980 4437 34989 4471
rect 34989 4437 35023 4471
rect 35023 4437 35032 4471
rect 34980 4428 35032 4437
rect 35348 4428 35400 4480
rect 35992 4428 36044 4480
rect 37004 4428 37056 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 11612 4156 11664 4208
rect 15752 4224 15804 4276
rect 15936 4224 15988 4276
rect 24676 4224 24728 4276
rect 14280 4199 14332 4208
rect 14280 4165 14289 4199
rect 14289 4165 14323 4199
rect 14323 4165 14332 4199
rect 14280 4156 14332 4165
rect 13452 4131 13504 4140
rect 13452 4097 13461 4131
rect 13461 4097 13495 4131
rect 13495 4097 13504 4131
rect 13452 4088 13504 4097
rect 15292 4131 15344 4140
rect 15292 4097 15301 4131
rect 15301 4097 15335 4131
rect 15335 4097 15344 4131
rect 15292 4088 15344 4097
rect 15844 4088 15896 4140
rect 16120 4131 16172 4140
rect 16120 4097 16129 4131
rect 16129 4097 16163 4131
rect 16163 4097 16172 4131
rect 16120 4088 16172 4097
rect 17960 4156 18012 4208
rect 18604 4156 18656 4208
rect 17040 4131 17092 4140
rect 17040 4097 17049 4131
rect 17049 4097 17083 4131
rect 17083 4097 17092 4131
rect 17040 4088 17092 4097
rect 17316 4088 17368 4140
rect 17592 4131 17644 4140
rect 17592 4097 17609 4131
rect 17609 4097 17643 4131
rect 17643 4097 17644 4131
rect 17592 4088 17644 4097
rect 18512 4088 18564 4140
rect 18788 4088 18840 4140
rect 19248 4088 19300 4140
rect 21824 4156 21876 4208
rect 33876 4224 33928 4276
rect 24952 4156 25004 4208
rect 29552 4156 29604 4208
rect 31300 4156 31352 4208
rect 36544 4224 36596 4276
rect 34888 4156 34940 4208
rect 12532 4020 12584 4072
rect 14556 4063 14608 4072
rect 14556 4029 14565 4063
rect 14565 4029 14599 4063
rect 14599 4029 14608 4063
rect 14556 4020 14608 4029
rect 16304 4020 16356 4072
rect 16580 4020 16632 4072
rect 17408 4020 17460 4072
rect 17684 4063 17736 4072
rect 17684 4029 17693 4063
rect 17693 4029 17727 4063
rect 17727 4029 17736 4063
rect 17684 4020 17736 4029
rect 13636 3952 13688 4004
rect 18052 3884 18104 3936
rect 18604 3927 18656 3936
rect 18604 3893 18613 3927
rect 18613 3893 18647 3927
rect 18647 3893 18656 3927
rect 18604 3884 18656 3893
rect 22008 4131 22060 4140
rect 22008 4097 22017 4131
rect 22017 4097 22051 4131
rect 22051 4097 22060 4131
rect 22008 4088 22060 4097
rect 24216 4131 24268 4140
rect 24216 4097 24225 4131
rect 24225 4097 24259 4131
rect 24259 4097 24268 4131
rect 24216 4088 24268 4097
rect 26424 4131 26476 4140
rect 26424 4097 26433 4131
rect 26433 4097 26467 4131
rect 26467 4097 26476 4131
rect 26424 4088 26476 4097
rect 26516 4131 26568 4140
rect 26516 4097 26525 4131
rect 26525 4097 26559 4131
rect 26559 4097 26568 4131
rect 26516 4088 26568 4097
rect 20720 4020 20772 4072
rect 22376 4020 22428 4072
rect 24492 4063 24544 4072
rect 23664 3952 23716 4004
rect 24216 3952 24268 4004
rect 22100 3884 22152 3936
rect 22468 3884 22520 3936
rect 24032 3884 24084 3936
rect 24492 4029 24501 4063
rect 24501 4029 24535 4063
rect 24535 4029 24544 4063
rect 24492 4020 24544 4029
rect 26332 4020 26384 4072
rect 27436 4020 27488 4072
rect 29368 4020 29420 4072
rect 31484 4131 31536 4140
rect 31484 4097 31493 4131
rect 31493 4097 31527 4131
rect 31527 4097 31536 4131
rect 31484 4088 31536 4097
rect 31668 4088 31720 4140
rect 33876 4088 33928 4140
rect 34612 4088 34664 4140
rect 36360 4156 36412 4208
rect 34980 4088 35032 4140
rect 35440 4088 35492 4140
rect 35808 4088 35860 4140
rect 30748 4020 30800 4072
rect 30840 4020 30892 4072
rect 31116 4020 31168 4072
rect 32588 4063 32640 4072
rect 26148 3952 26200 4004
rect 26424 3952 26476 4004
rect 28816 3952 28868 4004
rect 25964 3927 26016 3936
rect 25964 3893 25973 3927
rect 25973 3893 26007 3927
rect 26007 3893 26016 3927
rect 25964 3884 26016 3893
rect 26700 3884 26752 3936
rect 29000 3884 29052 3936
rect 29276 3927 29328 3936
rect 29276 3893 29285 3927
rect 29285 3893 29319 3927
rect 29319 3893 29328 3927
rect 29276 3884 29328 3893
rect 32128 3952 32180 4004
rect 32588 4029 32597 4063
rect 32597 4029 32631 4063
rect 32631 4029 32640 4063
rect 32588 4020 32640 4029
rect 33140 4020 33192 4072
rect 34520 3952 34572 4004
rect 36636 3952 36688 4004
rect 37648 3952 37700 4004
rect 33784 3884 33836 3936
rect 33876 3884 33928 3936
rect 34152 3884 34204 3936
rect 34704 3884 34756 3936
rect 35900 3927 35952 3936
rect 35900 3893 35909 3927
rect 35909 3893 35943 3927
rect 35943 3893 35952 3927
rect 35900 3884 35952 3893
rect 36176 3884 36228 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2320 3723 2372 3732
rect 2320 3689 2329 3723
rect 2329 3689 2363 3723
rect 2363 3689 2372 3723
rect 2320 3680 2372 3689
rect 10968 3680 11020 3732
rect 11612 3723 11664 3732
rect 11612 3689 11621 3723
rect 11621 3689 11655 3723
rect 11655 3689 11664 3723
rect 11612 3680 11664 3689
rect 12256 3723 12308 3732
rect 12256 3689 12265 3723
rect 12265 3689 12299 3723
rect 12299 3689 12308 3723
rect 12256 3680 12308 3689
rect 14280 3680 14332 3732
rect 14188 3612 14240 3664
rect 2780 3476 2832 3528
rect 11796 3476 11848 3528
rect 12900 3544 12952 3596
rect 12992 3476 13044 3528
rect 13728 3476 13780 3528
rect 14280 3519 14332 3528
rect 14280 3485 14289 3519
rect 14289 3485 14323 3519
rect 14323 3485 14332 3519
rect 14280 3476 14332 3485
rect 17500 3544 17552 3596
rect 18604 3544 18656 3596
rect 19156 3544 19208 3596
rect 21548 3544 21600 3596
rect 22100 3680 22152 3732
rect 23020 3680 23072 3732
rect 23204 3723 23256 3732
rect 23204 3689 23213 3723
rect 23213 3689 23247 3723
rect 23247 3689 23256 3723
rect 23204 3680 23256 3689
rect 21916 3612 21968 3664
rect 22928 3544 22980 3596
rect 17132 3519 17184 3528
rect 17132 3485 17141 3519
rect 17141 3485 17175 3519
rect 17175 3485 17184 3519
rect 17132 3476 17184 3485
rect 17408 3476 17460 3528
rect 17868 3519 17920 3528
rect 17868 3485 17877 3519
rect 17877 3485 17911 3519
rect 17911 3485 17920 3519
rect 17868 3476 17920 3485
rect 18512 3519 18564 3528
rect 18512 3485 18521 3519
rect 18521 3485 18555 3519
rect 18555 3485 18564 3519
rect 18512 3476 18564 3485
rect 1676 3383 1728 3392
rect 1676 3349 1685 3383
rect 1685 3349 1719 3383
rect 1719 3349 1728 3383
rect 1676 3340 1728 3349
rect 16948 3408 17000 3460
rect 18144 3408 18196 3460
rect 18696 3408 18748 3460
rect 12992 3340 13044 3392
rect 16764 3340 16816 3392
rect 18880 3340 18932 3392
rect 19432 3340 19484 3392
rect 23940 3476 23992 3528
rect 28816 3680 28868 3732
rect 31668 3680 31720 3732
rect 31944 3723 31996 3732
rect 31944 3689 31953 3723
rect 31953 3689 31987 3723
rect 31987 3689 31996 3723
rect 31944 3680 31996 3689
rect 32036 3680 32088 3732
rect 33232 3680 33284 3732
rect 34244 3723 34296 3732
rect 34244 3689 34253 3723
rect 34253 3689 34287 3723
rect 34287 3689 34296 3723
rect 34244 3680 34296 3689
rect 26424 3612 26476 3664
rect 27896 3612 27948 3664
rect 29644 3612 29696 3664
rect 29920 3612 29972 3664
rect 31576 3612 31628 3664
rect 32312 3612 32364 3664
rect 33784 3612 33836 3664
rect 36820 3612 36872 3664
rect 24308 3544 24360 3596
rect 24584 3544 24636 3596
rect 26332 3544 26384 3596
rect 26516 3544 26568 3596
rect 31208 3544 31260 3596
rect 31484 3587 31536 3596
rect 31484 3553 31493 3587
rect 31493 3553 31527 3587
rect 31527 3553 31536 3587
rect 31484 3544 31536 3553
rect 34060 3544 34112 3596
rect 37556 3544 37608 3596
rect 24216 3476 24268 3528
rect 29000 3519 29052 3528
rect 19984 3408 20036 3460
rect 20904 3408 20956 3460
rect 22192 3408 22244 3460
rect 22560 3451 22612 3460
rect 22560 3417 22569 3451
rect 22569 3417 22603 3451
rect 22603 3417 22612 3451
rect 22560 3408 22612 3417
rect 27068 3451 27120 3460
rect 27068 3417 27077 3451
rect 27077 3417 27111 3451
rect 27111 3417 27120 3451
rect 27068 3408 27120 3417
rect 27252 3408 27304 3460
rect 29000 3485 29009 3519
rect 29009 3485 29043 3519
rect 29043 3485 29052 3519
rect 29000 3476 29052 3485
rect 29828 3476 29880 3528
rect 34244 3476 34296 3528
rect 36636 3476 36688 3528
rect 36820 3519 36872 3528
rect 36820 3485 36829 3519
rect 36829 3485 36863 3519
rect 36863 3485 36872 3519
rect 36820 3476 36872 3485
rect 21180 3340 21232 3392
rect 23848 3383 23900 3392
rect 23848 3349 23857 3383
rect 23857 3349 23891 3383
rect 23891 3349 23900 3383
rect 23848 3340 23900 3349
rect 23940 3340 23992 3392
rect 26700 3340 26752 3392
rect 28080 3383 28132 3392
rect 28080 3349 28089 3383
rect 28089 3349 28123 3383
rect 28123 3349 28132 3383
rect 28080 3340 28132 3349
rect 29736 3340 29788 3392
rect 30564 3340 30616 3392
rect 30932 3408 30984 3460
rect 31300 3408 31352 3460
rect 31576 3408 31628 3460
rect 33324 3408 33376 3460
rect 33416 3451 33468 3460
rect 33416 3417 33425 3451
rect 33425 3417 33459 3451
rect 33459 3417 33468 3451
rect 33416 3408 33468 3417
rect 33876 3408 33928 3460
rect 35992 3408 36044 3460
rect 34980 3383 35032 3392
rect 34980 3349 34989 3383
rect 34989 3349 35023 3383
rect 35023 3349 35032 3383
rect 34980 3340 35032 3349
rect 35624 3383 35676 3392
rect 35624 3349 35633 3383
rect 35633 3349 35667 3383
rect 35667 3349 35676 3383
rect 35624 3340 35676 3349
rect 36268 3383 36320 3392
rect 36268 3349 36277 3383
rect 36277 3349 36311 3383
rect 36311 3349 36320 3383
rect 36268 3340 36320 3349
rect 37556 3383 37608 3392
rect 37556 3349 37565 3383
rect 37565 3349 37599 3383
rect 37599 3349 37608 3383
rect 37556 3340 37608 3349
rect 38200 3383 38252 3392
rect 38200 3349 38209 3383
rect 38209 3349 38243 3383
rect 38243 3349 38252 3383
rect 38200 3340 38252 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2320 3000 2372 3052
rect 11612 3136 11664 3188
rect 12532 3179 12584 3188
rect 12532 3145 12541 3179
rect 12541 3145 12575 3179
rect 12575 3145 12584 3179
rect 12532 3136 12584 3145
rect 16580 3136 16632 3188
rect 16948 3179 17000 3188
rect 16948 3145 16957 3179
rect 16957 3145 16991 3179
rect 16991 3145 17000 3179
rect 16948 3136 17000 3145
rect 10600 3111 10652 3120
rect 10600 3077 10609 3111
rect 10609 3077 10643 3111
rect 10643 3077 10652 3111
rect 10600 3068 10652 3077
rect 13636 3068 13688 3120
rect 10048 3000 10100 3052
rect 11796 3043 11848 3052
rect 11796 3009 11805 3043
rect 11805 3009 11839 3043
rect 11839 3009 11848 3043
rect 11796 3000 11848 3009
rect 12440 3043 12492 3052
rect 12440 3009 12449 3043
rect 12449 3009 12483 3043
rect 12483 3009 12492 3043
rect 12440 3000 12492 3009
rect 14004 3043 14056 3052
rect 14004 3009 14013 3043
rect 14013 3009 14047 3043
rect 14047 3009 14056 3043
rect 14004 3000 14056 3009
rect 14280 3000 14332 3052
rect 16120 3068 16172 3120
rect 15752 3000 15804 3052
rect 21272 3136 21324 3188
rect 21364 3136 21416 3188
rect 22192 3136 22244 3188
rect 17776 3111 17828 3120
rect 17776 3077 17785 3111
rect 17785 3077 17819 3111
rect 17819 3077 17828 3111
rect 17776 3068 17828 3077
rect 19064 3068 19116 3120
rect 20260 3068 20312 3120
rect 24032 3068 24084 3120
rect 27804 3068 27856 3120
rect 28080 3136 28132 3188
rect 29276 3136 29328 3188
rect 28908 3068 28960 3120
rect 29368 3068 29420 3120
rect 29736 3068 29788 3120
rect 17500 3043 17552 3052
rect 14188 2975 14240 2984
rect 14188 2941 14197 2975
rect 14197 2941 14231 2975
rect 14231 2941 14240 2975
rect 14188 2932 14240 2941
rect 17500 3009 17509 3043
rect 17509 3009 17543 3043
rect 17543 3009 17552 3043
rect 17500 3000 17552 3009
rect 19156 3000 19208 3052
rect 21088 3000 21140 3052
rect 22008 3043 22060 3052
rect 22008 3009 22017 3043
rect 22017 3009 22051 3043
rect 22051 3009 22060 3043
rect 22008 3000 22060 3009
rect 23388 3000 23440 3052
rect 24584 3043 24636 3052
rect 24584 3009 24593 3043
rect 24593 3009 24627 3043
rect 24627 3009 24636 3043
rect 24584 3000 24636 3009
rect 26240 3000 26292 3052
rect 27252 3043 27304 3052
rect 17408 2932 17460 2984
rect 17868 2932 17920 2984
rect 19984 2932 20036 2984
rect 21272 2932 21324 2984
rect 23664 2932 23716 2984
rect 25228 2932 25280 2984
rect 27252 3009 27261 3043
rect 27261 3009 27295 3043
rect 27295 3009 27304 3043
rect 27252 3000 27304 3009
rect 27988 3000 28040 3052
rect 31484 3068 31536 3120
rect 32220 3136 32272 3188
rect 36084 3136 36136 3188
rect 37556 3136 37608 3188
rect 32680 3068 32732 3120
rect 37280 3068 37332 3120
rect 37740 3068 37792 3120
rect 31760 3043 31812 3052
rect 26792 2932 26844 2984
rect 31300 2932 31352 2984
rect 19248 2907 19300 2916
rect 19248 2873 19257 2907
rect 19257 2873 19291 2907
rect 19291 2873 19300 2907
rect 19248 2864 19300 2873
rect 23572 2864 23624 2916
rect 31760 3009 31769 3043
rect 31769 3009 31803 3043
rect 31803 3009 31812 3043
rect 31760 3000 31812 3009
rect 34612 3000 34664 3052
rect 35808 3000 35860 3052
rect 36084 3000 36136 3052
rect 31484 2932 31536 2984
rect 31760 2864 31812 2916
rect 1308 2796 1360 2848
rect 2780 2796 2832 2848
rect 3056 2839 3108 2848
rect 3056 2805 3065 2839
rect 3065 2805 3099 2839
rect 3099 2805 3108 2839
rect 3056 2796 3108 2805
rect 9680 2839 9732 2848
rect 9680 2805 9689 2839
rect 9689 2805 9723 2839
rect 9723 2805 9732 2839
rect 9680 2796 9732 2805
rect 11888 2839 11940 2848
rect 11888 2805 11897 2839
rect 11897 2805 11931 2839
rect 11931 2805 11940 2839
rect 11888 2796 11940 2805
rect 12440 2796 12492 2848
rect 21364 2796 21416 2848
rect 21548 2796 21600 2848
rect 30196 2796 30248 2848
rect 30288 2796 30340 2848
rect 30564 2796 30616 2848
rect 34336 2864 34388 2916
rect 34428 2864 34480 2916
rect 34244 2796 34296 2848
rect 34520 2796 34572 2848
rect 34704 2796 34756 2848
rect 37372 3000 37424 3052
rect 36636 2839 36688 2848
rect 36636 2805 36645 2839
rect 36645 2805 36679 2839
rect 36679 2805 36688 2839
rect 36636 2796 36688 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 10048 2635 10100 2644
rect 10048 2601 10057 2635
rect 10057 2601 10091 2635
rect 10091 2601 10100 2635
rect 10048 2592 10100 2601
rect 12900 2635 12952 2644
rect 12900 2601 12909 2635
rect 12909 2601 12943 2635
rect 12943 2601 12952 2635
rect 12900 2592 12952 2601
rect 16764 2592 16816 2644
rect 19064 2592 19116 2644
rect 20076 2592 20128 2644
rect 20996 2592 21048 2644
rect 23664 2592 23716 2644
rect 30380 2592 30432 2644
rect 31116 2592 31168 2644
rect 10600 2524 10652 2576
rect 13360 2524 13412 2576
rect 19984 2524 20036 2576
rect 2504 2456 2556 2508
rect 4068 2499 4120 2508
rect 4068 2465 4077 2499
rect 4077 2465 4111 2499
rect 4111 2465 4120 2499
rect 4068 2456 4120 2465
rect 20 2388 72 2440
rect 3056 2388 3108 2440
rect 9772 2456 9824 2508
rect 6552 2431 6604 2440
rect 6552 2397 6561 2431
rect 6561 2397 6595 2431
rect 6595 2397 6604 2431
rect 6552 2388 6604 2397
rect 9680 2388 9732 2440
rect 11060 2388 11112 2440
rect 14004 2388 14056 2440
rect 17040 2456 17092 2508
rect 17592 2499 17644 2508
rect 17592 2465 17601 2499
rect 17601 2465 17635 2499
rect 17635 2465 17644 2499
rect 17592 2456 17644 2465
rect 22008 2456 22060 2508
rect 24584 2456 24636 2508
rect 25964 2456 26016 2508
rect 29736 2499 29788 2508
rect 29736 2465 29745 2499
rect 29745 2465 29779 2499
rect 29779 2465 29788 2499
rect 29736 2456 29788 2465
rect 31392 2456 31444 2508
rect 16856 2388 16908 2440
rect 17408 2431 17460 2440
rect 17408 2397 17417 2431
rect 17417 2397 17451 2431
rect 17451 2397 17460 2431
rect 17408 2388 17460 2397
rect 18880 2431 18932 2440
rect 18880 2397 18889 2431
rect 18889 2397 18923 2431
rect 18923 2397 18932 2431
rect 18880 2388 18932 2397
rect 27068 2388 27120 2440
rect 27436 2431 27488 2440
rect 27436 2397 27445 2431
rect 27445 2397 27479 2431
rect 27479 2397 27488 2431
rect 27436 2388 27488 2397
rect 3240 2295 3292 2304
rect 3240 2261 3249 2295
rect 3249 2261 3283 2295
rect 3283 2261 3292 2295
rect 3240 2252 3292 2261
rect 4528 2252 4580 2304
rect 6460 2252 6512 2304
rect 8392 2252 8444 2304
rect 13544 2320 13596 2372
rect 14556 2363 14608 2372
rect 14556 2329 14565 2363
rect 14565 2329 14599 2363
rect 14599 2329 14608 2363
rect 14556 2320 14608 2329
rect 20628 2320 20680 2372
rect 11612 2252 11664 2304
rect 14832 2252 14884 2304
rect 16764 2252 16816 2304
rect 18972 2252 19024 2304
rect 23388 2320 23440 2372
rect 23572 2320 23624 2372
rect 26792 2320 26844 2372
rect 27712 2363 27764 2372
rect 26976 2252 27028 2304
rect 27712 2329 27721 2363
rect 27721 2329 27755 2363
rect 27755 2329 27764 2363
rect 27712 2320 27764 2329
rect 29920 2320 29972 2372
rect 31300 2320 31352 2372
rect 34704 2592 34756 2644
rect 32588 2524 32640 2576
rect 33784 2499 33836 2508
rect 33784 2465 33793 2499
rect 33793 2465 33827 2499
rect 33827 2465 33836 2499
rect 33784 2456 33836 2465
rect 34060 2499 34112 2508
rect 34060 2465 34069 2499
rect 34069 2465 34103 2499
rect 34103 2465 34112 2499
rect 34060 2456 34112 2465
rect 35808 2456 35860 2508
rect 37648 2456 37700 2508
rect 38384 2456 38436 2508
rect 36636 2431 36688 2440
rect 33324 2320 33376 2372
rect 33692 2320 33744 2372
rect 36636 2397 36645 2431
rect 36645 2397 36679 2431
rect 36679 2397 36688 2431
rect 36636 2388 36688 2397
rect 39304 2388 39356 2440
rect 34152 2252 34204 2304
rect 35440 2252 35492 2304
rect 37188 2252 37240 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 21824 2048 21876 2100
rect 26792 2048 26844 2100
rect 26884 2048 26936 2100
rect 35624 2048 35676 2100
rect 14556 1980 14608 2032
rect 32404 1980 32456 2032
rect 21640 1912 21692 1964
rect 26884 1912 26936 1964
rect 26976 1912 27028 1964
rect 35348 1912 35400 1964
rect 11888 1844 11940 1896
rect 23572 1844 23624 1896
rect 19064 1776 19116 1828
rect 35900 1844 35952 1896
rect 29920 1776 29972 1828
rect 37004 1776 37056 1828
rect 27712 1708 27764 1760
rect 33508 1708 33560 1760
rect 34244 1708 34296 1760
rect 32404 1640 32456 1692
rect 34612 1640 34664 1692
<< metal2 >>
rect 1306 39200 1362 39800
rect 2594 39200 2650 39800
rect 2870 39536 2926 39545
rect 2870 39471 2926 39480
rect 1320 37346 1348 39200
rect 1674 37496 1730 37505
rect 1674 37431 1730 37440
rect 1320 37318 1440 37346
rect 1412 37262 1440 37318
rect 1400 37256 1452 37262
rect 1400 37198 1452 37204
rect 1688 36854 1716 37431
rect 2504 37256 2556 37262
rect 2504 37198 2556 37204
rect 2608 37210 2636 39200
rect 1768 37120 1820 37126
rect 1768 37062 1820 37068
rect 1676 36848 1728 36854
rect 1676 36790 1728 36796
rect 1674 36136 1730 36145
rect 1674 36071 1730 36080
rect 1688 36038 1716 36071
rect 1676 36032 1728 36038
rect 1676 35974 1728 35980
rect 1676 34400 1728 34406
rect 1676 34342 1728 34348
rect 1688 34105 1716 34342
rect 1674 34096 1730 34105
rect 1674 34031 1730 34040
rect 1676 32224 1728 32230
rect 1676 32166 1728 32172
rect 1688 32065 1716 32166
rect 1674 32056 1730 32065
rect 1674 31991 1730 32000
rect 1674 30696 1730 30705
rect 1674 30631 1676 30640
rect 1728 30631 1730 30640
rect 1676 30602 1728 30608
rect 1688 30394 1716 30602
rect 1676 30388 1728 30394
rect 1676 30330 1728 30336
rect 1584 29164 1636 29170
rect 1584 29106 1636 29112
rect 1596 28694 1624 29106
rect 1584 28688 1636 28694
rect 1582 28656 1584 28665
rect 1636 28656 1638 28665
rect 1582 28591 1638 28600
rect 1676 26784 1728 26790
rect 1676 26726 1728 26732
rect 1688 26625 1716 26726
rect 1674 26616 1730 26625
rect 1674 26551 1730 26560
rect 1584 25288 1636 25294
rect 1582 25256 1584 25265
rect 1636 25256 1638 25265
rect 1582 25191 1638 25200
rect 1596 24954 1624 25191
rect 1584 24948 1636 24954
rect 1584 24890 1636 24896
rect 1584 23656 1636 23662
rect 1584 23598 1636 23604
rect 1596 23254 1624 23598
rect 1584 23248 1636 23254
rect 1582 23216 1584 23225
rect 1636 23216 1638 23225
rect 1582 23151 1638 23160
rect 1780 21706 1808 37062
rect 2136 36644 2188 36650
rect 2136 36586 2188 36592
rect 1860 36168 1912 36174
rect 1860 36110 1912 36116
rect 1872 34746 1900 36110
rect 1860 34740 1912 34746
rect 1860 34682 1912 34688
rect 2044 34604 2096 34610
rect 2044 34546 2096 34552
rect 1952 30728 2004 30734
rect 1952 30670 2004 30676
rect 1964 26234 1992 30670
rect 1872 26206 1992 26234
rect 1872 23662 1900 26206
rect 2056 25498 2084 34546
rect 2044 25492 2096 25498
rect 2044 25434 2096 25440
rect 1952 25288 2004 25294
rect 1952 25230 2004 25236
rect 1860 23656 1912 23662
rect 1860 23598 1912 23604
rect 1596 21678 1808 21706
rect 1596 17202 1624 21678
rect 1768 21548 1820 21554
rect 1768 21490 1820 21496
rect 1676 21344 1728 21350
rect 1676 21286 1728 21292
rect 1688 21185 1716 21286
rect 1674 21176 1730 21185
rect 1780 21146 1808 21490
rect 1674 21111 1730 21120
rect 1768 21140 1820 21146
rect 1768 21082 1820 21088
rect 1674 19816 1730 19825
rect 1674 19751 1676 19760
rect 1728 19751 1730 19760
rect 1676 19722 1728 19728
rect 1688 19514 1716 19722
rect 1676 19508 1728 19514
rect 1676 19450 1728 19456
rect 1872 18766 1900 23598
rect 1964 20942 1992 25230
rect 1952 20936 2004 20942
rect 1952 20878 2004 20884
rect 1964 19378 1992 20878
rect 1952 19372 2004 19378
rect 1952 19314 2004 19320
rect 1860 18760 1912 18766
rect 1860 18702 1912 18708
rect 2148 18426 2176 36586
rect 2516 30938 2544 37198
rect 2608 37182 2820 37210
rect 2792 37126 2820 37182
rect 2780 37120 2832 37126
rect 2780 37062 2832 37068
rect 2884 36922 2912 39471
rect 4526 39200 4582 39800
rect 6458 39200 6514 39800
rect 7746 39200 7802 39800
rect 9678 39200 9734 39800
rect 11610 39200 11666 39800
rect 12898 39200 12954 39800
rect 14830 39200 14886 39800
rect 16762 39200 16818 39800
rect 18050 39200 18106 39800
rect 19982 39200 20038 39800
rect 21914 39200 21970 39800
rect 23202 39200 23258 39800
rect 25134 39200 25190 39800
rect 27066 39200 27122 39800
rect 28354 39200 28410 39800
rect 30286 39200 30342 39800
rect 32218 39200 32274 39800
rect 33506 39200 33562 39800
rect 35438 39200 35494 39800
rect 37370 39200 37426 39800
rect 38658 39200 38714 39800
rect 4540 37754 4568 39200
rect 4540 37726 4660 37754
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4632 37126 4660 37726
rect 6472 37262 6500 39200
rect 6552 37324 6604 37330
rect 6552 37266 6604 37272
rect 6460 37256 6512 37262
rect 6460 37198 6512 37204
rect 4620 37120 4672 37126
rect 4620 37062 4672 37068
rect 5448 37120 5500 37126
rect 5448 37062 5500 37068
rect 2872 36916 2924 36922
rect 2872 36858 2924 36864
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 2504 30932 2556 30938
rect 2504 30874 2556 30880
rect 2228 30660 2280 30666
rect 2228 30602 2280 30608
rect 2240 20466 2268 30602
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 5460 29510 5488 37062
rect 5448 29504 5500 29510
rect 5448 29446 5500 29452
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 2228 20460 2280 20466
rect 2228 20402 2280 20408
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 2136 18420 2188 18426
rect 2136 18362 2188 18368
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1688 17785 1716 18022
rect 1674 17776 1730 17785
rect 1674 17711 1730 17720
rect 1584 17196 1636 17202
rect 1584 17138 1636 17144
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 1688 15745 1716 15846
rect 1674 15736 1730 15745
rect 1674 15671 1730 15680
rect 2424 15638 2452 15846
rect 2412 15632 2464 15638
rect 2412 15574 2464 15580
rect 1952 15360 2004 15366
rect 1952 15302 2004 15308
rect 1584 14408 1636 14414
rect 1582 14376 1584 14385
rect 1636 14376 1638 14385
rect 1582 14311 1638 14320
rect 1596 14074 1624 14311
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1688 12345 1716 12582
rect 1674 12336 1730 12345
rect 1674 12271 1730 12280
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1688 10305 1716 10406
rect 1674 10296 1730 10305
rect 1674 10231 1730 10240
rect 1872 9110 1900 12242
rect 1860 9104 1912 9110
rect 1860 9046 1912 9052
rect 1674 8936 1730 8945
rect 1674 8871 1676 8880
rect 1728 8871 1730 8880
rect 1676 8842 1728 8848
rect 1688 8634 1716 8842
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1688 6905 1716 7142
rect 1964 6914 1992 15302
rect 4080 14618 4108 18226
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 1674 6896 1730 6905
rect 1674 6831 1730 6840
rect 1872 6886 1992 6914
rect 1872 5234 1900 6886
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1688 4865 1716 4966
rect 1674 4856 1730 4865
rect 1674 4791 1730 4800
rect 2332 3738 2360 13330
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 4080 9654 4108 12786
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 5552 11150 5580 14350
rect 6564 11898 6592 37266
rect 7760 37126 7788 39200
rect 9692 37262 9720 39200
rect 11520 37324 11572 37330
rect 11520 37266 11572 37272
rect 8116 37256 8168 37262
rect 8116 37198 8168 37204
rect 9680 37256 9732 37262
rect 9680 37198 9732 37204
rect 7748 37120 7800 37126
rect 7748 37062 7800 37068
rect 8128 36922 8156 37198
rect 10692 37188 10744 37194
rect 10692 37130 10744 37136
rect 8116 36916 8168 36922
rect 8116 36858 8168 36864
rect 10704 36786 10732 37130
rect 10692 36780 10744 36786
rect 10692 36722 10744 36728
rect 11532 35894 11560 37266
rect 11624 36786 11652 39200
rect 12912 37330 12940 39200
rect 12900 37324 12952 37330
rect 12900 37266 12952 37272
rect 14844 37126 14872 39200
rect 15200 37256 15252 37262
rect 15200 37198 15252 37204
rect 14832 37120 14884 37126
rect 14832 37062 14884 37068
rect 11612 36780 11664 36786
rect 11612 36722 11664 36728
rect 11624 36378 11652 36722
rect 11980 36712 12032 36718
rect 11980 36654 12032 36660
rect 11612 36372 11664 36378
rect 11612 36314 11664 36320
rect 11532 35866 11652 35894
rect 9128 32428 9180 32434
rect 9128 32370 9180 32376
rect 6828 26988 6880 26994
rect 6828 26930 6880 26936
rect 6840 21690 6868 26930
rect 9140 25498 9168 32370
rect 9128 25492 9180 25498
rect 9128 25434 9180 25440
rect 7840 25152 7892 25158
rect 7840 25094 7892 25100
rect 9772 25152 9824 25158
rect 9772 25094 9824 25100
rect 6828 21684 6880 21690
rect 6828 21626 6880 21632
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5736 10674 5764 11494
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2516 7410 2544 8434
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 1688 3398 1716 3431
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 2332 3058 2360 3674
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 1308 2848 1360 2854
rect 1308 2790 1360 2796
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 32 800 60 2382
rect 1320 800 1348 2790
rect 2516 2514 2544 7346
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 6380 6798 6408 11086
rect 7852 7449 7880 25094
rect 8300 17128 8352 17134
rect 8300 17070 8352 17076
rect 8312 12306 8340 17070
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 7838 7440 7894 7449
rect 7838 7375 7894 7384
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 2792 3534 2820 5510
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 2792 1465 2820 2790
rect 3068 2446 3096 2790
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4066 2544 4122 2553
rect 4066 2479 4068 2488
rect 4120 2479 4122 2488
rect 4068 2450 4120 2456
rect 6564 2446 6592 6598
rect 9784 6390 9812 25094
rect 10876 13796 10928 13802
rect 10876 13738 10928 13744
rect 10888 13394 10916 13738
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9692 2446 9720 2790
rect 9784 2514 9812 4966
rect 10060 3058 10088 7346
rect 10980 3738 11008 9590
rect 11624 4214 11652 35866
rect 11992 27470 12020 36654
rect 13084 34536 13136 34542
rect 13084 34478 13136 34484
rect 11980 27464 12032 27470
rect 11980 27406 12032 27412
rect 13096 20806 13124 34478
rect 15212 28150 15240 37198
rect 15568 37188 15620 37194
rect 15568 37130 15620 37136
rect 15580 28558 15608 37130
rect 16776 37126 16804 39200
rect 17316 37392 17368 37398
rect 17316 37334 17368 37340
rect 17132 37256 17184 37262
rect 17132 37198 17184 37204
rect 16764 37120 16816 37126
rect 16764 37062 16816 37068
rect 15568 28552 15620 28558
rect 15568 28494 15620 28500
rect 15660 28416 15712 28422
rect 15660 28358 15712 28364
rect 15200 28144 15252 28150
rect 15200 28086 15252 28092
rect 15568 27328 15620 27334
rect 15568 27270 15620 27276
rect 13544 21344 13596 21350
rect 13544 21286 13596 21292
rect 13084 20800 13136 20806
rect 13084 20742 13136 20748
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11716 16726 11744 17138
rect 11704 16720 11756 16726
rect 11704 16662 11756 16668
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 11888 5228 11940 5234
rect 11808 5188 11888 5216
rect 11808 4622 11836 5188
rect 11888 5170 11940 5176
rect 12438 5128 12494 5137
rect 12912 5114 12940 9862
rect 13096 9654 13124 17274
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13372 12986 13400 13262
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13372 12434 13400 12922
rect 13372 12406 13492 12434
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13372 10470 13400 11086
rect 13360 10464 13412 10470
rect 13360 10406 13412 10412
rect 13084 9648 13136 9654
rect 13084 9590 13136 9596
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 13096 5302 13124 5510
rect 13084 5296 13136 5302
rect 13084 5238 13136 5244
rect 12912 5086 13032 5114
rect 12438 5063 12440 5072
rect 12492 5063 12494 5072
rect 12440 5034 12492 5040
rect 12346 4856 12402 4865
rect 12346 4791 12348 4800
rect 12400 4791 12402 4800
rect 12348 4762 12400 4768
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11612 4208 11664 4214
rect 11612 4150 11664 4156
rect 11624 3738 11652 4150
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 10600 3120 10652 3126
rect 10600 3062 10652 3068
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 10060 2650 10088 2994
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 10612 2582 10640 3062
rect 10980 2802 11008 3674
rect 11624 3194 11652 3674
rect 11808 3534 11836 4558
rect 12254 4176 12310 4185
rect 12254 4111 12310 4120
rect 12268 3738 12296 4111
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11808 3058 11836 3470
rect 12544 3194 12572 4014
rect 12900 3596 12952 3602
rect 12900 3538 12952 3544
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12452 2854 12480 2994
rect 11888 2848 11940 2854
rect 10980 2774 11100 2802
rect 11888 2790 11940 2796
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 10600 2576 10652 2582
rect 10600 2518 10652 2524
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 11072 2446 11100 2774
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 3252 800 3280 2246
rect 4540 800 4568 2246
rect 6472 800 6500 2246
rect 8404 800 8432 2246
rect 9692 800 9720 2382
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11624 800 11652 2246
rect 11900 1902 11928 2790
rect 12912 2650 12940 3538
rect 13004 3534 13032 5086
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 13004 3398 13032 3470
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 13372 2582 13400 10406
rect 13464 9654 13492 12406
rect 13556 11150 13584 21286
rect 14740 16108 14792 16114
rect 14740 16050 14792 16056
rect 14752 15026 14780 16050
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 13728 14272 13780 14278
rect 13648 14232 13728 14260
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13452 9648 13504 9654
rect 13452 9590 13504 9596
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13464 5234 13492 5646
rect 13556 5370 13584 8910
rect 13648 7546 13676 14232
rect 13728 14214 13780 14220
rect 14016 14074 14044 14554
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13740 13530 13768 13874
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13740 12442 13768 13466
rect 13820 13252 13872 13258
rect 13820 13194 13872 13200
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13832 10470 13860 13194
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 14108 10198 14136 14350
rect 14752 13433 14780 14962
rect 15580 13734 15608 27270
rect 15672 17814 15700 28358
rect 17144 28218 17172 37198
rect 17132 28212 17184 28218
rect 17132 28154 17184 28160
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 15660 17808 15712 17814
rect 15660 17750 15712 17756
rect 15672 16794 15700 17750
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 16580 17604 16632 17610
rect 16580 17546 16632 17552
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 16028 15904 16080 15910
rect 16028 15846 16080 15852
rect 16040 15162 16068 15846
rect 16210 15464 16266 15473
rect 16210 15399 16212 15408
rect 16264 15399 16266 15408
rect 16212 15370 16264 15376
rect 16028 15156 16080 15162
rect 16028 15098 16080 15104
rect 15752 14884 15804 14890
rect 15752 14826 15804 14832
rect 15764 14346 15792 14826
rect 15752 14340 15804 14346
rect 15752 14282 15804 14288
rect 16040 14074 16068 15098
rect 16212 15088 16264 15094
rect 16212 15030 16264 15036
rect 16120 14544 16172 14550
rect 16120 14486 16172 14492
rect 16132 14346 16160 14486
rect 16120 14340 16172 14346
rect 16120 14282 16172 14288
rect 16224 14074 16252 15030
rect 16592 14958 16620 17546
rect 16868 17202 16896 17614
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16672 17060 16724 17066
rect 16672 17002 16724 17008
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16028 14068 16080 14074
rect 16028 14010 16080 14016
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 16316 13870 16344 14010
rect 16396 14000 16448 14006
rect 16448 13948 16620 13954
rect 16396 13942 16620 13948
rect 16408 13938 16620 13942
rect 16408 13932 16632 13938
rect 16408 13926 16580 13932
rect 16580 13874 16632 13880
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 15568 13728 15620 13734
rect 15752 13728 15804 13734
rect 15620 13676 15700 13682
rect 15568 13670 15700 13676
rect 15752 13670 15804 13676
rect 15580 13654 15700 13670
rect 15672 13530 15700 13654
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 14738 13424 14794 13433
rect 14738 13359 14794 13368
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14292 11762 14320 12378
rect 14476 12238 14504 12922
rect 15672 12918 15700 13466
rect 15764 13394 15792 13670
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15856 12918 15884 13126
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 15844 12912 15896 12918
rect 15844 12854 15896 12860
rect 16028 12912 16080 12918
rect 16028 12854 16080 12860
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14936 12102 14964 12786
rect 15752 12708 15804 12714
rect 15752 12650 15804 12656
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14292 11014 14320 11086
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14648 10736 14700 10742
rect 14648 10678 14700 10684
rect 14660 10266 14688 10678
rect 14830 10568 14886 10577
rect 14830 10503 14886 10512
rect 14648 10260 14700 10266
rect 14648 10202 14700 10208
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 14096 10192 14148 10198
rect 14752 10146 14780 10202
rect 14096 10134 14148 10140
rect 14108 8566 14136 10134
rect 14568 10118 14780 10146
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 14096 8560 14148 8566
rect 14096 8502 14148 8508
rect 14108 8362 14136 8502
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 14200 7478 14228 9522
rect 14278 9072 14334 9081
rect 14278 9007 14334 9016
rect 14292 8974 14320 9007
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14384 8634 14412 8774
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14568 8566 14596 10118
rect 14556 8560 14608 8566
rect 14556 8502 14608 8508
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14188 7472 14240 7478
rect 14188 7414 14240 7420
rect 13820 6384 13872 6390
rect 13820 6326 13872 6332
rect 13544 5364 13596 5370
rect 13544 5306 13596 5312
rect 13452 5228 13504 5234
rect 13452 5170 13504 5176
rect 13464 4622 13492 5170
rect 13832 4826 13860 6326
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14476 5710 14504 6054
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14370 5400 14426 5409
rect 14370 5335 14426 5344
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13924 4622 13952 5170
rect 14384 5030 14412 5335
rect 14476 5234 14504 5646
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13912 4616 13964 4622
rect 13912 4558 13964 4564
rect 13464 4146 13492 4558
rect 14280 4208 14332 4214
rect 14280 4150 14332 4156
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13636 4004 13688 4010
rect 13636 3946 13688 3952
rect 13648 3126 13676 3946
rect 14292 3738 14320 4150
rect 14568 4078 14596 8366
rect 14648 7948 14700 7954
rect 14648 7890 14700 7896
rect 14660 6730 14688 7890
rect 14648 6724 14700 6730
rect 14648 6666 14700 6672
rect 14660 5778 14688 6666
rect 14844 5914 14872 10503
rect 14936 9674 14964 12038
rect 15212 11898 15240 12038
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15764 11830 15792 12650
rect 16040 12238 16068 12854
rect 16488 12640 16540 12646
rect 16488 12582 16540 12588
rect 15844 12232 15896 12238
rect 15842 12200 15844 12209
rect 16028 12232 16080 12238
rect 15896 12200 15898 12209
rect 16028 12174 16080 12180
rect 15842 12135 15898 12144
rect 15752 11824 15804 11830
rect 15752 11766 15804 11772
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15016 11076 15068 11082
rect 15016 11018 15068 11024
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 15028 10606 15056 11018
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 15120 10538 15148 11018
rect 15488 11014 15516 11290
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15476 11008 15528 11014
rect 15476 10950 15528 10956
rect 15108 10532 15160 10538
rect 15108 10474 15160 10480
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 14936 9646 15056 9674
rect 14924 9580 14976 9586
rect 14924 9522 14976 9528
rect 14936 8974 14964 9522
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 15028 7954 15056 9646
rect 15120 8838 15148 9862
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15212 8294 15240 10950
rect 15488 9518 15516 10950
rect 15476 9512 15528 9518
rect 15290 9480 15346 9489
rect 15476 9454 15528 9460
rect 15290 9415 15346 9424
rect 15200 8288 15252 8294
rect 15200 8230 15252 8236
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 15028 7546 15056 7890
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 15304 6866 15332 9415
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 15488 6458 15516 7686
rect 15580 7206 15608 11698
rect 16040 11626 16068 12174
rect 16304 12164 16356 12170
rect 16304 12106 16356 12112
rect 16316 11937 16344 12106
rect 16302 11928 16358 11937
rect 16302 11863 16358 11872
rect 16396 11688 16448 11694
rect 16396 11630 16448 11636
rect 15660 11620 15712 11626
rect 15660 11562 15712 11568
rect 16028 11620 16080 11626
rect 16028 11562 16080 11568
rect 15672 11354 15700 11562
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15844 10532 15896 10538
rect 15844 10474 15896 10480
rect 15658 10160 15714 10169
rect 15856 10130 15884 10474
rect 15658 10095 15660 10104
rect 15712 10095 15714 10104
rect 15844 10124 15896 10130
rect 15660 10066 15712 10072
rect 15844 10066 15896 10072
rect 15660 9988 15712 9994
rect 15660 9930 15712 9936
rect 15672 9761 15700 9930
rect 15658 9752 15714 9761
rect 15658 9687 15714 9696
rect 15936 9036 15988 9042
rect 15936 8978 15988 8984
rect 15948 8906 15976 8978
rect 15936 8900 15988 8906
rect 15936 8842 15988 8848
rect 15844 8832 15896 8838
rect 15844 8774 15896 8780
rect 15752 8560 15804 8566
rect 15752 8502 15804 8508
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15764 6866 15792 8502
rect 15856 8430 15884 8774
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15844 6724 15896 6730
rect 15844 6666 15896 6672
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 15014 5672 15070 5681
rect 15014 5607 15070 5616
rect 15028 5370 15056 5607
rect 15016 5364 15068 5370
rect 15016 5306 15068 5312
rect 15856 5234 15884 6666
rect 16040 5778 16068 11562
rect 16408 11218 16436 11630
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 16500 11082 16528 12582
rect 16684 12209 16712 17002
rect 16960 16046 16988 19314
rect 17224 16516 17276 16522
rect 17224 16458 17276 16464
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 16960 14958 16988 15982
rect 17236 15570 17264 16458
rect 17224 15564 17276 15570
rect 17224 15506 17276 15512
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16764 14884 16816 14890
rect 16764 14826 16816 14832
rect 16670 12200 16726 12209
rect 16670 12135 16726 12144
rect 16684 11370 16712 12135
rect 16776 12050 16804 14826
rect 17236 14550 17264 15506
rect 17224 14544 17276 14550
rect 17224 14486 17276 14492
rect 17040 14408 17092 14414
rect 17040 14350 17092 14356
rect 16948 13864 17000 13870
rect 16948 13806 17000 13812
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16868 12209 16896 12242
rect 16854 12200 16910 12209
rect 16960 12170 16988 13806
rect 17052 12782 17080 14350
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 16854 12135 16910 12144
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16776 12022 16896 12050
rect 16684 11342 16804 11370
rect 16488 11076 16540 11082
rect 16488 11018 16540 11024
rect 16776 11014 16804 11342
rect 16764 11008 16816 11014
rect 16764 10950 16816 10956
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16132 10470 16160 10610
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16132 9722 16160 10406
rect 16868 10169 16896 12022
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 17052 10674 17080 11494
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 16854 10160 16910 10169
rect 16854 10095 16910 10104
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16592 9926 16620 9998
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16316 9489 16344 9522
rect 16302 9480 16358 9489
rect 16302 9415 16358 9424
rect 16396 8288 16448 8294
rect 16394 8256 16396 8265
rect 16448 8256 16450 8265
rect 16394 8191 16450 8200
rect 16500 6730 16528 9862
rect 16592 9654 16620 9862
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 16672 9444 16724 9450
rect 16672 9386 16724 9392
rect 16764 9444 16816 9450
rect 16764 9386 16816 9392
rect 16684 9353 16712 9386
rect 16670 9344 16726 9353
rect 16670 9279 16726 9288
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16580 8560 16632 8566
rect 16580 8502 16632 8508
rect 16592 6866 16620 8502
rect 16684 8294 16712 8910
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 16684 8022 16712 8230
rect 16672 8016 16724 8022
rect 16672 7958 16724 7964
rect 16776 7410 16804 9386
rect 17052 9178 17080 9590
rect 17144 9518 17172 13874
rect 17236 13297 17264 14486
rect 17222 13288 17278 13297
rect 17328 13258 17356 37334
rect 18064 37126 18092 39200
rect 18420 37256 18472 37262
rect 18420 37198 18472 37204
rect 18052 37120 18104 37126
rect 18052 37062 18104 37068
rect 18432 28762 18460 37198
rect 19996 37126 20024 39200
rect 21928 37330 21956 39200
rect 21916 37324 21968 37330
rect 21916 37266 21968 37272
rect 23216 37262 23244 39200
rect 25148 37262 25176 39200
rect 20352 37256 20404 37262
rect 20352 37198 20404 37204
rect 22284 37256 22336 37262
rect 22284 37198 22336 37204
rect 23204 37256 23256 37262
rect 23204 37198 23256 37204
rect 25136 37256 25188 37262
rect 25136 37198 25188 37204
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 18420 28756 18472 28762
rect 18420 28698 18472 28704
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 18512 28076 18564 28082
rect 18512 28018 18564 28024
rect 18524 27334 18552 28018
rect 18512 27328 18564 27334
rect 18512 27270 18564 27276
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 20364 24206 20392 37198
rect 22296 36786 22324 37198
rect 23216 36922 23244 37198
rect 26332 37188 26384 37194
rect 26332 37130 26384 37136
rect 25412 37120 25464 37126
rect 25412 37062 25464 37068
rect 23204 36916 23256 36922
rect 23204 36858 23256 36864
rect 22284 36780 22336 36786
rect 22284 36722 22336 36728
rect 22296 28082 22324 36722
rect 23664 29504 23716 29510
rect 23664 29446 23716 29452
rect 23112 28416 23164 28422
rect 23112 28358 23164 28364
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22928 27872 22980 27878
rect 22928 27814 22980 27820
rect 21456 27328 21508 27334
rect 21456 27270 21508 27276
rect 20352 24200 20404 24206
rect 20352 24142 20404 24148
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 21272 21344 21324 21350
rect 21272 21286 21324 21292
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19444 18970 19472 19654
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 18328 18692 18380 18698
rect 18328 18634 18380 18640
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17512 18358 17540 18566
rect 17500 18352 17552 18358
rect 17500 18294 17552 18300
rect 17592 18352 17644 18358
rect 17592 18294 17644 18300
rect 17604 17882 17632 18294
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17592 17876 17644 17882
rect 17592 17818 17644 17824
rect 17684 17128 17736 17134
rect 17684 17070 17736 17076
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17420 15434 17448 16934
rect 17696 16794 17724 17070
rect 17776 17060 17828 17066
rect 17776 17002 17828 17008
rect 17684 16788 17736 16794
rect 17684 16730 17736 16736
rect 17788 16658 17816 17002
rect 17776 16652 17828 16658
rect 17776 16594 17828 16600
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17788 15434 17816 15846
rect 17408 15428 17460 15434
rect 17408 15370 17460 15376
rect 17776 15428 17828 15434
rect 17776 15370 17828 15376
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 17420 14414 17448 14894
rect 17592 14884 17644 14890
rect 17592 14826 17644 14832
rect 17500 14612 17552 14618
rect 17500 14554 17552 14560
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17420 13870 17448 14214
rect 17512 13938 17540 14554
rect 17604 14482 17632 14826
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17592 14272 17644 14278
rect 17592 14214 17644 14220
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17222 13223 17278 13232
rect 17316 13252 17368 13258
rect 17316 13194 17368 13200
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 17236 12889 17264 13126
rect 17328 12986 17356 13194
rect 17316 12980 17368 12986
rect 17316 12922 17368 12928
rect 17222 12880 17278 12889
rect 17222 12815 17278 12824
rect 17316 12776 17368 12782
rect 17316 12718 17368 12724
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 17040 9172 17092 9178
rect 17040 9114 17092 9120
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 16856 9104 16908 9110
rect 17144 9058 17172 9114
rect 16908 9052 17172 9058
rect 16856 9046 17172 9052
rect 16868 9030 17172 9046
rect 17236 8906 17264 10542
rect 17328 9926 17356 12718
rect 17512 12594 17540 13330
rect 17604 12918 17632 14214
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17592 12912 17644 12918
rect 17592 12854 17644 12860
rect 17512 12566 17632 12594
rect 17604 12306 17632 12566
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 17696 11830 17724 13262
rect 17684 11824 17736 11830
rect 17684 11766 17736 11772
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17420 11218 17448 11494
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17420 10130 17448 11154
rect 17788 10538 17816 15370
rect 17880 12986 17908 18022
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 18064 16182 18092 16934
rect 18156 16250 18184 18158
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18248 16726 18276 17478
rect 18236 16720 18288 16726
rect 18236 16662 18288 16668
rect 18144 16244 18196 16250
rect 18144 16186 18196 16192
rect 18052 16176 18104 16182
rect 18052 16118 18104 16124
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 17972 13802 18000 15030
rect 18064 14958 18092 16118
rect 18156 14958 18184 16186
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 18340 14362 18368 18634
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 19892 18216 19944 18222
rect 19890 18184 19892 18193
rect 19944 18184 19946 18193
rect 20180 18154 20208 18226
rect 19890 18119 19946 18128
rect 19984 18148 20036 18154
rect 19904 18086 19932 18119
rect 19984 18090 20036 18096
rect 20168 18148 20220 18154
rect 20168 18090 20220 18096
rect 19892 18080 19944 18086
rect 19892 18022 19944 18028
rect 19432 17808 19484 17814
rect 19432 17750 19484 17756
rect 19340 17536 19392 17542
rect 19340 17478 19392 17484
rect 19352 16998 19380 17478
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19352 16810 19380 16934
rect 19260 16782 19380 16810
rect 18788 16448 18840 16454
rect 18788 16390 18840 16396
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 18708 15570 18736 15982
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 18604 15428 18656 15434
rect 18604 15370 18656 15376
rect 18616 15162 18644 15370
rect 18800 15366 18828 16390
rect 19260 15994 19288 16782
rect 19340 16720 19392 16726
rect 19340 16662 19392 16668
rect 19352 16114 19380 16662
rect 19444 16232 19472 17750
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19996 16522 20024 18090
rect 20272 17814 20300 18566
rect 20260 17808 20312 17814
rect 20260 17750 20312 17756
rect 20168 17536 20220 17542
rect 20168 17478 20220 17484
rect 19984 16516 20036 16522
rect 19984 16458 20036 16464
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19444 16204 19564 16232
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 18972 15972 19024 15978
rect 19260 15966 19380 15994
rect 19352 15960 19380 15966
rect 19352 15932 19472 15960
rect 18972 15914 19024 15920
rect 18880 15428 18932 15434
rect 18880 15370 18932 15376
rect 18788 15360 18840 15366
rect 18788 15302 18840 15308
rect 18604 15156 18656 15162
rect 18604 15098 18656 15104
rect 18248 14346 18368 14362
rect 18892 14346 18920 15370
rect 18052 14340 18104 14346
rect 18052 14282 18104 14288
rect 18236 14340 18368 14346
rect 18288 14334 18368 14340
rect 18880 14340 18932 14346
rect 18236 14282 18288 14288
rect 18880 14282 18932 14288
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 18064 13258 18092 14282
rect 18248 13394 18276 14282
rect 18512 13456 18564 13462
rect 18512 13398 18564 13404
rect 18788 13456 18840 13462
rect 18788 13398 18840 13404
rect 18236 13388 18288 13394
rect 18236 13330 18288 13336
rect 18052 13252 18104 13258
rect 18052 13194 18104 13200
rect 18328 13252 18380 13258
rect 18328 13194 18380 13200
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17880 12374 17908 12718
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17880 11812 17908 12310
rect 17960 11824 18012 11830
rect 17880 11784 17960 11812
rect 17960 11766 18012 11772
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 17972 11082 18000 11630
rect 18156 11370 18184 12378
rect 18236 12300 18288 12306
rect 18236 12242 18288 12248
rect 18064 11342 18184 11370
rect 18064 11150 18092 11342
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 17960 11076 18012 11082
rect 17960 11018 18012 11024
rect 17868 11008 17920 11014
rect 17868 10950 17920 10956
rect 17776 10532 17828 10538
rect 17776 10474 17828 10480
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 17776 9988 17828 9994
rect 17776 9930 17828 9936
rect 17316 9920 17368 9926
rect 17788 9897 17816 9930
rect 17316 9862 17368 9868
rect 17774 9888 17830 9897
rect 17224 8900 17276 8906
rect 17224 8842 17276 8848
rect 17040 8560 17092 8566
rect 17040 8502 17092 8508
rect 17052 8090 17080 8502
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 17236 8022 17264 8842
rect 17224 8016 17276 8022
rect 17224 7958 17276 7964
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16488 6724 16540 6730
rect 16488 6666 16540 6672
rect 16578 6624 16634 6633
rect 16578 6559 16634 6568
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 15936 5636 15988 5642
rect 15936 5578 15988 5584
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 15844 5228 15896 5234
rect 15844 5170 15896 5176
rect 14648 5092 14700 5098
rect 14648 5034 14700 5040
rect 14660 4826 14688 5034
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14936 4622 14964 5170
rect 15948 4826 15976 5578
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 15292 4616 15344 4622
rect 15844 4616 15896 4622
rect 15292 4558 15344 4564
rect 15842 4584 15844 4593
rect 15896 4584 15898 4593
rect 15304 4146 15332 4558
rect 16040 4554 16068 4762
rect 15842 4519 15898 4528
rect 16028 4548 16080 4554
rect 15752 4276 15804 4282
rect 15752 4218 15804 4224
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14188 3664 14240 3670
rect 14188 3606 14240 3612
rect 13728 3528 13780 3534
rect 13726 3496 13728 3505
rect 13780 3496 13782 3505
rect 13726 3431 13782 3440
rect 13636 3120 13688 3126
rect 13636 3062 13688 3068
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 13360 2576 13412 2582
rect 13360 2518 13412 2524
rect 14016 2446 14044 2994
rect 14200 2990 14228 3606
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14292 3058 14320 3470
rect 15764 3058 15792 4218
rect 15856 4146 15884 4519
rect 16028 4490 16080 4496
rect 16132 4486 16160 6054
rect 16304 5772 16356 5778
rect 16304 5714 16356 5720
rect 15936 4480 15988 4486
rect 15936 4422 15988 4428
rect 16120 4480 16172 4486
rect 16120 4422 16172 4428
rect 15948 4282 15976 4422
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 16132 4146 16160 4422
rect 15844 4140 15896 4146
rect 15844 4082 15896 4088
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16132 4049 16160 4082
rect 16316 4078 16344 5714
rect 16592 5370 16620 6559
rect 16684 5574 16712 7278
rect 16960 6186 16988 7822
rect 17224 7472 17276 7478
rect 17224 7414 17276 7420
rect 17132 7268 17184 7274
rect 17132 7210 17184 7216
rect 17040 6248 17092 6254
rect 17040 6190 17092 6196
rect 16948 6180 17000 6186
rect 16948 6122 17000 6128
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 16764 5364 16816 5370
rect 16764 5306 16816 5312
rect 16776 5166 16804 5306
rect 17052 5234 17080 6190
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16672 4616 16724 4622
rect 16670 4584 16672 4593
rect 16724 4584 16726 4593
rect 16670 4519 16726 4528
rect 16304 4072 16356 4078
rect 16118 4040 16174 4049
rect 16304 4014 16356 4020
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16118 3975 16174 3984
rect 16132 3126 16160 3975
rect 16592 3194 16620 4014
rect 16764 3392 16816 3398
rect 16764 3334 16816 3340
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 16120 3120 16172 3126
rect 16120 3062 16172 3068
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 16776 2650 16804 3334
rect 16764 2644 16816 2650
rect 16764 2586 16816 2592
rect 16868 2446 16896 4966
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 16948 3460 17000 3466
rect 16948 3402 17000 3408
rect 16960 3194 16988 3402
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 17052 2514 17080 4082
rect 17144 3534 17172 7210
rect 17236 5846 17264 7414
rect 17328 7274 17356 9862
rect 17774 9823 17830 9832
rect 17592 9716 17644 9722
rect 17592 9658 17644 9664
rect 17604 9518 17632 9658
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 17420 8634 17448 9454
rect 17880 9382 17908 10950
rect 18248 10606 18276 12242
rect 18340 11218 18368 13194
rect 18524 12170 18552 13398
rect 18800 13258 18828 13398
rect 18788 13252 18840 13258
rect 18788 13194 18840 13200
rect 18892 12714 18920 14282
rect 18984 14006 19012 15914
rect 19156 15088 19208 15094
rect 19156 15030 19208 15036
rect 19064 15020 19116 15026
rect 19064 14962 19116 14968
rect 18972 14000 19024 14006
rect 18972 13942 19024 13948
rect 19076 13938 19104 14962
rect 19064 13932 19116 13938
rect 19064 13874 19116 13880
rect 19062 13288 19118 13297
rect 19062 13223 19118 13232
rect 19076 12782 19104 13223
rect 19064 12776 19116 12782
rect 19064 12718 19116 12724
rect 18880 12708 18932 12714
rect 18880 12650 18932 12656
rect 19168 12442 19196 15030
rect 19248 14816 19300 14822
rect 19248 14758 19300 14764
rect 19260 13190 19288 14758
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19248 13184 19300 13190
rect 19248 13126 19300 13132
rect 19352 12918 19380 13806
rect 19444 13734 19472 15932
rect 19536 15570 19564 16204
rect 20180 16182 20208 17478
rect 20168 16176 20220 16182
rect 20168 16118 20220 16124
rect 19800 16108 19852 16114
rect 19800 16050 19852 16056
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 19812 15570 19840 16050
rect 19524 15564 19576 15570
rect 19524 15506 19576 15512
rect 19800 15564 19852 15570
rect 19800 15506 19852 15512
rect 19524 15428 19576 15434
rect 19708 15428 19760 15434
rect 19576 15388 19708 15416
rect 19524 15370 19576 15376
rect 19708 15370 19760 15376
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19996 14482 20024 16050
rect 20076 15156 20128 15162
rect 20076 15098 20128 15104
rect 19984 14476 20036 14482
rect 19984 14418 20036 14424
rect 20088 14414 20116 15098
rect 20364 15094 20392 20742
rect 20904 18080 20956 18086
rect 20904 18022 20956 18028
rect 20442 17912 20498 17921
rect 20442 17847 20498 17856
rect 20456 17678 20484 17847
rect 20444 17672 20496 17678
rect 20444 17614 20496 17620
rect 20916 17610 20944 18022
rect 20812 17604 20864 17610
rect 20812 17546 20864 17552
rect 20904 17604 20956 17610
rect 20904 17546 20956 17552
rect 21088 17604 21140 17610
rect 21088 17546 21140 17552
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20548 16998 20576 17138
rect 20536 16992 20588 16998
rect 20536 16934 20588 16940
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 20534 16008 20590 16017
rect 20534 15943 20590 15952
rect 20548 15910 20576 15943
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 20640 15502 20668 16186
rect 20628 15496 20680 15502
rect 20628 15438 20680 15444
rect 20732 15094 20760 16934
rect 20824 16454 20852 17546
rect 20996 17128 21048 17134
rect 20996 17070 21048 17076
rect 21008 16658 21036 17070
rect 20996 16652 21048 16658
rect 20996 16594 21048 16600
rect 20812 16448 20864 16454
rect 20812 16390 20864 16396
rect 21100 15978 21128 17546
rect 21284 17202 21312 21286
rect 21364 19168 21416 19174
rect 21364 19110 21416 19116
rect 21376 18834 21404 19110
rect 21364 18828 21416 18834
rect 21364 18770 21416 18776
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 21468 16561 21496 27270
rect 22836 22976 22888 22982
rect 22836 22918 22888 22924
rect 22652 21888 22704 21894
rect 22652 21830 22704 21836
rect 22008 20800 22060 20806
rect 22008 20742 22060 20748
rect 22020 20466 22048 20742
rect 22008 20460 22060 20466
rect 22008 20402 22060 20408
rect 21916 19372 21968 19378
rect 22020 19360 22048 20402
rect 22376 20256 22428 20262
rect 22376 20198 22428 20204
rect 22388 19922 22416 20198
rect 22376 19916 22428 19922
rect 22376 19858 22428 19864
rect 22192 19712 22244 19718
rect 22192 19654 22244 19660
rect 22100 19508 22152 19514
rect 22100 19450 22152 19456
rect 21968 19332 22048 19360
rect 21916 19314 21968 19320
rect 21916 19236 21968 19242
rect 21916 19178 21968 19184
rect 21928 18630 21956 19178
rect 22020 18698 22048 19332
rect 22112 18970 22140 19450
rect 22204 19378 22232 19654
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 22100 18964 22152 18970
rect 22100 18906 22152 18912
rect 22664 18834 22692 21830
rect 22652 18828 22704 18834
rect 22652 18770 22704 18776
rect 22008 18692 22060 18698
rect 22008 18634 22060 18640
rect 22468 18692 22520 18698
rect 22468 18634 22520 18640
rect 21916 18624 21968 18630
rect 21916 18566 21968 18572
rect 21548 18284 21600 18290
rect 21548 18226 21600 18232
rect 21560 16794 21588 18226
rect 21732 17604 21784 17610
rect 21732 17546 21784 17552
rect 21640 17332 21692 17338
rect 21640 17274 21692 17280
rect 21652 16794 21680 17274
rect 21744 17134 21772 17546
rect 21928 17338 21956 18566
rect 22098 17912 22154 17921
rect 22098 17847 22154 17856
rect 21916 17332 21968 17338
rect 21916 17274 21968 17280
rect 21732 17128 21784 17134
rect 21732 17070 21784 17076
rect 21824 17128 21876 17134
rect 21824 17070 21876 17076
rect 21548 16788 21600 16794
rect 21548 16730 21600 16736
rect 21640 16788 21692 16794
rect 21640 16730 21692 16736
rect 21454 16552 21510 16561
rect 21454 16487 21510 16496
rect 20812 15972 20864 15978
rect 20812 15914 20864 15920
rect 21088 15972 21140 15978
rect 21088 15914 21140 15920
rect 20352 15088 20404 15094
rect 20352 15030 20404 15036
rect 20536 15088 20588 15094
rect 20536 15030 20588 15036
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19982 14104 20038 14113
rect 20088 14074 20116 14214
rect 19982 14039 19984 14048
rect 20036 14039 20038 14048
rect 20076 14068 20128 14074
rect 19984 14010 20036 14016
rect 20076 14010 20128 14016
rect 19432 13728 19484 13734
rect 19432 13670 19484 13676
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 19536 13394 19564 13670
rect 19524 13388 19576 13394
rect 19524 13330 19576 13336
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 20548 12782 20576 15030
rect 20824 14906 20852 15914
rect 20904 15904 20956 15910
rect 20904 15846 20956 15852
rect 20916 15638 20944 15846
rect 21468 15638 21496 16487
rect 20904 15632 20956 15638
rect 20904 15574 20956 15580
rect 21456 15632 21508 15638
rect 21456 15574 21508 15580
rect 21088 15360 21140 15366
rect 21272 15360 21324 15366
rect 21088 15302 21140 15308
rect 21270 15328 21272 15337
rect 21324 15328 21326 15337
rect 20732 14878 20852 14906
rect 20996 14952 21048 14958
rect 20996 14894 21048 14900
rect 20628 14544 20680 14550
rect 20626 14512 20628 14521
rect 20680 14512 20682 14521
rect 20626 14447 20682 14456
rect 20628 13932 20680 13938
rect 20628 13874 20680 13880
rect 20168 12776 20220 12782
rect 20168 12718 20220 12724
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 19340 12368 19392 12374
rect 19340 12310 19392 12316
rect 18512 12164 18564 12170
rect 18512 12106 18564 12112
rect 18880 12164 18932 12170
rect 18880 12106 18932 12112
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 18616 11218 18644 11630
rect 18788 11620 18840 11626
rect 18788 11562 18840 11568
rect 18328 11212 18380 11218
rect 18328 11154 18380 11160
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 18144 10532 18196 10538
rect 18144 10474 18196 10480
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17500 9036 17552 9042
rect 17500 8978 17552 8984
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17512 8362 17540 8978
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 17500 8356 17552 8362
rect 17500 8298 17552 8304
rect 17604 8090 17632 8502
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17408 7472 17460 7478
rect 17408 7414 17460 7420
rect 17316 7268 17368 7274
rect 17316 7210 17368 7216
rect 17316 6928 17368 6934
rect 17316 6870 17368 6876
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17222 4584 17278 4593
rect 17222 4519 17224 4528
rect 17276 4519 17278 4528
rect 17224 4490 17276 4496
rect 17328 4146 17356 6870
rect 17420 5914 17448 7414
rect 17788 6769 17816 8910
rect 17972 8401 18000 9590
rect 18064 9450 18092 9590
rect 18052 9444 18104 9450
rect 18052 9386 18104 9392
rect 17958 8392 18014 8401
rect 17958 8327 18014 8336
rect 17960 8016 18012 8022
rect 17960 7958 18012 7964
rect 17972 7546 18000 7958
rect 18156 7818 18184 10474
rect 18234 9752 18290 9761
rect 18234 9687 18290 9696
rect 18144 7812 18196 7818
rect 18144 7754 18196 7760
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17774 6760 17830 6769
rect 17774 6695 17776 6704
rect 17828 6695 17830 6704
rect 17776 6666 17828 6672
rect 17788 6118 17816 6666
rect 17958 6352 18014 6361
rect 17958 6287 18014 6296
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17682 5808 17738 5817
rect 17682 5743 17738 5752
rect 17408 5296 17460 5302
rect 17408 5238 17460 5244
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17420 4078 17448 5238
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 17604 4146 17632 4558
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17408 4072 17460 4078
rect 17408 4014 17460 4020
rect 17500 3596 17552 3602
rect 17500 3538 17552 3544
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17420 2990 17448 3470
rect 17512 3058 17540 3538
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 17420 2446 17448 2926
rect 17604 2514 17632 4082
rect 17696 4078 17724 5743
rect 17788 5030 17816 6054
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 17684 4072 17736 4078
rect 17684 4014 17736 4020
rect 17788 3126 17816 4966
rect 17972 4214 18000 6287
rect 17960 4208 18012 4214
rect 17960 4150 18012 4156
rect 17866 4040 17922 4049
rect 17866 3975 17922 3984
rect 17880 3534 17908 3975
rect 18064 3942 18092 7686
rect 18248 6934 18276 9687
rect 18340 8090 18368 11018
rect 18512 10736 18564 10742
rect 18512 10678 18564 10684
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18432 10266 18460 10542
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18418 9888 18474 9897
rect 18418 9823 18474 9832
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 18236 6928 18288 6934
rect 18142 6896 18198 6905
rect 18236 6870 18288 6876
rect 18142 6831 18198 6840
rect 18156 6798 18184 6831
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 18340 5166 18368 7482
rect 18432 6866 18460 9823
rect 18524 9110 18552 10678
rect 18616 9761 18644 11154
rect 18800 10266 18828 11562
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 18892 10198 18920 12106
rect 19246 11248 19302 11257
rect 19246 11183 19302 11192
rect 19064 11076 19116 11082
rect 19064 11018 19116 11024
rect 19076 10742 19104 11018
rect 19064 10736 19116 10742
rect 19064 10678 19116 10684
rect 18880 10192 18932 10198
rect 18880 10134 18932 10140
rect 18602 9752 18658 9761
rect 18602 9687 18658 9696
rect 19156 9512 19208 9518
rect 19156 9454 19208 9460
rect 18512 9104 18564 9110
rect 18512 9046 18564 9052
rect 18604 9104 18656 9110
rect 18604 9046 18656 9052
rect 18616 8922 18644 9046
rect 18524 8906 18644 8922
rect 19168 8906 19196 9454
rect 19260 9450 19288 11183
rect 19352 10826 19380 12310
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19798 11792 19854 11801
rect 19798 11727 19800 11736
rect 19852 11727 19854 11736
rect 19800 11698 19852 11704
rect 19812 11121 19840 11698
rect 19996 11234 20024 12038
rect 20088 11558 20116 12582
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 19996 11206 20116 11234
rect 20180 11218 20208 12718
rect 20260 12708 20312 12714
rect 20260 12650 20312 12656
rect 20272 11898 20300 12650
rect 20640 12481 20668 13874
rect 20626 12472 20682 12481
rect 20626 12407 20682 12416
rect 20732 12306 20760 14878
rect 21008 14346 21036 14894
rect 21100 14346 21128 15302
rect 21270 15263 21326 15272
rect 21180 14884 21232 14890
rect 21180 14826 21232 14832
rect 20996 14340 21048 14346
rect 20996 14282 21048 14288
rect 21088 14340 21140 14346
rect 21088 14282 21140 14288
rect 20812 14000 20864 14006
rect 20812 13942 20864 13948
rect 20824 13394 20852 13942
rect 20904 13796 20956 13802
rect 20904 13738 20956 13744
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 20916 13258 20944 13738
rect 21192 13394 21220 14826
rect 21456 13524 21508 13530
rect 21456 13466 21508 13472
rect 21180 13388 21232 13394
rect 21180 13330 21232 13336
rect 20904 13252 20956 13258
rect 20904 13194 20956 13200
rect 21180 13184 21232 13190
rect 21180 13126 21232 13132
rect 20720 12300 20772 12306
rect 20720 12242 20772 12248
rect 21086 12200 21142 12209
rect 21192 12170 21220 13126
rect 21468 12918 21496 13466
rect 21456 12912 21508 12918
rect 21456 12854 21508 12860
rect 21560 12434 21588 16730
rect 21640 16108 21692 16114
rect 21640 16050 21692 16056
rect 21652 15570 21680 16050
rect 21640 15564 21692 15570
rect 21640 15506 21692 15512
rect 21652 14113 21680 15506
rect 21744 15366 21772 17070
rect 21732 15360 21784 15366
rect 21732 15302 21784 15308
rect 21732 14884 21784 14890
rect 21732 14826 21784 14832
rect 21744 14346 21772 14826
rect 21732 14340 21784 14346
rect 21732 14282 21784 14288
rect 21638 14104 21694 14113
rect 21638 14039 21694 14048
rect 21652 13938 21680 14039
rect 21640 13932 21692 13938
rect 21640 13874 21692 13880
rect 21836 12434 21864 17070
rect 21916 15632 21968 15638
rect 21916 15574 21968 15580
rect 21928 13394 21956 15574
rect 22112 15026 22140 17847
rect 22192 17264 22244 17270
rect 22192 17206 22244 17212
rect 22204 16522 22232 17206
rect 22284 16720 22336 16726
rect 22284 16662 22336 16668
rect 22192 16516 22244 16522
rect 22192 16458 22244 16464
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 22204 15162 22232 15438
rect 22192 15156 22244 15162
rect 22192 15098 22244 15104
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 22100 14612 22152 14618
rect 22100 14554 22152 14560
rect 22112 14414 22140 14554
rect 22296 14521 22324 16662
rect 22376 15360 22428 15366
rect 22376 15302 22428 15308
rect 22282 14512 22338 14521
rect 22282 14447 22338 14456
rect 22008 14408 22060 14414
rect 22006 14376 22008 14385
rect 22100 14408 22152 14414
rect 22060 14376 22062 14385
rect 22100 14350 22152 14356
rect 22006 14311 22062 14320
rect 22100 14272 22152 14278
rect 22100 14214 22152 14220
rect 21916 13388 21968 13394
rect 21916 13330 21968 13336
rect 21376 12406 21588 12434
rect 21744 12406 21864 12434
rect 21086 12135 21142 12144
rect 21180 12164 21232 12170
rect 20812 12096 20864 12102
rect 20812 12038 20864 12044
rect 20260 11892 20312 11898
rect 20260 11834 20312 11840
rect 20824 11830 20852 12038
rect 20812 11824 20864 11830
rect 20812 11766 20864 11772
rect 20996 11824 21048 11830
rect 20996 11766 21048 11772
rect 21008 11529 21036 11766
rect 20994 11520 21050 11529
rect 20994 11455 21050 11464
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 20812 11280 20864 11286
rect 21008 11257 21036 11290
rect 20812 11222 20864 11228
rect 20994 11248 21050 11257
rect 19798 11112 19854 11121
rect 20088 11082 20116 11206
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 19798 11047 19854 11056
rect 20076 11076 20128 11082
rect 20076 11018 20128 11024
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19352 10798 19472 10826
rect 19340 10736 19392 10742
rect 19340 10678 19392 10684
rect 19248 9444 19300 9450
rect 19248 9386 19300 9392
rect 18512 8900 18644 8906
rect 18564 8894 18644 8900
rect 18696 8900 18748 8906
rect 18512 8842 18564 8848
rect 18696 8842 18748 8848
rect 18788 8900 18840 8906
rect 18788 8842 18840 8848
rect 19156 8900 19208 8906
rect 19156 8842 19208 8848
rect 18708 8634 18736 8842
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 18512 8560 18564 8566
rect 18512 8502 18564 8508
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 18524 6633 18552 8502
rect 18616 8362 18644 8570
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18696 8016 18748 8022
rect 18696 7958 18748 7964
rect 18708 7886 18736 7958
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18510 6624 18566 6633
rect 18510 6559 18566 6568
rect 18708 6458 18736 7822
rect 18800 7546 18828 8842
rect 18970 8392 19026 8401
rect 18970 8327 19026 8336
rect 18880 8288 18932 8294
rect 18880 8230 18932 8236
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 18788 7200 18840 7206
rect 18788 7142 18840 7148
rect 18800 7002 18828 7142
rect 18788 6996 18840 7002
rect 18788 6938 18840 6944
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18604 5568 18656 5574
rect 18604 5510 18656 5516
rect 18328 5160 18380 5166
rect 18328 5102 18380 5108
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17776 3120 17828 3126
rect 17776 3062 17828 3068
rect 17880 2990 17908 3470
rect 18156 3466 18184 4966
rect 18616 4486 18644 5510
rect 18604 4480 18656 4486
rect 18604 4422 18656 4428
rect 18616 4214 18644 4422
rect 18604 4208 18656 4214
rect 18604 4150 18656 4156
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18524 3534 18552 4082
rect 18616 3942 18644 4150
rect 18800 4146 18828 6734
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 18604 3936 18656 3942
rect 18604 3878 18656 3884
rect 18616 3602 18644 3878
rect 18604 3596 18656 3602
rect 18604 3538 18656 3544
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18144 3460 18196 3466
rect 18144 3402 18196 3408
rect 18696 3460 18748 3466
rect 18696 3402 18748 3408
rect 17868 2984 17920 2990
rect 17868 2926 17920 2932
rect 17592 2508 17644 2514
rect 17592 2450 17644 2456
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 13544 2372 13596 2378
rect 13544 2314 13596 2320
rect 14556 2372 14608 2378
rect 14556 2314 14608 2320
rect 11888 1896 11940 1902
rect 11888 1838 11940 1844
rect 13556 800 13584 2314
rect 14568 2038 14596 2314
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 14556 2032 14608 2038
rect 14556 1974 14608 1980
rect 14844 800 14872 2246
rect 16776 800 16804 2246
rect 18708 800 18736 3402
rect 18892 3398 18920 8230
rect 18880 3392 18932 3398
rect 18880 3334 18932 3340
rect 18878 2680 18934 2689
rect 18878 2615 18934 2624
rect 18892 2446 18920 2615
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 18984 2310 19012 8327
rect 19168 7546 19196 8842
rect 19260 8498 19288 9386
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 19260 7478 19288 8434
rect 19352 8090 19380 10678
rect 19444 10305 19472 10798
rect 20076 10736 20128 10742
rect 20076 10678 20128 10684
rect 19616 10600 19668 10606
rect 19616 10542 19668 10548
rect 19430 10296 19486 10305
rect 19628 10266 19656 10542
rect 20088 10470 20116 10678
rect 20260 10668 20312 10674
rect 20260 10610 20312 10616
rect 20272 10470 20300 10610
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 20350 10432 20406 10441
rect 20350 10367 20406 10376
rect 19430 10231 19486 10240
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 20076 10056 20128 10062
rect 20076 9998 20128 10004
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19984 9648 20036 9654
rect 19982 9616 19984 9625
rect 20036 9616 20038 9625
rect 19982 9551 20038 9560
rect 19708 9376 19760 9382
rect 19708 9318 19760 9324
rect 19720 8906 19748 9318
rect 19708 8900 19760 8906
rect 19708 8842 19760 8848
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19892 8628 19944 8634
rect 19996 8616 20024 9551
rect 19944 8588 20024 8616
rect 19892 8570 19944 8576
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19248 7472 19300 7478
rect 19062 7440 19118 7449
rect 19248 7414 19300 7420
rect 19062 7375 19064 7384
rect 19116 7375 19118 7384
rect 19064 7346 19116 7352
rect 19076 5914 19104 7346
rect 19156 6928 19208 6934
rect 19156 6870 19208 6876
rect 19064 5908 19116 5914
rect 19064 5850 19116 5856
rect 19064 5636 19116 5642
rect 19064 5578 19116 5584
rect 19076 4049 19104 5578
rect 19168 4865 19196 6870
rect 19248 6792 19300 6798
rect 19246 6760 19248 6769
rect 19300 6760 19302 6769
rect 19246 6695 19302 6704
rect 19352 6118 19380 7822
rect 19444 6866 19472 8570
rect 20088 8242 20116 9998
rect 20166 8936 20222 8945
rect 20166 8871 20222 8880
rect 20180 8362 20208 8871
rect 20168 8356 20220 8362
rect 20168 8298 20220 8304
rect 20088 8214 20208 8242
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19996 7206 20024 7822
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 19984 7200 20036 7206
rect 19984 7142 20036 7148
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19708 6792 19760 6798
rect 19444 6740 19708 6746
rect 19444 6734 19760 6740
rect 19444 6718 19748 6734
rect 19444 6390 19472 6718
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19996 6458 20024 7142
rect 20088 6934 20116 7346
rect 20076 6928 20128 6934
rect 20076 6870 20128 6876
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 19432 6384 19484 6390
rect 19432 6326 19484 6332
rect 19524 6316 19576 6322
rect 19524 6258 19576 6264
rect 19628 6310 20116 6338
rect 19432 6180 19484 6186
rect 19432 6122 19484 6128
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19260 5914 19288 6054
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19246 5264 19302 5273
rect 19246 5199 19302 5208
rect 19260 5166 19288 5199
rect 19248 5160 19300 5166
rect 19248 5102 19300 5108
rect 19248 5024 19300 5030
rect 19248 4966 19300 4972
rect 19154 4856 19210 4865
rect 19154 4791 19210 4800
rect 19260 4486 19288 4966
rect 19352 4758 19380 5714
rect 19444 5250 19472 6122
rect 19536 6089 19564 6258
rect 19628 6254 19656 6310
rect 19616 6248 19668 6254
rect 19616 6190 19668 6196
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 20088 6202 20116 6310
rect 20180 6202 20208 8214
rect 20260 7744 20312 7750
rect 20258 7712 20260 7721
rect 20312 7712 20314 7721
rect 20258 7647 20314 7656
rect 20364 6905 20392 10367
rect 20732 10282 20760 10950
rect 20824 10606 20852 11222
rect 20994 11183 21050 11192
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 20548 10254 20760 10282
rect 20548 10198 20576 10254
rect 20536 10192 20588 10198
rect 20536 10134 20588 10140
rect 20626 10160 20682 10169
rect 20626 10095 20682 10104
rect 20812 10124 20864 10130
rect 20534 9888 20590 9897
rect 20534 9823 20590 9832
rect 20444 9648 20496 9654
rect 20444 9590 20496 9596
rect 20350 6896 20406 6905
rect 20260 6860 20312 6866
rect 20350 6831 20406 6840
rect 20260 6802 20312 6808
rect 20272 6769 20300 6802
rect 20258 6760 20314 6769
rect 20258 6695 20314 6704
rect 19616 6112 19668 6118
rect 19522 6080 19578 6089
rect 19616 6054 19668 6060
rect 19522 6015 19578 6024
rect 19628 5574 19656 6054
rect 19996 5658 20024 6190
rect 20088 6174 20300 6202
rect 20272 5710 20300 6174
rect 20168 5704 20220 5710
rect 19996 5630 20116 5658
rect 20168 5646 20220 5652
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 19616 5568 19668 5574
rect 19616 5510 19668 5516
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19444 5222 19564 5250
rect 19340 4752 19392 4758
rect 19340 4694 19392 4700
rect 19430 4720 19486 4729
rect 19430 4655 19486 4664
rect 19444 4622 19472 4655
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19248 4480 19300 4486
rect 19536 4468 19564 5222
rect 19892 5228 19944 5234
rect 19892 5170 19944 5176
rect 19904 5098 19932 5170
rect 19892 5092 19944 5098
rect 19892 5034 19944 5040
rect 19708 5024 19760 5030
rect 19708 4966 19760 4972
rect 19720 4758 19748 4966
rect 19708 4752 19760 4758
rect 19708 4694 19760 4700
rect 19248 4422 19300 4428
rect 19444 4440 19564 4468
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19062 4040 19118 4049
rect 19062 3975 19118 3984
rect 19156 3596 19208 3602
rect 19156 3538 19208 3544
rect 19064 3120 19116 3126
rect 19064 3062 19116 3068
rect 19076 2650 19104 3062
rect 19168 3058 19196 3538
rect 19156 3052 19208 3058
rect 19156 2994 19208 3000
rect 19260 2922 19288 4082
rect 19444 3398 19472 4440
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19996 3505 20024 5510
rect 20088 5098 20116 5630
rect 20076 5092 20128 5098
rect 20076 5034 20128 5040
rect 19982 3496 20038 3505
rect 19982 3431 19984 3440
rect 20036 3431 20038 3440
rect 19984 3402 20036 3408
rect 19432 3392 19484 3398
rect 19996 3371 20024 3402
rect 19432 3334 19484 3340
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19982 3088 20038 3097
rect 19982 3023 20038 3032
rect 19996 2990 20024 3023
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19248 2916 19300 2922
rect 19248 2858 19300 2864
rect 20088 2650 20116 5034
rect 20180 4486 20208 5646
rect 20364 4758 20392 6831
rect 20456 5681 20484 9590
rect 20548 9110 20576 9823
rect 20536 9104 20588 9110
rect 20536 9046 20588 9052
rect 20640 7886 20668 10095
rect 20812 10066 20864 10072
rect 20720 9988 20772 9994
rect 20720 9930 20772 9936
rect 20732 9518 20760 9930
rect 20720 9512 20772 9518
rect 20720 9454 20772 9460
rect 20718 8528 20774 8537
rect 20718 8463 20774 8472
rect 20732 8430 20760 8463
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20824 8022 20852 10066
rect 20996 9512 21048 9518
rect 20916 9472 20996 9500
rect 20916 8974 20944 9472
rect 20996 9454 21048 9460
rect 20904 8968 20956 8974
rect 20904 8910 20956 8916
rect 20916 8566 20944 8910
rect 20904 8560 20956 8566
rect 20904 8502 20956 8508
rect 20812 8016 20864 8022
rect 20812 7958 20864 7964
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20640 7342 20668 7822
rect 20812 7812 20864 7818
rect 20812 7754 20864 7760
rect 20904 7812 20956 7818
rect 20904 7754 20956 7760
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20628 5704 20680 5710
rect 20442 5672 20498 5681
rect 20628 5646 20680 5652
rect 20442 5607 20498 5616
rect 20640 5409 20668 5646
rect 20626 5400 20682 5409
rect 20626 5335 20682 5344
rect 20352 4752 20404 4758
rect 20352 4694 20404 4700
rect 20260 4684 20312 4690
rect 20260 4626 20312 4632
rect 20272 4554 20300 4626
rect 20260 4548 20312 4554
rect 20260 4490 20312 4496
rect 20168 4480 20220 4486
rect 20168 4422 20220 4428
rect 20732 4078 20760 6598
rect 20824 5545 20852 7754
rect 20916 7721 20944 7754
rect 20902 7712 20958 7721
rect 20902 7647 20958 7656
rect 20996 6180 21048 6186
rect 20996 6122 21048 6128
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 20916 5642 20944 5850
rect 20904 5636 20956 5642
rect 20904 5578 20956 5584
rect 20810 5536 20866 5545
rect 20810 5471 20866 5480
rect 20824 5166 20852 5471
rect 20812 5160 20864 5166
rect 20812 5102 20864 5108
rect 21008 4672 21036 6122
rect 20916 4644 21036 4672
rect 20916 4554 20944 4644
rect 21100 4570 21128 12135
rect 21180 12106 21232 12112
rect 21376 9674 21404 12406
rect 21456 11620 21508 11626
rect 21456 11562 21508 11568
rect 21468 11150 21496 11562
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 21640 11076 21692 11082
rect 21640 11018 21692 11024
rect 21548 10804 21600 10810
rect 21548 10746 21600 10752
rect 21560 10713 21588 10746
rect 21546 10704 21602 10713
rect 21546 10639 21602 10648
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 21560 9722 21588 10542
rect 21284 9646 21404 9674
rect 21548 9716 21600 9722
rect 21548 9658 21600 9664
rect 21284 8537 21312 9646
rect 21270 8528 21326 8537
rect 21270 8463 21326 8472
rect 21180 8424 21232 8430
rect 21180 8366 21232 8372
rect 21456 8424 21508 8430
rect 21456 8366 21508 8372
rect 21192 8129 21220 8366
rect 21362 8256 21418 8265
rect 21362 8191 21418 8200
rect 21178 8120 21234 8129
rect 21178 8055 21234 8064
rect 21192 5914 21220 8055
rect 21376 7954 21404 8191
rect 21364 7948 21416 7954
rect 21364 7890 21416 7896
rect 21180 5908 21232 5914
rect 21180 5850 21232 5856
rect 20904 4548 20956 4554
rect 20904 4490 20956 4496
rect 21008 4542 21128 4570
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 20904 3460 20956 3466
rect 20904 3402 20956 3408
rect 20916 3233 20944 3402
rect 20902 3224 20958 3233
rect 20902 3159 20958 3168
rect 20260 3120 20312 3126
rect 21008 3074 21036 4542
rect 21086 4448 21142 4457
rect 21086 4383 21142 4392
rect 20312 3068 21036 3074
rect 20260 3062 21036 3068
rect 20272 3046 21036 3062
rect 21100 3058 21128 4383
rect 21178 3632 21234 3641
rect 21178 3567 21234 3576
rect 21192 3398 21220 3567
rect 21180 3392 21232 3398
rect 21180 3334 21232 3340
rect 21376 3194 21404 7890
rect 21468 7410 21496 8366
rect 21652 8090 21680 11018
rect 21744 11014 21772 12406
rect 21928 12374 21956 13330
rect 21916 12368 21968 12374
rect 21916 12310 21968 12316
rect 22008 11892 22060 11898
rect 22008 11834 22060 11840
rect 22020 11778 22048 11834
rect 22112 11830 22140 14214
rect 22296 13841 22324 14447
rect 22282 13832 22338 13841
rect 22282 13767 22338 13776
rect 21928 11750 22048 11778
rect 22100 11824 22152 11830
rect 22100 11766 22152 11772
rect 21824 11688 21876 11694
rect 21824 11630 21876 11636
rect 21732 11008 21784 11014
rect 21732 10950 21784 10956
rect 21744 9042 21772 10950
rect 21836 10266 21864 11630
rect 21928 11558 21956 11750
rect 21916 11552 21968 11558
rect 21916 11494 21968 11500
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 22020 11218 22048 11494
rect 22008 11212 22060 11218
rect 22008 11154 22060 11160
rect 22098 10976 22154 10985
rect 22098 10911 22154 10920
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 21914 10296 21970 10305
rect 21824 10260 21876 10266
rect 21914 10231 21970 10240
rect 21824 10202 21876 10208
rect 21928 10198 21956 10231
rect 21916 10192 21968 10198
rect 21916 10134 21968 10140
rect 22020 10146 22048 10610
rect 22112 10470 22140 10911
rect 22190 10704 22246 10713
rect 22190 10639 22246 10648
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22204 10266 22232 10639
rect 22296 10470 22324 13767
rect 22284 10464 22336 10470
rect 22284 10406 22336 10412
rect 22388 10282 22416 15302
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 22296 10254 22416 10282
rect 21824 10124 21876 10130
rect 21824 10066 21876 10072
rect 22020 10118 22140 10146
rect 21836 9761 21864 10066
rect 21916 10056 21968 10062
rect 21914 10024 21916 10033
rect 21968 10024 21970 10033
rect 21914 9959 21970 9968
rect 21822 9752 21878 9761
rect 21822 9687 21878 9696
rect 21916 9648 21968 9654
rect 21916 9590 21968 9596
rect 21928 9353 21956 9590
rect 22020 9518 22048 10118
rect 22008 9512 22060 9518
rect 22112 9500 22140 10118
rect 22192 10124 22244 10130
rect 22192 10066 22244 10072
rect 22204 9926 22232 10066
rect 22192 9920 22244 9926
rect 22192 9862 22244 9868
rect 22296 9602 22324 10254
rect 22480 9738 22508 18634
rect 22664 18358 22692 18770
rect 22744 18692 22796 18698
rect 22744 18634 22796 18640
rect 22652 18352 22704 18358
rect 22652 18294 22704 18300
rect 22652 18216 22704 18222
rect 22652 18158 22704 18164
rect 22664 17610 22692 18158
rect 22756 17882 22784 18634
rect 22848 18222 22876 22918
rect 22836 18216 22888 18222
rect 22836 18158 22888 18164
rect 22744 17876 22796 17882
rect 22744 17818 22796 17824
rect 22652 17604 22704 17610
rect 22652 17546 22704 17552
rect 22560 16992 22612 16998
rect 22560 16934 22612 16940
rect 22572 16046 22600 16934
rect 22940 16454 22968 27814
rect 23124 22094 23152 28358
rect 23676 26926 23704 29446
rect 24768 28008 24820 28014
rect 24768 27950 24820 27956
rect 23664 26920 23716 26926
rect 23664 26862 23716 26868
rect 23676 23322 23704 26862
rect 23664 23316 23716 23322
rect 23664 23258 23716 23264
rect 23676 23118 23704 23258
rect 23664 23112 23716 23118
rect 23664 23054 23716 23060
rect 23032 22066 23152 22094
rect 22928 16448 22980 16454
rect 22928 16390 22980 16396
rect 22560 16040 22612 16046
rect 22560 15982 22612 15988
rect 22652 15156 22704 15162
rect 22652 15098 22704 15104
rect 22664 12434 22692 15098
rect 22928 14884 22980 14890
rect 22928 14826 22980 14832
rect 22744 13728 22796 13734
rect 22744 13670 22796 13676
rect 22756 12986 22784 13670
rect 22940 13462 22968 14826
rect 23032 13462 23060 22066
rect 23112 20460 23164 20466
rect 23112 20402 23164 20408
rect 23124 19990 23152 20402
rect 24780 19990 24808 27950
rect 24860 27940 24912 27946
rect 24860 27882 24912 27888
rect 24872 20466 24900 27882
rect 24952 20936 25004 20942
rect 24952 20878 25004 20884
rect 24964 20466 24992 20878
rect 25424 20806 25452 37062
rect 25688 33516 25740 33522
rect 25688 33458 25740 33464
rect 25596 29028 25648 29034
rect 25596 28970 25648 28976
rect 25608 28218 25636 28970
rect 25596 28212 25648 28218
rect 25596 28154 25648 28160
rect 25608 22098 25636 28154
rect 25596 22092 25648 22098
rect 25596 22034 25648 22040
rect 25700 21690 25728 33458
rect 26344 28218 26372 37130
rect 27080 37126 27108 39200
rect 27160 37256 27212 37262
rect 27160 37198 27212 37204
rect 27344 37256 27396 37262
rect 27344 37198 27396 37204
rect 27068 37120 27120 37126
rect 27068 37062 27120 37068
rect 26976 30728 27028 30734
rect 26976 30670 27028 30676
rect 26332 28212 26384 28218
rect 26332 28154 26384 28160
rect 26424 27328 26476 27334
rect 26424 27270 26476 27276
rect 25688 21684 25740 21690
rect 25688 21626 25740 21632
rect 25136 20800 25188 20806
rect 25136 20742 25188 20748
rect 25412 20800 25464 20806
rect 25412 20742 25464 20748
rect 24860 20460 24912 20466
rect 24860 20402 24912 20408
rect 24952 20460 25004 20466
rect 24952 20402 25004 20408
rect 24860 20256 24912 20262
rect 24860 20198 24912 20204
rect 23112 19984 23164 19990
rect 23112 19926 23164 19932
rect 24768 19984 24820 19990
rect 24768 19926 24820 19932
rect 23124 19718 23152 19926
rect 23756 19848 23808 19854
rect 23756 19790 23808 19796
rect 23112 19712 23164 19718
rect 23112 19654 23164 19660
rect 23124 17882 23152 19654
rect 23768 18834 23796 19790
rect 24032 19712 24084 19718
rect 24032 19654 24084 19660
rect 24676 19712 24728 19718
rect 24676 19654 24728 19660
rect 24044 19446 24072 19654
rect 24032 19440 24084 19446
rect 24032 19382 24084 19388
rect 24308 19372 24360 19378
rect 24308 19314 24360 19320
rect 23756 18828 23808 18834
rect 23756 18770 23808 18776
rect 23296 18692 23348 18698
rect 23296 18634 23348 18640
rect 23112 17876 23164 17882
rect 23112 17818 23164 17824
rect 23308 16182 23336 18634
rect 23388 18352 23440 18358
rect 23388 18294 23440 18300
rect 23400 17338 23428 18294
rect 24032 18216 24084 18222
rect 24032 18158 24084 18164
rect 23570 17368 23626 17377
rect 23388 17332 23440 17338
rect 23570 17303 23626 17312
rect 23388 17274 23440 17280
rect 23480 16992 23532 16998
rect 23480 16934 23532 16940
rect 23296 16176 23348 16182
rect 23296 16118 23348 16124
rect 23112 15632 23164 15638
rect 23308 15586 23336 16118
rect 23112 15574 23164 15580
rect 23124 14550 23152 15574
rect 23216 15558 23336 15586
rect 23112 14544 23164 14550
rect 23112 14486 23164 14492
rect 22928 13456 22980 13462
rect 22928 13398 22980 13404
rect 23020 13456 23072 13462
rect 23020 13398 23072 13404
rect 22744 12980 22796 12986
rect 22744 12922 22796 12928
rect 23032 12782 23060 13398
rect 23124 13394 23152 14486
rect 23216 14278 23244 15558
rect 23296 15496 23348 15502
rect 23296 15438 23348 15444
rect 23308 14618 23336 15438
rect 23492 15094 23520 16934
rect 23584 16658 23612 17303
rect 23572 16652 23624 16658
rect 23572 16594 23624 16600
rect 23756 16652 23808 16658
rect 23756 16594 23808 16600
rect 23664 16584 23716 16590
rect 23664 16526 23716 16532
rect 23676 15502 23704 16526
rect 23768 16454 23796 16594
rect 23756 16448 23808 16454
rect 23756 16390 23808 16396
rect 23848 16176 23900 16182
rect 23848 16118 23900 16124
rect 23860 15706 23888 16118
rect 24044 16046 24072 18158
rect 24216 17808 24268 17814
rect 24216 17750 24268 17756
rect 24124 16720 24176 16726
rect 24124 16662 24176 16668
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 23848 15700 23900 15706
rect 23848 15642 23900 15648
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23480 15088 23532 15094
rect 23480 15030 23532 15036
rect 23296 14612 23348 14618
rect 23296 14554 23348 14560
rect 23204 14272 23256 14278
rect 23204 14214 23256 14220
rect 23492 14074 23520 15030
rect 23572 14816 23624 14822
rect 23572 14758 23624 14764
rect 23584 14482 23612 14758
rect 23676 14618 23704 15438
rect 24136 14890 24164 16662
rect 24124 14884 24176 14890
rect 24124 14826 24176 14832
rect 23756 14816 23808 14822
rect 23756 14758 23808 14764
rect 23664 14612 23716 14618
rect 23664 14554 23716 14560
rect 23572 14476 23624 14482
rect 23572 14418 23624 14424
rect 23768 14414 23796 14758
rect 23940 14544 23992 14550
rect 23940 14486 23992 14492
rect 23756 14408 23808 14414
rect 23756 14350 23808 14356
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23848 14000 23900 14006
rect 23294 13968 23350 13977
rect 23848 13942 23900 13948
rect 23294 13903 23296 13912
rect 23348 13903 23350 13912
rect 23296 13874 23348 13880
rect 23480 13864 23532 13870
rect 23480 13806 23532 13812
rect 23756 13864 23808 13870
rect 23756 13806 23808 13812
rect 23388 13796 23440 13802
rect 23388 13738 23440 13744
rect 23112 13388 23164 13394
rect 23112 13330 23164 13336
rect 23296 13388 23348 13394
rect 23296 13330 23348 13336
rect 23204 13252 23256 13258
rect 23204 13194 23256 13200
rect 23216 12986 23244 13194
rect 23204 12980 23256 12986
rect 23204 12922 23256 12928
rect 23020 12776 23072 12782
rect 23020 12718 23072 12724
rect 23032 12434 23060 12718
rect 22664 12406 22784 12434
rect 23032 12406 23152 12434
rect 22652 11076 22704 11082
rect 22652 11018 22704 11024
rect 22560 10736 22612 10742
rect 22560 10678 22612 10684
rect 22572 10198 22600 10678
rect 22664 10606 22692 11018
rect 22652 10600 22704 10606
rect 22652 10542 22704 10548
rect 22652 10464 22704 10470
rect 22652 10406 22704 10412
rect 22560 10192 22612 10198
rect 22560 10134 22612 10140
rect 22480 9710 22600 9738
rect 22572 9625 22600 9710
rect 22558 9616 22614 9625
rect 22296 9574 22508 9602
rect 22284 9512 22336 9518
rect 22112 9472 22284 9500
rect 22008 9454 22060 9460
rect 22284 9454 22336 9460
rect 21914 9344 21970 9353
rect 21914 9279 21970 9288
rect 21732 9036 21784 9042
rect 21732 8978 21784 8984
rect 21640 8084 21692 8090
rect 21640 8026 21692 8032
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 21652 6322 21680 7346
rect 21744 7290 21772 8978
rect 22020 8634 22048 9454
rect 22100 9376 22152 9382
rect 22100 9318 22152 9324
rect 22112 9217 22140 9318
rect 22098 9208 22154 9217
rect 22098 9143 22154 9152
rect 22192 9036 22244 9042
rect 22192 8978 22244 8984
rect 22098 8664 22154 8673
rect 22008 8628 22060 8634
rect 22098 8599 22154 8608
rect 22008 8570 22060 8576
rect 22006 8528 22062 8537
rect 22006 8463 22062 8472
rect 22020 8430 22048 8463
rect 22008 8424 22060 8430
rect 21822 8392 21878 8401
rect 22008 8366 22060 8372
rect 22112 8362 22140 8599
rect 21822 8327 21824 8336
rect 21876 8327 21878 8336
rect 22100 8356 22152 8362
rect 21824 8298 21876 8304
rect 22100 8298 22152 8304
rect 22204 7478 22232 8978
rect 22480 8650 22508 9574
rect 22558 9551 22614 9560
rect 22388 8622 22508 8650
rect 22388 7834 22416 8622
rect 22388 7818 22508 7834
rect 22388 7812 22520 7818
rect 22388 7806 22468 7812
rect 22468 7754 22520 7760
rect 22192 7472 22244 7478
rect 22192 7414 22244 7420
rect 22376 7336 22428 7342
rect 21744 7262 21864 7290
rect 22376 7278 22428 7284
rect 21730 7168 21786 7177
rect 21730 7103 21786 7112
rect 21744 6866 21772 7103
rect 21732 6860 21784 6866
rect 21732 6802 21784 6808
rect 21732 6384 21784 6390
rect 21732 6326 21784 6332
rect 21640 6316 21692 6322
rect 21640 6258 21692 6264
rect 21548 6180 21600 6186
rect 21548 6122 21600 6128
rect 21560 5914 21588 6122
rect 21652 6118 21680 6258
rect 21744 6225 21772 6326
rect 21730 6216 21786 6225
rect 21730 6151 21786 6160
rect 21836 6118 21864 7262
rect 21916 7200 21968 7206
rect 22100 7200 22152 7206
rect 21916 7142 21968 7148
rect 22098 7168 22100 7177
rect 22152 7168 22154 7177
rect 21928 7041 21956 7142
rect 22098 7103 22154 7112
rect 22388 7041 22416 7278
rect 21914 7032 21970 7041
rect 21914 6967 21970 6976
rect 22374 7032 22430 7041
rect 22374 6967 22430 6976
rect 22376 6928 22428 6934
rect 22376 6870 22428 6876
rect 22192 6724 22244 6730
rect 22192 6666 22244 6672
rect 21916 6656 21968 6662
rect 21916 6598 21968 6604
rect 21640 6112 21692 6118
rect 21640 6054 21692 6060
rect 21824 6112 21876 6118
rect 21824 6054 21876 6060
rect 21548 5908 21600 5914
rect 21548 5850 21600 5856
rect 21456 5704 21508 5710
rect 21456 5646 21508 5652
rect 21468 5370 21496 5646
rect 21836 5574 21864 6054
rect 21928 5953 21956 6598
rect 22204 6186 22232 6666
rect 22388 6662 22416 6870
rect 22572 6866 22600 9551
rect 22664 7206 22692 10406
rect 22756 10266 22784 12406
rect 22928 12368 22980 12374
rect 22928 12310 22980 12316
rect 22836 11280 22888 11286
rect 22834 11248 22836 11257
rect 22888 11248 22890 11257
rect 22834 11183 22890 11192
rect 22836 10736 22888 10742
rect 22836 10678 22888 10684
rect 22848 10577 22876 10678
rect 22834 10568 22890 10577
rect 22834 10503 22890 10512
rect 22744 10260 22796 10266
rect 22744 10202 22796 10208
rect 22940 9897 22968 12310
rect 23124 12306 23152 12406
rect 23112 12300 23164 12306
rect 23112 12242 23164 12248
rect 23308 11898 23336 13330
rect 23400 12782 23428 13738
rect 23492 12918 23520 13806
rect 23480 12912 23532 12918
rect 23480 12854 23532 12860
rect 23388 12776 23440 12782
rect 23388 12718 23440 12724
rect 23296 11892 23348 11898
rect 23296 11834 23348 11840
rect 23492 11286 23520 12854
rect 23768 12434 23796 13806
rect 23676 12406 23796 12434
rect 23572 12300 23624 12306
rect 23572 12242 23624 12248
rect 23584 12102 23612 12242
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23480 11280 23532 11286
rect 23480 11222 23532 11228
rect 23478 11112 23534 11121
rect 23204 11076 23256 11082
rect 23478 11047 23534 11056
rect 23204 11018 23256 11024
rect 23112 10260 23164 10266
rect 23112 10202 23164 10208
rect 22926 9888 22982 9897
rect 22926 9823 22982 9832
rect 22742 9752 22798 9761
rect 22742 9687 22798 9696
rect 22652 7200 22704 7206
rect 22652 7142 22704 7148
rect 22560 6860 22612 6866
rect 22560 6802 22612 6808
rect 22468 6792 22520 6798
rect 22468 6734 22520 6740
rect 22376 6656 22428 6662
rect 22376 6598 22428 6604
rect 22480 6322 22508 6734
rect 22756 6662 22784 9687
rect 23124 9042 23152 10202
rect 23112 9036 23164 9042
rect 23112 8978 23164 8984
rect 23110 8800 23166 8809
rect 23110 8735 23166 8744
rect 22926 8120 22982 8129
rect 22926 8055 22982 8064
rect 22940 7546 22968 8055
rect 23124 7818 23152 8735
rect 23112 7812 23164 7818
rect 23112 7754 23164 7760
rect 22928 7540 22980 7546
rect 22928 7482 22980 7488
rect 22744 6656 22796 6662
rect 22744 6598 22796 6604
rect 22468 6316 22520 6322
rect 22468 6258 22520 6264
rect 22192 6180 22244 6186
rect 22192 6122 22244 6128
rect 22374 6080 22430 6089
rect 22374 6015 22430 6024
rect 21914 5944 21970 5953
rect 21914 5879 21970 5888
rect 22098 5944 22154 5953
rect 22098 5879 22100 5888
rect 22152 5879 22154 5888
rect 22100 5850 22152 5856
rect 21824 5568 21876 5574
rect 21824 5510 21876 5516
rect 22190 5400 22246 5409
rect 21456 5364 21508 5370
rect 22190 5335 22246 5344
rect 21456 5306 21508 5312
rect 21468 5234 21496 5306
rect 22204 5302 22232 5335
rect 22192 5296 22244 5302
rect 21638 5264 21694 5273
rect 21456 5228 21508 5234
rect 22192 5238 22244 5244
rect 21638 5199 21694 5208
rect 21456 5170 21508 5176
rect 21468 4690 21496 5170
rect 21652 5166 21680 5199
rect 21640 5160 21692 5166
rect 21640 5102 21692 5108
rect 22192 5160 22244 5166
rect 22192 5102 22244 5108
rect 22204 5030 22232 5102
rect 22192 5024 22244 5030
rect 22192 4966 22244 4972
rect 22388 4758 22416 6015
rect 22468 5364 22520 5370
rect 22468 5306 22520 5312
rect 22480 5030 22508 5306
rect 23124 5302 23152 7754
rect 23216 7750 23244 11018
rect 23388 8968 23440 8974
rect 23388 8910 23440 8916
rect 23400 8129 23428 8910
rect 23386 8120 23442 8129
rect 23386 8055 23442 8064
rect 23204 7744 23256 7750
rect 23204 7686 23256 7692
rect 23388 7744 23440 7750
rect 23388 7686 23440 7692
rect 23400 7206 23428 7686
rect 23388 7200 23440 7206
rect 23388 7142 23440 7148
rect 23296 6996 23348 7002
rect 23296 6938 23348 6944
rect 23204 6384 23256 6390
rect 23204 6326 23256 6332
rect 23112 5296 23164 5302
rect 23112 5238 23164 5244
rect 23216 5234 23244 6326
rect 23308 5846 23336 6938
rect 23296 5840 23348 5846
rect 23296 5782 23348 5788
rect 23204 5228 23256 5234
rect 23204 5170 23256 5176
rect 22560 5092 22612 5098
rect 22560 5034 22612 5040
rect 22468 5024 22520 5030
rect 22468 4966 22520 4972
rect 22376 4752 22428 4758
rect 22428 4712 22508 4740
rect 22376 4694 22428 4700
rect 21456 4684 21508 4690
rect 21456 4626 21508 4632
rect 21640 4548 21692 4554
rect 21640 4490 21692 4496
rect 21548 3596 21600 3602
rect 21548 3538 21600 3544
rect 21272 3188 21324 3194
rect 21272 3130 21324 3136
rect 21364 3188 21416 3194
rect 21364 3130 21416 3136
rect 21008 2650 21036 3046
rect 21088 3052 21140 3058
rect 21088 2994 21140 3000
rect 21284 2990 21312 3130
rect 21272 2984 21324 2990
rect 21272 2926 21324 2932
rect 21362 2952 21418 2961
rect 21362 2887 21418 2896
rect 21376 2854 21404 2887
rect 21560 2854 21588 3538
rect 21364 2848 21416 2854
rect 21364 2790 21416 2796
rect 21548 2848 21600 2854
rect 21548 2790 21600 2796
rect 19064 2644 19116 2650
rect 19064 2586 19116 2592
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 20996 2644 21048 2650
rect 20996 2586 21048 2592
rect 18972 2304 19024 2310
rect 18972 2246 19024 2252
rect 19076 1834 19104 2586
rect 19984 2576 20036 2582
rect 19984 2518 20036 2524
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19064 1828 19116 1834
rect 19064 1770 19116 1776
rect 19996 800 20024 2518
rect 20626 2408 20682 2417
rect 20626 2343 20628 2352
rect 20680 2343 20682 2352
rect 20628 2314 20680 2320
rect 21652 1970 21680 4490
rect 21824 4208 21876 4214
rect 21824 4150 21876 4156
rect 21836 2106 21864 4150
rect 22008 4140 22060 4146
rect 22008 4082 22060 4088
rect 21916 3664 21968 3670
rect 21916 3606 21968 3612
rect 21824 2100 21876 2106
rect 21824 2042 21876 2048
rect 21640 1964 21692 1970
rect 21640 1906 21692 1912
rect 21928 800 21956 3606
rect 22020 3058 22048 4082
rect 22376 4072 22428 4078
rect 22374 4040 22376 4049
rect 22428 4040 22430 4049
rect 22374 3975 22430 3984
rect 22480 3942 22508 4712
rect 22100 3936 22152 3942
rect 22098 3904 22100 3913
rect 22468 3936 22520 3942
rect 22152 3904 22154 3913
rect 22468 3878 22520 3884
rect 22098 3839 22154 3848
rect 22100 3732 22152 3738
rect 22100 3674 22152 3680
rect 22112 3641 22140 3674
rect 22098 3632 22154 3641
rect 22098 3567 22154 3576
rect 22572 3466 22600 5034
rect 23020 5024 23072 5030
rect 22926 4992 22982 5001
rect 23020 4966 23072 4972
rect 22926 4927 22982 4936
rect 22836 4820 22888 4826
rect 22836 4762 22888 4768
rect 22848 4554 22876 4762
rect 22836 4548 22888 4554
rect 22836 4490 22888 4496
rect 22940 3602 22968 4927
rect 23032 4826 23060 4966
rect 23020 4820 23072 4826
rect 23020 4762 23072 4768
rect 23020 4616 23072 4622
rect 23020 4558 23072 4564
rect 23032 3738 23060 4558
rect 23202 4040 23258 4049
rect 23202 3975 23258 3984
rect 23216 3738 23244 3975
rect 23020 3732 23072 3738
rect 23020 3674 23072 3680
rect 23204 3732 23256 3738
rect 23204 3674 23256 3680
rect 22928 3596 22980 3602
rect 22928 3538 22980 3544
rect 22192 3460 22244 3466
rect 22192 3402 22244 3408
rect 22560 3460 22612 3466
rect 22560 3402 22612 3408
rect 22204 3369 22232 3402
rect 22190 3360 22246 3369
rect 22190 3295 22246 3304
rect 22190 3224 22246 3233
rect 22190 3159 22192 3168
rect 22244 3159 22246 3168
rect 22192 3130 22244 3136
rect 22008 3052 22060 3058
rect 22008 2994 22060 3000
rect 22020 2514 22048 2994
rect 23308 2774 23336 5782
rect 23492 4865 23520 11047
rect 23676 10826 23704 12406
rect 23756 12164 23808 12170
rect 23756 12106 23808 12112
rect 23768 11665 23796 12106
rect 23754 11656 23810 11665
rect 23754 11591 23810 11600
rect 23860 11354 23888 13942
rect 23952 11830 23980 14486
rect 24136 14113 24164 14826
rect 24122 14104 24178 14113
rect 24122 14039 24178 14048
rect 24136 13530 24164 14039
rect 24124 13524 24176 13530
rect 24124 13466 24176 13472
rect 24030 13424 24086 13433
rect 24030 13359 24086 13368
rect 23940 11824 23992 11830
rect 23940 11766 23992 11772
rect 23848 11348 23900 11354
rect 23848 11290 23900 11296
rect 23756 11144 23808 11150
rect 23756 11086 23808 11092
rect 23584 10798 23704 10826
rect 23584 9489 23612 10798
rect 23664 10736 23716 10742
rect 23664 10678 23716 10684
rect 23570 9480 23626 9489
rect 23570 9415 23626 9424
rect 23676 9178 23704 10678
rect 23664 9172 23716 9178
rect 23664 9114 23716 9120
rect 23664 9036 23716 9042
rect 23664 8978 23716 8984
rect 23676 8838 23704 8978
rect 23768 8838 23796 11086
rect 24044 10062 24072 13359
rect 24124 12436 24176 12442
rect 24124 12378 24176 12384
rect 24136 10538 24164 12378
rect 24228 11121 24256 17750
rect 24320 17678 24348 19314
rect 24492 18080 24544 18086
rect 24492 18022 24544 18028
rect 24504 17746 24532 18022
rect 24492 17740 24544 17746
rect 24492 17682 24544 17688
rect 24308 17672 24360 17678
rect 24308 17614 24360 17620
rect 24584 17264 24636 17270
rect 24584 17206 24636 17212
rect 24308 16992 24360 16998
rect 24308 16934 24360 16940
rect 24320 14482 24348 16934
rect 24400 16448 24452 16454
rect 24400 16390 24452 16396
rect 24412 16250 24440 16390
rect 24400 16244 24452 16250
rect 24400 16186 24452 16192
rect 24308 14476 24360 14482
rect 24308 14418 24360 14424
rect 24320 12434 24348 14418
rect 24596 14414 24624 17206
rect 24584 14408 24636 14414
rect 24584 14350 24636 14356
rect 24492 12436 24544 12442
rect 24320 12406 24440 12434
rect 24308 11824 24360 11830
rect 24308 11766 24360 11772
rect 24214 11112 24270 11121
rect 24214 11047 24270 11056
rect 24124 10532 24176 10538
rect 24124 10474 24176 10480
rect 24032 10056 24084 10062
rect 24032 9998 24084 10004
rect 23848 9648 23900 9654
rect 23848 9590 23900 9596
rect 23664 8832 23716 8838
rect 23664 8774 23716 8780
rect 23756 8832 23808 8838
rect 23756 8774 23808 8780
rect 23768 8673 23796 8774
rect 23754 8664 23810 8673
rect 23754 8599 23810 8608
rect 23572 7812 23624 7818
rect 23572 7754 23624 7760
rect 23478 4856 23534 4865
rect 23478 4791 23534 4800
rect 23386 3088 23442 3097
rect 23386 3023 23388 3032
rect 23440 3023 23442 3032
rect 23388 2994 23440 3000
rect 23584 2922 23612 7754
rect 23756 6112 23808 6118
rect 23756 6054 23808 6060
rect 23768 5914 23796 6054
rect 23664 5908 23716 5914
rect 23664 5850 23716 5856
rect 23756 5908 23808 5914
rect 23756 5850 23808 5856
rect 23676 4010 23704 5850
rect 23860 5574 23888 9590
rect 24044 9382 24072 9998
rect 24228 9654 24256 11047
rect 24320 10198 24348 11766
rect 24308 10192 24360 10198
rect 24308 10134 24360 10140
rect 24216 9648 24268 9654
rect 24216 9590 24268 9596
rect 24124 9580 24176 9586
rect 24124 9522 24176 9528
rect 24032 9376 24084 9382
rect 24032 9318 24084 9324
rect 23940 8900 23992 8906
rect 23940 8842 23992 8848
rect 23952 6186 23980 8842
rect 24044 8430 24072 9318
rect 24032 8424 24084 8430
rect 24032 8366 24084 8372
rect 24136 7313 24164 9522
rect 24308 9512 24360 9518
rect 24308 9454 24360 9460
rect 24216 9104 24268 9110
rect 24216 9046 24268 9052
rect 24122 7304 24178 7313
rect 24122 7239 24178 7248
rect 24228 6458 24256 9046
rect 24320 8945 24348 9454
rect 24306 8936 24362 8945
rect 24412 8906 24440 12406
rect 24492 12378 24544 12384
rect 24504 11898 24532 12378
rect 24596 12306 24624 14350
rect 24688 12434 24716 19654
rect 24780 19310 24808 19926
rect 24768 19304 24820 19310
rect 24768 19246 24820 19252
rect 24780 17134 24808 19246
rect 24872 18902 24900 20198
rect 25148 19310 25176 20742
rect 26148 20460 26200 20466
rect 26148 20402 26200 20408
rect 26056 20392 26108 20398
rect 26056 20334 26108 20340
rect 25228 20256 25280 20262
rect 25228 20198 25280 20204
rect 25136 19304 25188 19310
rect 25136 19246 25188 19252
rect 24860 18896 24912 18902
rect 24860 18838 24912 18844
rect 25240 18834 25268 20198
rect 26068 20058 26096 20334
rect 26056 20052 26108 20058
rect 26056 19994 26108 20000
rect 26160 19854 26188 20402
rect 26148 19848 26200 19854
rect 26148 19790 26200 19796
rect 25780 19304 25832 19310
rect 25780 19246 25832 19252
rect 25228 18828 25280 18834
rect 25228 18770 25280 18776
rect 25136 18692 25188 18698
rect 25136 18634 25188 18640
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24964 17134 24992 18566
rect 24768 17128 24820 17134
rect 24768 17070 24820 17076
rect 24952 17128 25004 17134
rect 24952 17070 25004 17076
rect 24768 16992 24820 16998
rect 24768 16934 24820 16940
rect 24860 16992 24912 16998
rect 24860 16934 24912 16940
rect 24780 16794 24808 16934
rect 24768 16788 24820 16794
rect 24768 16730 24820 16736
rect 24872 16522 24900 16934
rect 24860 16516 24912 16522
rect 24860 16458 24912 16464
rect 24964 16266 24992 17070
rect 25148 16402 25176 18634
rect 25596 17604 25648 17610
rect 25596 17546 25648 17552
rect 25504 17128 25556 17134
rect 25504 17070 25556 17076
rect 24780 16250 24992 16266
rect 24768 16244 24992 16250
rect 24820 16238 24992 16244
rect 24768 16186 24820 16192
rect 24964 15094 24992 16238
rect 25056 16374 25176 16402
rect 24952 15088 25004 15094
rect 24952 15030 25004 15036
rect 24860 15020 24912 15026
rect 24860 14962 24912 14968
rect 24872 13734 24900 14962
rect 25056 14958 25084 16374
rect 25412 16176 25464 16182
rect 25412 16118 25464 16124
rect 25424 15706 25452 16118
rect 25412 15700 25464 15706
rect 25412 15642 25464 15648
rect 25228 15428 25280 15434
rect 25228 15370 25280 15376
rect 25412 15428 25464 15434
rect 25516 15416 25544 17070
rect 25464 15388 25544 15416
rect 25412 15370 25464 15376
rect 25044 14952 25096 14958
rect 25044 14894 25096 14900
rect 24860 13728 24912 13734
rect 24860 13670 24912 13676
rect 24768 13184 24820 13190
rect 24768 13126 24820 13132
rect 24780 12782 24808 13126
rect 24768 12776 24820 12782
rect 24768 12718 24820 12724
rect 24872 12434 24900 13670
rect 24688 12406 24808 12434
rect 24872 12406 24992 12434
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 24584 12164 24636 12170
rect 24584 12106 24636 12112
rect 24492 11892 24544 11898
rect 24492 11834 24544 11840
rect 24596 11286 24624 12106
rect 24584 11280 24636 11286
rect 24584 11222 24636 11228
rect 24584 11076 24636 11082
rect 24584 11018 24636 11024
rect 24596 10985 24624 11018
rect 24582 10976 24638 10985
rect 24582 10911 24638 10920
rect 24676 9920 24728 9926
rect 24676 9862 24728 9868
rect 24490 9752 24546 9761
rect 24490 9687 24546 9696
rect 24306 8871 24362 8880
rect 24400 8900 24452 8906
rect 24320 7750 24348 8871
rect 24400 8842 24452 8848
rect 24308 7744 24360 7750
rect 24308 7686 24360 7692
rect 24412 6866 24440 8842
rect 24400 6860 24452 6866
rect 24400 6802 24452 6808
rect 24504 6746 24532 9687
rect 24688 9178 24716 9862
rect 24780 9178 24808 12406
rect 24860 11824 24912 11830
rect 24860 11766 24912 11772
rect 24872 10266 24900 11766
rect 24964 11218 24992 12406
rect 24952 11212 25004 11218
rect 24952 11154 25004 11160
rect 25056 10742 25084 14894
rect 25134 14376 25190 14385
rect 25134 14311 25190 14320
rect 25148 13954 25176 14311
rect 25240 14074 25268 15370
rect 25608 15094 25636 17546
rect 25792 17542 25820 19246
rect 26056 18896 26108 18902
rect 26056 18838 26108 18844
rect 25964 18080 26016 18086
rect 25964 18022 26016 18028
rect 25780 17536 25832 17542
rect 25780 17478 25832 17484
rect 25976 17338 26004 18022
rect 26068 17678 26096 18838
rect 26056 17672 26108 17678
rect 26054 17640 26056 17649
rect 26108 17640 26110 17649
rect 26054 17575 26110 17584
rect 25964 17332 26016 17338
rect 25964 17274 26016 17280
rect 25976 16658 26004 17274
rect 25964 16652 26016 16658
rect 25964 16594 26016 16600
rect 25778 16552 25834 16561
rect 25778 16487 25780 16496
rect 25832 16487 25834 16496
rect 25780 16458 25832 16464
rect 25688 15972 25740 15978
rect 25688 15914 25740 15920
rect 25596 15088 25648 15094
rect 25596 15030 25648 15036
rect 25412 14476 25464 14482
rect 25412 14418 25464 14424
rect 25228 14068 25280 14074
rect 25228 14010 25280 14016
rect 25148 13926 25268 13954
rect 25136 13864 25188 13870
rect 25136 13806 25188 13812
rect 25148 12306 25176 13806
rect 25240 12434 25268 13926
rect 25320 13932 25372 13938
rect 25320 13874 25372 13880
rect 25332 12918 25360 13874
rect 25424 13870 25452 14418
rect 25504 14408 25556 14414
rect 25502 14376 25504 14385
rect 25556 14376 25558 14385
rect 25502 14311 25558 14320
rect 25608 14278 25636 15030
rect 25700 15026 25728 15914
rect 25964 15904 26016 15910
rect 25964 15846 26016 15852
rect 25872 15428 25924 15434
rect 25872 15370 25924 15376
rect 25688 15020 25740 15026
rect 25688 14962 25740 14968
rect 25688 14612 25740 14618
rect 25688 14554 25740 14560
rect 25596 14272 25648 14278
rect 25596 14214 25648 14220
rect 25700 13870 25728 14554
rect 25412 13864 25464 13870
rect 25412 13806 25464 13812
rect 25688 13864 25740 13870
rect 25688 13806 25740 13812
rect 25412 13456 25464 13462
rect 25412 13398 25464 13404
rect 25320 12912 25372 12918
rect 25320 12854 25372 12860
rect 25240 12406 25360 12434
rect 25136 12300 25188 12306
rect 25136 12242 25188 12248
rect 25134 12064 25190 12073
rect 25134 11999 25190 12008
rect 25148 11830 25176 11999
rect 25136 11824 25188 11830
rect 25188 11784 25268 11812
rect 25136 11766 25188 11772
rect 25134 11384 25190 11393
rect 25134 11319 25190 11328
rect 25148 11082 25176 11319
rect 25240 11218 25268 11784
rect 25228 11212 25280 11218
rect 25228 11154 25280 11160
rect 25136 11076 25188 11082
rect 25136 11018 25188 11024
rect 25228 11076 25280 11082
rect 25228 11018 25280 11024
rect 25044 10736 25096 10742
rect 25044 10678 25096 10684
rect 24860 10260 24912 10266
rect 24860 10202 24912 10208
rect 25240 10130 25268 11018
rect 25228 10124 25280 10130
rect 25228 10066 25280 10072
rect 25044 10056 25096 10062
rect 25044 9998 25096 10004
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 24676 9172 24728 9178
rect 24676 9114 24728 9120
rect 24768 9172 24820 9178
rect 24768 9114 24820 9120
rect 24768 8968 24820 8974
rect 24964 8956 24992 9658
rect 25056 9654 25084 9998
rect 25044 9648 25096 9654
rect 25332 9602 25360 12406
rect 25424 11257 25452 13398
rect 25780 13388 25832 13394
rect 25780 13330 25832 13336
rect 25686 13288 25742 13297
rect 25686 13223 25688 13232
rect 25740 13223 25742 13232
rect 25688 13194 25740 13200
rect 25792 12918 25820 13330
rect 25884 13190 25912 15370
rect 25976 14482 26004 15846
rect 26056 14952 26108 14958
rect 26056 14894 26108 14900
rect 25964 14476 26016 14482
rect 25964 14418 26016 14424
rect 26068 13870 26096 14894
rect 26056 13864 26108 13870
rect 26056 13806 26108 13812
rect 25964 13252 26016 13258
rect 25964 13194 26016 13200
rect 25872 13184 25924 13190
rect 25872 13126 25924 13132
rect 25780 12912 25832 12918
rect 25780 12854 25832 12860
rect 25872 12776 25924 12782
rect 25976 12764 26004 13194
rect 25924 12736 26004 12764
rect 26056 12776 26108 12782
rect 25872 12718 25924 12724
rect 26056 12718 26108 12724
rect 25596 12640 25648 12646
rect 25596 12582 25648 12588
rect 25608 12434 25636 12582
rect 25608 12406 25820 12434
rect 25410 11248 25466 11257
rect 25410 11183 25466 11192
rect 25424 10742 25452 11183
rect 25412 10736 25464 10742
rect 25412 10678 25464 10684
rect 25044 9590 25096 9596
rect 25056 9042 25084 9590
rect 25148 9574 25360 9602
rect 25044 9036 25096 9042
rect 25044 8978 25096 8984
rect 24820 8928 24992 8956
rect 24768 8910 24820 8916
rect 24584 7880 24636 7886
rect 24584 7822 24636 7828
rect 24412 6718 24532 6746
rect 24308 6656 24360 6662
rect 24308 6598 24360 6604
rect 24320 6458 24348 6598
rect 24216 6452 24268 6458
rect 24216 6394 24268 6400
rect 24308 6452 24360 6458
rect 24308 6394 24360 6400
rect 23940 6180 23992 6186
rect 23940 6122 23992 6128
rect 23848 5568 23900 5574
rect 23848 5510 23900 5516
rect 24032 5296 24084 5302
rect 24032 5238 24084 5244
rect 24044 5098 24072 5238
rect 24124 5228 24176 5234
rect 24124 5170 24176 5176
rect 24032 5092 24084 5098
rect 24032 5034 24084 5040
rect 24136 4826 24164 5170
rect 24228 4826 24256 6394
rect 24308 5568 24360 5574
rect 24308 5510 24360 5516
rect 24320 5273 24348 5510
rect 24412 5302 24440 6718
rect 24596 6254 24624 7822
rect 24780 7818 24808 8910
rect 24860 8492 24912 8498
rect 24860 8434 24912 8440
rect 24872 7857 24900 8434
rect 25148 8412 25176 9574
rect 25320 9512 25372 9518
rect 25320 9454 25372 9460
rect 25228 9376 25280 9382
rect 25228 9318 25280 9324
rect 25240 8537 25268 9318
rect 25332 8974 25360 9454
rect 25320 8968 25372 8974
rect 25320 8910 25372 8916
rect 25688 8968 25740 8974
rect 25688 8910 25740 8916
rect 25226 8528 25282 8537
rect 25226 8463 25282 8472
rect 25332 8430 25360 8910
rect 25700 8566 25728 8910
rect 25688 8560 25740 8566
rect 25688 8502 25740 8508
rect 25228 8424 25280 8430
rect 25148 8384 25228 8412
rect 24858 7848 24914 7857
rect 24768 7812 24820 7818
rect 24858 7783 24914 7792
rect 24768 7754 24820 7760
rect 24780 7721 24808 7754
rect 24766 7712 24822 7721
rect 24766 7647 24822 7656
rect 24952 7472 25004 7478
rect 24952 7414 25004 7420
rect 24860 6656 24912 6662
rect 24688 6616 24860 6644
rect 24584 6248 24636 6254
rect 24584 6190 24636 6196
rect 24596 6118 24624 6190
rect 24584 6112 24636 6118
rect 24584 6054 24636 6060
rect 24584 5568 24636 5574
rect 24582 5536 24584 5545
rect 24636 5536 24638 5545
rect 24582 5471 24638 5480
rect 24400 5296 24452 5302
rect 24306 5264 24362 5273
rect 24400 5238 24452 5244
rect 24306 5199 24362 5208
rect 24124 4820 24176 4826
rect 24124 4762 24176 4768
rect 24216 4820 24268 4826
rect 24216 4762 24268 4768
rect 23756 4684 23808 4690
rect 23756 4626 23808 4632
rect 23768 4486 23796 4626
rect 23756 4480 23808 4486
rect 23756 4422 23808 4428
rect 24136 4128 24164 4762
rect 24688 4758 24716 6616
rect 24860 6598 24912 6604
rect 24768 5840 24820 5846
rect 24768 5782 24820 5788
rect 24780 5137 24808 5782
rect 24964 5166 24992 7414
rect 25148 6934 25176 8384
rect 25228 8366 25280 8372
rect 25320 8424 25372 8430
rect 25320 8366 25372 8372
rect 25228 7200 25280 7206
rect 25228 7142 25280 7148
rect 25136 6928 25188 6934
rect 25136 6870 25188 6876
rect 25240 6390 25268 7142
rect 25792 6769 25820 12406
rect 25884 12306 25912 12718
rect 26068 12646 26096 12718
rect 26056 12640 26108 12646
rect 26056 12582 26108 12588
rect 26160 12434 26188 19790
rect 26332 19712 26384 19718
rect 26332 19654 26384 19660
rect 26240 19372 26292 19378
rect 26240 19314 26292 19320
rect 26252 17202 26280 19314
rect 26344 19310 26372 19654
rect 26332 19304 26384 19310
rect 26332 19246 26384 19252
rect 26332 17536 26384 17542
rect 26332 17478 26384 17484
rect 26240 17196 26292 17202
rect 26240 17138 26292 17144
rect 26240 16244 26292 16250
rect 26240 16186 26292 16192
rect 26252 14482 26280 16186
rect 26344 14804 26372 17478
rect 26436 17202 26464 27270
rect 26608 19780 26660 19786
rect 26608 19722 26660 19728
rect 26516 18624 26568 18630
rect 26516 18566 26568 18572
rect 26528 17377 26556 18566
rect 26514 17368 26570 17377
rect 26514 17303 26570 17312
rect 26424 17196 26476 17202
rect 26424 17138 26476 17144
rect 26516 17196 26568 17202
rect 26516 17138 26568 17144
rect 26436 15570 26464 17138
rect 26424 15564 26476 15570
rect 26424 15506 26476 15512
rect 26424 14816 26476 14822
rect 26344 14776 26424 14804
rect 26424 14758 26476 14764
rect 26240 14476 26292 14482
rect 26240 14418 26292 14424
rect 26332 12640 26384 12646
rect 26332 12582 26384 12588
rect 26344 12442 26372 12582
rect 26068 12406 26188 12434
rect 26332 12436 26384 12442
rect 25872 12300 25924 12306
rect 25872 12242 25924 12248
rect 25964 7472 26016 7478
rect 26068 7460 26096 12406
rect 26332 12378 26384 12384
rect 26424 12436 26476 12442
rect 26424 12378 26476 12384
rect 26148 12300 26200 12306
rect 26148 12242 26200 12248
rect 26160 11218 26188 12242
rect 26436 12170 26464 12378
rect 26424 12164 26476 12170
rect 26424 12106 26476 12112
rect 26240 11824 26292 11830
rect 26240 11766 26292 11772
rect 26252 11218 26280 11766
rect 26528 11336 26556 17138
rect 26620 13954 26648 19722
rect 26700 19712 26752 19718
rect 26700 19654 26752 19660
rect 26712 19378 26740 19654
rect 26700 19372 26752 19378
rect 26700 19314 26752 19320
rect 26988 18970 27016 30670
rect 27172 26234 27200 37198
rect 27356 32570 27384 37198
rect 28368 37126 28396 39200
rect 30300 37126 30328 39200
rect 30380 37256 30432 37262
rect 30380 37198 30432 37204
rect 30656 37256 30708 37262
rect 30656 37198 30708 37204
rect 28356 37120 28408 37126
rect 28356 37062 28408 37068
rect 30288 37120 30340 37126
rect 30288 37062 30340 37068
rect 30392 35834 30420 37198
rect 30380 35828 30432 35834
rect 30380 35770 30432 35776
rect 28540 35692 28592 35698
rect 28540 35634 28592 35640
rect 27344 32564 27396 32570
rect 27344 32506 27396 32512
rect 28552 32366 28580 35634
rect 28540 32360 28592 32366
rect 28540 32302 28592 32308
rect 28552 28082 28580 32302
rect 28632 32224 28684 32230
rect 28632 32166 28684 32172
rect 28540 28076 28592 28082
rect 28540 28018 28592 28024
rect 27080 26206 27200 26234
rect 26976 18964 27028 18970
rect 26976 18906 27028 18912
rect 26700 18624 26752 18630
rect 26700 18566 26752 18572
rect 26712 18290 26740 18566
rect 26700 18284 26752 18290
rect 26700 18226 26752 18232
rect 26792 17740 26844 17746
rect 26792 17682 26844 17688
rect 26804 16998 26832 17682
rect 26884 17672 26936 17678
rect 26884 17614 26936 17620
rect 26896 17202 26924 17614
rect 26884 17196 26936 17202
rect 26884 17138 26936 17144
rect 26792 16992 26844 16998
rect 26792 16934 26844 16940
rect 26700 16516 26752 16522
rect 26700 16458 26752 16464
rect 26712 16250 26740 16458
rect 26700 16244 26752 16250
rect 26700 16186 26752 16192
rect 26792 16040 26844 16046
rect 26792 15982 26844 15988
rect 26698 15056 26754 15065
rect 26698 14991 26700 15000
rect 26752 14991 26754 15000
rect 26700 14962 26752 14968
rect 26804 14550 26832 15982
rect 26976 15360 27028 15366
rect 26976 15302 27028 15308
rect 26884 14884 26936 14890
rect 26884 14826 26936 14832
rect 26792 14544 26844 14550
rect 26792 14486 26844 14492
rect 26896 14074 26924 14826
rect 26988 14550 27016 15302
rect 26976 14544 27028 14550
rect 26976 14486 27028 14492
rect 26988 14074 27016 14486
rect 26884 14068 26936 14074
rect 26884 14010 26936 14016
rect 26976 14068 27028 14074
rect 26976 14010 27028 14016
rect 26620 13926 26924 13954
rect 26608 13864 26660 13870
rect 26608 13806 26660 13812
rect 26620 11540 26648 13806
rect 26620 11512 26740 11540
rect 26528 11308 26648 11336
rect 26514 11248 26570 11257
rect 26148 11212 26200 11218
rect 26148 11154 26200 11160
rect 26240 11212 26292 11218
rect 26514 11183 26570 11192
rect 26240 11154 26292 11160
rect 26424 10532 26476 10538
rect 26424 10474 26476 10480
rect 26436 10441 26464 10474
rect 26422 10432 26478 10441
rect 26422 10367 26478 10376
rect 26146 10296 26202 10305
rect 26146 10231 26148 10240
rect 26200 10231 26202 10240
rect 26148 10202 26200 10208
rect 26160 9178 26188 10202
rect 26528 9518 26556 11183
rect 26516 9512 26568 9518
rect 26516 9454 26568 9460
rect 26148 9172 26200 9178
rect 26148 9114 26200 9120
rect 26240 9036 26292 9042
rect 26240 8978 26292 8984
rect 26252 8430 26280 8978
rect 26424 8900 26476 8906
rect 26424 8842 26476 8848
rect 26240 8424 26292 8430
rect 26240 8366 26292 8372
rect 26016 7432 26096 7460
rect 25964 7414 26016 7420
rect 25872 7336 25924 7342
rect 25872 7278 25924 7284
rect 25778 6760 25834 6769
rect 25778 6695 25834 6704
rect 25228 6384 25280 6390
rect 25228 6326 25280 6332
rect 25792 5302 25820 6695
rect 25884 5658 25912 7278
rect 26068 7002 26096 7432
rect 26252 7410 26280 8366
rect 26436 8362 26464 8842
rect 26528 8838 26556 9454
rect 26516 8832 26568 8838
rect 26516 8774 26568 8780
rect 26424 8356 26476 8362
rect 26424 8298 26476 8304
rect 26240 7404 26292 7410
rect 26240 7346 26292 7352
rect 26332 7336 26384 7342
rect 26332 7278 26384 7284
rect 26056 6996 26108 7002
rect 26056 6938 26108 6944
rect 26148 6860 26200 6866
rect 26148 6802 26200 6808
rect 26056 6316 26108 6322
rect 26056 6258 26108 6264
rect 26068 5914 26096 6258
rect 26160 5930 26188 6802
rect 26344 6746 26372 7278
rect 26252 6730 26464 6746
rect 26240 6724 26464 6730
rect 26292 6718 26464 6724
rect 26240 6666 26292 6672
rect 26436 6662 26464 6718
rect 26424 6656 26476 6662
rect 26424 6598 26476 6604
rect 26620 6458 26648 11308
rect 26712 7342 26740 11512
rect 26790 11112 26846 11121
rect 26790 11047 26846 11056
rect 26804 11014 26832 11047
rect 26792 11008 26844 11014
rect 26792 10950 26844 10956
rect 26896 10198 26924 13926
rect 26988 12918 27016 14010
rect 26976 12912 27028 12918
rect 26976 12854 27028 12860
rect 27080 11354 27108 26206
rect 27804 24200 27856 24206
rect 27804 24142 27856 24148
rect 27816 22094 27844 24142
rect 27724 22066 27844 22094
rect 27528 20800 27580 20806
rect 27528 20742 27580 20748
rect 27160 19372 27212 19378
rect 27160 19314 27212 19320
rect 27172 18193 27200 19314
rect 27344 19168 27396 19174
rect 27344 19110 27396 19116
rect 27252 18760 27304 18766
rect 27252 18702 27304 18708
rect 27158 18184 27214 18193
rect 27158 18119 27214 18128
rect 27172 13870 27200 18119
rect 27264 17921 27292 18702
rect 27250 17912 27306 17921
rect 27250 17847 27306 17856
rect 27356 17762 27384 19110
rect 27540 17882 27568 20742
rect 27620 19168 27672 19174
rect 27620 19110 27672 19116
rect 27632 18698 27660 19110
rect 27620 18692 27672 18698
rect 27620 18634 27672 18640
rect 27528 17876 27580 17882
rect 27528 17818 27580 17824
rect 27264 17734 27384 17762
rect 27264 16454 27292 17734
rect 27540 17678 27568 17818
rect 27528 17672 27580 17678
rect 27528 17614 27580 17620
rect 27436 17536 27488 17542
rect 27436 17478 27488 17484
rect 27528 17536 27580 17542
rect 27528 17478 27580 17484
rect 27344 16992 27396 16998
rect 27344 16934 27396 16940
rect 27252 16448 27304 16454
rect 27252 16390 27304 16396
rect 27264 15994 27292 16390
rect 27356 16182 27384 16934
rect 27344 16176 27396 16182
rect 27344 16118 27396 16124
rect 27448 16046 27476 17478
rect 27540 17134 27568 17478
rect 27528 17128 27580 17134
rect 27528 17070 27580 17076
rect 27436 16040 27488 16046
rect 27264 15966 27384 15994
rect 27528 16040 27580 16046
rect 27436 15982 27488 15988
rect 27526 16008 27528 16017
rect 27580 16008 27582 16017
rect 27252 15360 27304 15366
rect 27252 15302 27304 15308
rect 27264 14958 27292 15302
rect 27252 14952 27304 14958
rect 27252 14894 27304 14900
rect 27250 14512 27306 14521
rect 27250 14447 27306 14456
rect 27264 14346 27292 14447
rect 27252 14340 27304 14346
rect 27252 14282 27304 14288
rect 27160 13864 27212 13870
rect 27160 13806 27212 13812
rect 27252 13728 27304 13734
rect 27252 13670 27304 13676
rect 27160 13524 27212 13530
rect 27160 13466 27212 13472
rect 27068 11348 27120 11354
rect 27068 11290 27120 11296
rect 27172 10690 27200 13466
rect 27264 13394 27292 13670
rect 27252 13388 27304 13394
rect 27252 13330 27304 13336
rect 27250 11520 27306 11529
rect 27250 11455 27306 11464
rect 27264 11354 27292 11455
rect 27252 11348 27304 11354
rect 27252 11290 27304 11296
rect 26988 10662 27200 10690
rect 26884 10192 26936 10198
rect 26884 10134 26936 10140
rect 26792 9172 26844 9178
rect 26792 9114 26844 9120
rect 26700 7336 26752 7342
rect 26700 7278 26752 7284
rect 26608 6452 26660 6458
rect 26608 6394 26660 6400
rect 26424 6384 26476 6390
rect 26424 6326 26476 6332
rect 26436 6118 26464 6326
rect 26608 6316 26660 6322
rect 26608 6258 26660 6264
rect 26514 6216 26570 6225
rect 26514 6151 26570 6160
rect 26528 6118 26556 6151
rect 26424 6112 26476 6118
rect 26424 6054 26476 6060
rect 26516 6112 26568 6118
rect 26516 6054 26568 6060
rect 25964 5908 26016 5914
rect 25964 5850 26016 5856
rect 26056 5908 26108 5914
rect 26160 5902 26464 5930
rect 26056 5850 26108 5856
rect 25976 5794 26004 5850
rect 25976 5766 26280 5794
rect 26436 5778 26464 5902
rect 25884 5642 26096 5658
rect 25884 5636 26108 5642
rect 25884 5630 26056 5636
rect 26056 5578 26108 5584
rect 25780 5296 25832 5302
rect 25134 5264 25190 5273
rect 25780 5238 25832 5244
rect 25134 5199 25190 5208
rect 25148 5166 25176 5199
rect 24952 5160 25004 5166
rect 24766 5128 24822 5137
rect 24952 5102 25004 5108
rect 25136 5160 25188 5166
rect 25136 5102 25188 5108
rect 24766 5063 24822 5072
rect 24860 4820 24912 4826
rect 24860 4762 24912 4768
rect 24676 4752 24728 4758
rect 24676 4694 24728 4700
rect 24872 4690 24900 4762
rect 24492 4684 24544 4690
rect 24492 4626 24544 4632
rect 24860 4684 24912 4690
rect 24860 4626 24912 4632
rect 24216 4140 24268 4146
rect 24136 4100 24216 4128
rect 24268 4100 24348 4128
rect 24216 4082 24268 4088
rect 23664 4004 23716 4010
rect 23664 3946 23716 3952
rect 24216 4004 24268 4010
rect 24216 3946 24268 3952
rect 24032 3936 24084 3942
rect 24032 3878 24084 3884
rect 23940 3528 23992 3534
rect 23940 3470 23992 3476
rect 23952 3398 23980 3470
rect 23848 3392 23900 3398
rect 23848 3334 23900 3340
rect 23940 3392 23992 3398
rect 23940 3334 23992 3340
rect 23664 2984 23716 2990
rect 23664 2926 23716 2932
rect 23572 2916 23624 2922
rect 23572 2858 23624 2864
rect 23308 2746 23428 2774
rect 22008 2508 22060 2514
rect 22008 2450 22060 2456
rect 23400 2378 23428 2746
rect 23676 2650 23704 2926
rect 23664 2644 23716 2650
rect 23664 2586 23716 2592
rect 23388 2372 23440 2378
rect 23388 2314 23440 2320
rect 23572 2372 23624 2378
rect 23572 2314 23624 2320
rect 23584 1902 23612 2314
rect 23572 1896 23624 1902
rect 23572 1838 23624 1844
rect 23860 800 23888 3334
rect 24044 3126 24072 3878
rect 24228 3534 24256 3946
rect 24320 3602 24348 4100
rect 24504 4078 24532 4626
rect 24676 4480 24728 4486
rect 24676 4422 24728 4428
rect 24688 4282 24716 4422
rect 24676 4276 24728 4282
rect 24676 4218 24728 4224
rect 24952 4208 25004 4214
rect 24950 4176 24952 4185
rect 25004 4176 25006 4185
rect 24950 4111 25006 4120
rect 24492 4072 24544 4078
rect 24492 4014 24544 4020
rect 26068 3992 26096 5578
rect 26148 4004 26200 4010
rect 26068 3964 26148 3992
rect 26148 3946 26200 3952
rect 25964 3936 26016 3942
rect 25964 3878 26016 3884
rect 24308 3596 24360 3602
rect 24308 3538 24360 3544
rect 24584 3596 24636 3602
rect 24584 3538 24636 3544
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24032 3120 24084 3126
rect 24032 3062 24084 3068
rect 24596 3058 24624 3538
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 24596 2514 24624 2994
rect 25228 2984 25280 2990
rect 25228 2926 25280 2932
rect 25240 2774 25268 2926
rect 25148 2746 25268 2774
rect 24584 2508 24636 2514
rect 24584 2450 24636 2456
rect 25148 800 25176 2746
rect 25976 2514 26004 3878
rect 26252 3058 26280 5766
rect 26424 5772 26476 5778
rect 26424 5714 26476 5720
rect 26332 5704 26384 5710
rect 26332 5646 26384 5652
rect 26344 4622 26372 5646
rect 26516 5296 26568 5302
rect 26516 5238 26568 5244
rect 26424 4820 26476 4826
rect 26424 4762 26476 4768
rect 26332 4616 26384 4622
rect 26332 4558 26384 4564
rect 26344 4078 26372 4558
rect 26436 4146 26464 4762
rect 26528 4146 26556 5238
rect 26424 4140 26476 4146
rect 26424 4082 26476 4088
rect 26516 4140 26568 4146
rect 26516 4082 26568 4088
rect 26332 4072 26384 4078
rect 26332 4014 26384 4020
rect 26344 3602 26372 4014
rect 26424 4004 26476 4010
rect 26424 3946 26476 3952
rect 26436 3670 26464 3946
rect 26620 3913 26648 6258
rect 26698 4856 26754 4865
rect 26698 4791 26700 4800
rect 26752 4791 26754 4800
rect 26700 4762 26752 4768
rect 26804 4729 26832 9114
rect 26988 6882 27016 10662
rect 27160 10600 27212 10606
rect 27160 10542 27212 10548
rect 27172 8838 27200 10542
rect 27252 9920 27304 9926
rect 27252 9862 27304 9868
rect 27264 9761 27292 9862
rect 27250 9752 27306 9761
rect 27250 9687 27306 9696
rect 27252 9104 27304 9110
rect 27252 9046 27304 9052
rect 27160 8832 27212 8838
rect 27160 8774 27212 8780
rect 27172 8430 27200 8774
rect 27160 8424 27212 8430
rect 27160 8366 27212 8372
rect 27068 8356 27120 8362
rect 27068 8298 27120 8304
rect 27080 7546 27108 8298
rect 27172 7886 27200 8366
rect 27160 7880 27212 7886
rect 27160 7822 27212 7828
rect 27068 7540 27120 7546
rect 27068 7482 27120 7488
rect 27172 7342 27200 7822
rect 27264 7750 27292 9046
rect 27252 7744 27304 7750
rect 27252 7686 27304 7692
rect 27356 7478 27384 15966
rect 27526 15943 27582 15952
rect 27540 15434 27568 15943
rect 27528 15428 27580 15434
rect 27528 15370 27580 15376
rect 27436 14340 27488 14346
rect 27436 14282 27488 14288
rect 27448 13682 27476 14282
rect 27620 14272 27672 14278
rect 27620 14214 27672 14220
rect 27632 13870 27660 14214
rect 27620 13864 27672 13870
rect 27620 13806 27672 13812
rect 27526 13696 27582 13705
rect 27448 13654 27526 13682
rect 27526 13631 27582 13640
rect 27540 13258 27568 13631
rect 27620 13388 27672 13394
rect 27620 13330 27672 13336
rect 27632 13297 27660 13330
rect 27618 13288 27674 13297
rect 27528 13252 27580 13258
rect 27618 13223 27674 13232
rect 27528 13194 27580 13200
rect 27436 12368 27488 12374
rect 27436 12310 27488 12316
rect 27448 11694 27476 12310
rect 27528 12164 27580 12170
rect 27528 12106 27580 12112
rect 27540 11694 27568 12106
rect 27436 11688 27488 11694
rect 27436 11630 27488 11636
rect 27528 11688 27580 11694
rect 27528 11630 27580 11636
rect 27724 11286 27752 22066
rect 28172 17672 28224 17678
rect 28172 17614 28224 17620
rect 28080 17196 28132 17202
rect 28080 17138 28132 17144
rect 27896 16992 27948 16998
rect 27896 16934 27948 16940
rect 27988 16992 28040 16998
rect 27988 16934 28040 16940
rect 27908 15570 27936 16934
rect 28000 16590 28028 16934
rect 27988 16584 28040 16590
rect 27988 16526 28040 16532
rect 27896 15564 27948 15570
rect 27896 15506 27948 15512
rect 28000 13938 28028 16526
rect 27988 13932 28040 13938
rect 27988 13874 28040 13880
rect 27896 12708 27948 12714
rect 27896 12650 27948 12656
rect 27802 11928 27858 11937
rect 27802 11863 27858 11872
rect 27712 11280 27764 11286
rect 27712 11222 27764 11228
rect 27816 11082 27844 11863
rect 27804 11076 27856 11082
rect 27804 11018 27856 11024
rect 27804 10736 27856 10742
rect 27804 10678 27856 10684
rect 27816 10062 27844 10678
rect 27804 10056 27856 10062
rect 27804 9998 27856 10004
rect 27436 9648 27488 9654
rect 27436 9590 27488 9596
rect 27344 7472 27396 7478
rect 27344 7414 27396 7420
rect 27160 7336 27212 7342
rect 27160 7278 27212 7284
rect 27342 7304 27398 7313
rect 26896 6854 27016 6882
rect 26896 6390 26924 6854
rect 27172 6798 27200 7278
rect 27342 7239 27398 7248
rect 27356 6866 27384 7239
rect 27344 6860 27396 6866
rect 27344 6802 27396 6808
rect 27160 6792 27212 6798
rect 27160 6734 27212 6740
rect 26884 6384 26936 6390
rect 26884 6326 26936 6332
rect 27068 6384 27120 6390
rect 27068 6326 27120 6332
rect 26896 5234 26924 6326
rect 26884 5228 26936 5234
rect 26884 5170 26936 5176
rect 26790 4720 26846 4729
rect 26790 4655 26846 4664
rect 26700 3936 26752 3942
rect 26606 3904 26662 3913
rect 26700 3878 26752 3884
rect 26606 3839 26662 3848
rect 26424 3664 26476 3670
rect 26424 3606 26476 3612
rect 26332 3596 26384 3602
rect 26332 3538 26384 3544
rect 26516 3596 26568 3602
rect 26516 3538 26568 3544
rect 26528 3233 26556 3538
rect 26712 3398 26740 3878
rect 27080 3466 27108 6326
rect 27172 6186 27200 6734
rect 27448 6497 27476 9590
rect 27528 8900 27580 8906
rect 27528 8842 27580 8848
rect 27540 8809 27568 8842
rect 27526 8800 27582 8809
rect 27526 8735 27582 8744
rect 27528 8560 27580 8566
rect 27528 8502 27580 8508
rect 27540 8430 27568 8502
rect 27528 8424 27580 8430
rect 27528 8366 27580 8372
rect 27526 8120 27582 8129
rect 27526 8055 27582 8064
rect 27434 6488 27490 6497
rect 27434 6423 27490 6432
rect 27160 6180 27212 6186
rect 27160 6122 27212 6128
rect 27172 5710 27200 6122
rect 27540 5778 27568 8055
rect 27620 7744 27672 7750
rect 27618 7712 27620 7721
rect 27672 7712 27674 7721
rect 27618 7647 27674 7656
rect 27528 5772 27580 5778
rect 27528 5714 27580 5720
rect 27160 5704 27212 5710
rect 27160 5646 27212 5652
rect 27436 4072 27488 4078
rect 27436 4014 27488 4020
rect 27068 3460 27120 3466
rect 27068 3402 27120 3408
rect 27252 3460 27304 3466
rect 27252 3402 27304 3408
rect 26700 3392 26752 3398
rect 26700 3334 26752 3340
rect 26514 3224 26570 3233
rect 26514 3159 26570 3168
rect 27264 3058 27292 3402
rect 26240 3052 26292 3058
rect 26240 2994 26292 3000
rect 27252 3052 27304 3058
rect 27252 2994 27304 3000
rect 26792 2984 26844 2990
rect 26790 2952 26792 2961
rect 26844 2952 26846 2961
rect 26790 2887 26846 2896
rect 25964 2508 26016 2514
rect 25964 2450 26016 2456
rect 27448 2446 27476 4014
rect 27908 3670 27936 12650
rect 27986 12472 28042 12481
rect 27986 12407 28042 12416
rect 28000 11121 28028 12407
rect 27986 11112 28042 11121
rect 27986 11047 28042 11056
rect 28000 8974 28028 11047
rect 27988 8968 28040 8974
rect 27988 8910 28040 8916
rect 27988 6656 28040 6662
rect 27988 6598 28040 6604
rect 28000 5166 28028 6598
rect 27988 5160 28040 5166
rect 27988 5102 28040 5108
rect 27896 3664 27948 3670
rect 27896 3606 27948 3612
rect 27802 3496 27858 3505
rect 28092 3482 28120 17138
rect 28184 17066 28212 17614
rect 28644 17202 28672 32166
rect 30668 30938 30696 37198
rect 32232 37126 32260 39200
rect 33520 37126 33548 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 33600 37256 33652 37262
rect 33600 37198 33652 37204
rect 34796 37256 34848 37262
rect 34796 37198 34848 37204
rect 32220 37120 32272 37126
rect 32220 37062 32272 37068
rect 33508 37120 33560 37126
rect 33508 37062 33560 37068
rect 33612 36922 33640 37198
rect 34808 37126 34836 37198
rect 35452 37126 35480 39200
rect 36818 38856 36874 38865
rect 36818 38791 36874 38800
rect 36832 37466 36860 38791
rect 36820 37460 36872 37466
rect 36820 37402 36872 37408
rect 36452 37188 36504 37194
rect 36452 37130 36504 37136
rect 34796 37120 34848 37126
rect 34796 37062 34848 37068
rect 35440 37120 35492 37126
rect 35440 37062 35492 37068
rect 36268 37120 36320 37126
rect 36268 37062 36320 37068
rect 33600 36916 33652 36922
rect 33600 36858 33652 36864
rect 30656 30932 30708 30938
rect 30656 30874 30708 30880
rect 30196 30252 30248 30258
rect 30196 30194 30248 30200
rect 30012 21548 30064 21554
rect 30012 21490 30064 21496
rect 30024 20806 30052 21490
rect 30012 20800 30064 20806
rect 30012 20742 30064 20748
rect 30208 18834 30236 30194
rect 33600 19372 33652 19378
rect 33600 19314 33652 19320
rect 30196 18828 30248 18834
rect 30196 18770 30248 18776
rect 29276 18624 29328 18630
rect 29276 18566 29328 18572
rect 29000 18080 29052 18086
rect 29000 18022 29052 18028
rect 28724 17604 28776 17610
rect 28724 17546 28776 17552
rect 28632 17196 28684 17202
rect 28632 17138 28684 17144
rect 28736 17134 28764 17546
rect 29012 17270 29040 18022
rect 29000 17264 29052 17270
rect 29000 17206 29052 17212
rect 28908 17196 28960 17202
rect 28908 17138 28960 17144
rect 28724 17128 28776 17134
rect 28724 17070 28776 17076
rect 28172 17060 28224 17066
rect 28172 17002 28224 17008
rect 28736 16538 28764 17070
rect 28920 16726 28948 17138
rect 28908 16720 28960 16726
rect 28908 16662 28960 16668
rect 28644 16510 28764 16538
rect 28448 16244 28500 16250
rect 28448 16186 28500 16192
rect 28172 15904 28224 15910
rect 28172 15846 28224 15852
rect 28184 15162 28212 15846
rect 28264 15496 28316 15502
rect 28264 15438 28316 15444
rect 28276 15337 28304 15438
rect 28262 15328 28318 15337
rect 28262 15263 28318 15272
rect 28172 15156 28224 15162
rect 28172 15098 28224 15104
rect 28276 15026 28304 15263
rect 28264 15020 28316 15026
rect 28264 14962 28316 14968
rect 28356 15020 28408 15026
rect 28356 14962 28408 14968
rect 28368 14822 28396 14962
rect 28356 14816 28408 14822
rect 28356 14758 28408 14764
rect 28460 14657 28488 16186
rect 28540 15632 28592 15638
rect 28540 15574 28592 15580
rect 28552 15434 28580 15574
rect 28540 15428 28592 15434
rect 28540 15370 28592 15376
rect 28538 15192 28594 15201
rect 28538 15127 28594 15136
rect 28446 14648 28502 14657
rect 28446 14583 28502 14592
rect 28448 14408 28500 14414
rect 28552 14396 28580 15127
rect 28644 14929 28672 16510
rect 29184 16448 29236 16454
rect 29184 16390 29236 16396
rect 29196 16114 29224 16390
rect 29184 16108 29236 16114
rect 29184 16050 29236 16056
rect 28724 15972 28776 15978
rect 28724 15914 28776 15920
rect 28736 15026 28764 15914
rect 28816 15904 28868 15910
rect 28816 15846 28868 15852
rect 28828 15706 28856 15846
rect 28816 15700 28868 15706
rect 28816 15642 28868 15648
rect 29092 15564 29144 15570
rect 29092 15506 29144 15512
rect 28814 15328 28870 15337
rect 28814 15263 28870 15272
rect 28998 15328 29054 15337
rect 28998 15263 29054 15272
rect 28828 15026 28856 15263
rect 28906 15192 28962 15201
rect 28906 15127 28962 15136
rect 28724 15020 28776 15026
rect 28724 14962 28776 14968
rect 28816 15020 28868 15026
rect 28920 15008 28948 15127
rect 29012 15008 29040 15263
rect 28920 14980 29040 15008
rect 28816 14962 28868 14968
rect 29104 14940 29132 15506
rect 29182 15464 29238 15473
rect 29182 15399 29238 15408
rect 28630 14920 28686 14929
rect 29012 14912 29132 14940
rect 28630 14855 28686 14864
rect 28816 14884 28868 14890
rect 28500 14368 28580 14396
rect 28448 14350 28500 14356
rect 28262 14104 28318 14113
rect 28262 14039 28264 14048
rect 28316 14039 28318 14048
rect 28264 14010 28316 14016
rect 28172 14000 28224 14006
rect 28540 14000 28592 14006
rect 28224 13948 28540 13954
rect 28172 13942 28592 13948
rect 28184 13926 28580 13942
rect 28172 13796 28224 13802
rect 28172 13738 28224 13744
rect 28184 13462 28212 13738
rect 28172 13456 28224 13462
rect 28172 13398 28224 13404
rect 28448 12708 28500 12714
rect 28448 12650 28500 12656
rect 28460 12442 28488 12650
rect 28448 12436 28500 12442
rect 28448 12378 28500 12384
rect 28540 12436 28592 12442
rect 28540 12378 28592 12384
rect 28356 12164 28408 12170
rect 28356 12106 28408 12112
rect 28448 12164 28500 12170
rect 28448 12106 28500 12112
rect 28264 11756 28316 11762
rect 28264 11698 28316 11704
rect 28170 11656 28226 11665
rect 28170 11591 28172 11600
rect 28224 11591 28226 11600
rect 28172 11562 28224 11568
rect 28172 10804 28224 10810
rect 28276 10792 28304 11698
rect 28368 11218 28396 12106
rect 28460 11608 28488 12106
rect 28552 12073 28580 12378
rect 28538 12064 28594 12073
rect 28538 11999 28594 12008
rect 28540 11620 28592 11626
rect 28460 11580 28540 11608
rect 28356 11212 28408 11218
rect 28356 11154 28408 11160
rect 28460 10985 28488 11580
rect 28540 11562 28592 11568
rect 28446 10976 28502 10985
rect 28446 10911 28502 10920
rect 28224 10764 28304 10792
rect 28172 10746 28224 10752
rect 28184 9674 28212 10746
rect 28184 9646 28304 9674
rect 28276 4690 28304 9646
rect 28644 8022 28672 14855
rect 28868 14844 28948 14872
rect 28816 14826 28868 14832
rect 28920 14770 28948 14844
rect 28828 14742 28948 14770
rect 28828 14618 28856 14742
rect 28906 14648 28962 14657
rect 28816 14612 28868 14618
rect 28906 14583 28908 14592
rect 28816 14554 28868 14560
rect 28960 14583 28962 14592
rect 28908 14554 28960 14560
rect 28906 14512 28962 14521
rect 28906 14447 28908 14456
rect 28960 14447 28962 14456
rect 28908 14418 28960 14424
rect 29012 14278 29040 14912
rect 29196 14657 29224 15399
rect 29182 14648 29238 14657
rect 29182 14583 29238 14592
rect 29196 14414 29224 14583
rect 29184 14408 29236 14414
rect 29184 14350 29236 14356
rect 29000 14272 29052 14278
rect 29000 14214 29052 14220
rect 28724 14000 28776 14006
rect 28724 13942 28776 13948
rect 28736 11898 28764 13942
rect 29184 13864 29236 13870
rect 28998 13832 29054 13841
rect 28908 13796 28960 13802
rect 28998 13767 29000 13776
rect 28908 13738 28960 13744
rect 29052 13767 29054 13776
rect 29182 13832 29184 13841
rect 29236 13832 29238 13841
rect 29182 13767 29238 13776
rect 29000 13738 29052 13744
rect 28920 13530 28948 13738
rect 29182 13696 29238 13705
rect 29182 13631 29238 13640
rect 28908 13524 28960 13530
rect 28908 13466 28960 13472
rect 28920 12850 28948 13466
rect 29000 13388 29052 13394
rect 29000 13330 29052 13336
rect 29012 13025 29040 13330
rect 29196 13258 29224 13631
rect 29184 13252 29236 13258
rect 29184 13194 29236 13200
rect 28998 13016 29054 13025
rect 28998 12951 29054 12960
rect 28998 12880 29054 12889
rect 28908 12844 28960 12850
rect 28998 12815 29000 12824
rect 28908 12786 28960 12792
rect 29052 12815 29054 12824
rect 29000 12786 29052 12792
rect 29184 12776 29236 12782
rect 29184 12718 29236 12724
rect 28998 12336 29054 12345
rect 28998 12271 29000 12280
rect 29052 12271 29054 12280
rect 29000 12242 29052 12248
rect 29000 12164 29052 12170
rect 29000 12106 29052 12112
rect 28724 11892 28776 11898
rect 28724 11834 28776 11840
rect 29012 11529 29040 12106
rect 29092 12096 29144 12102
rect 29090 12064 29092 12073
rect 29144 12064 29146 12073
rect 29090 11999 29146 12008
rect 29090 11792 29146 11801
rect 29090 11727 29092 11736
rect 29144 11727 29146 11736
rect 29092 11698 29144 11704
rect 29092 11552 29144 11558
rect 28998 11520 29054 11529
rect 29092 11494 29144 11500
rect 28998 11455 29054 11464
rect 29104 11354 29132 11494
rect 29196 11393 29224 12718
rect 29182 11384 29238 11393
rect 29092 11348 29144 11354
rect 29182 11319 29238 11328
rect 29092 11290 29144 11296
rect 29090 11248 29146 11257
rect 29090 11183 29146 11192
rect 29104 11150 29132 11183
rect 28724 11144 28776 11150
rect 28724 11086 28776 11092
rect 29092 11144 29144 11150
rect 29092 11086 29144 11092
rect 29184 11144 29236 11150
rect 29184 11086 29236 11092
rect 28736 9722 28764 11086
rect 29196 11014 29224 11086
rect 29184 11008 29236 11014
rect 29184 10950 29236 10956
rect 29000 10192 29052 10198
rect 29000 10134 29052 10140
rect 28908 9988 28960 9994
rect 28908 9930 28960 9936
rect 28920 9874 28948 9930
rect 29012 9874 29040 10134
rect 29092 9988 29144 9994
rect 29092 9930 29144 9936
rect 28920 9846 29040 9874
rect 28724 9716 28776 9722
rect 28724 9658 28776 9664
rect 28632 8016 28684 8022
rect 28632 7958 28684 7964
rect 28644 7274 28672 7958
rect 28632 7268 28684 7274
rect 28632 7210 28684 7216
rect 28356 6452 28408 6458
rect 28356 6394 28408 6400
rect 28368 6186 28396 6394
rect 28736 6390 28764 9658
rect 29012 8650 29040 9846
rect 29104 8838 29132 9930
rect 29092 8832 29144 8838
rect 29092 8774 29144 8780
rect 29012 8622 29224 8650
rect 29000 7744 29052 7750
rect 29000 7686 29052 7692
rect 29012 7562 29040 7686
rect 28920 7534 29040 7562
rect 28920 7274 28948 7534
rect 29000 7404 29052 7410
rect 29000 7346 29052 7352
rect 28908 7268 28960 7274
rect 28908 7210 28960 7216
rect 29012 7002 29040 7346
rect 29000 6996 29052 7002
rect 29000 6938 29052 6944
rect 29000 6792 29052 6798
rect 29000 6734 29052 6740
rect 28816 6656 28868 6662
rect 28814 6624 28816 6633
rect 28908 6656 28960 6662
rect 28868 6624 28870 6633
rect 28908 6598 28960 6604
rect 28814 6559 28870 6568
rect 28724 6384 28776 6390
rect 28724 6326 28776 6332
rect 28356 6180 28408 6186
rect 28356 6122 28408 6128
rect 28920 5778 28948 6598
rect 29012 6458 29040 6734
rect 29000 6452 29052 6458
rect 29000 6394 29052 6400
rect 28908 5772 28960 5778
rect 28908 5714 28960 5720
rect 29012 5642 29040 6394
rect 29092 6384 29144 6390
rect 29090 6352 29092 6361
rect 29144 6352 29146 6361
rect 29090 6287 29146 6296
rect 29000 5636 29052 5642
rect 29000 5578 29052 5584
rect 29012 4690 29040 5578
rect 28264 4684 28316 4690
rect 28264 4626 28316 4632
rect 29000 4684 29052 4690
rect 29000 4626 29052 4632
rect 29196 4554 29224 8622
rect 29288 8430 29316 18566
rect 29460 18080 29512 18086
rect 29460 18022 29512 18028
rect 29472 17066 29500 18022
rect 30288 17332 30340 17338
rect 30288 17274 30340 17280
rect 30012 17128 30064 17134
rect 30012 17070 30064 17076
rect 29460 17060 29512 17066
rect 29460 17002 29512 17008
rect 29368 15904 29420 15910
rect 29368 15846 29420 15852
rect 29380 14550 29408 15846
rect 29828 15496 29880 15502
rect 29828 15438 29880 15444
rect 29920 15496 29972 15502
rect 29920 15438 29972 15444
rect 29458 15328 29514 15337
rect 29458 15263 29514 15272
rect 29472 15162 29500 15263
rect 29460 15156 29512 15162
rect 29460 15098 29512 15104
rect 29552 14884 29604 14890
rect 29552 14826 29604 14832
rect 29368 14544 29420 14550
rect 29368 14486 29420 14492
rect 29460 14544 29512 14550
rect 29460 14486 29512 14492
rect 29368 14408 29420 14414
rect 29366 14376 29368 14385
rect 29420 14376 29422 14385
rect 29366 14311 29422 14320
rect 29472 14090 29500 14486
rect 29564 14278 29592 14826
rect 29644 14816 29696 14822
rect 29644 14758 29696 14764
rect 29552 14272 29604 14278
rect 29552 14214 29604 14220
rect 29380 14062 29500 14090
rect 29276 8424 29328 8430
rect 29276 8366 29328 8372
rect 29288 7206 29316 8366
rect 29276 7200 29328 7206
rect 29274 7168 29276 7177
rect 29328 7168 29330 7177
rect 29274 7103 29330 7112
rect 29274 6352 29330 6361
rect 29274 6287 29276 6296
rect 29328 6287 29330 6296
rect 29276 6258 29328 6264
rect 28908 4548 28960 4554
rect 28908 4490 28960 4496
rect 29184 4548 29236 4554
rect 29184 4490 29236 4496
rect 28816 4004 28868 4010
rect 28816 3946 28868 3952
rect 28828 3738 28856 3946
rect 28816 3732 28868 3738
rect 28816 3674 28868 3680
rect 27802 3431 27858 3440
rect 28000 3454 28120 3482
rect 27816 3126 27844 3431
rect 27804 3120 27856 3126
rect 27804 3062 27856 3068
rect 28000 3058 28028 3454
rect 28080 3392 28132 3398
rect 28080 3334 28132 3340
rect 28092 3194 28120 3334
rect 28080 3188 28132 3194
rect 28080 3130 28132 3136
rect 28920 3126 28948 4490
rect 29000 4480 29052 4486
rect 29000 4422 29052 4428
rect 29012 3942 29040 4422
rect 29380 4078 29408 14062
rect 29460 14000 29512 14006
rect 29460 13942 29512 13948
rect 29550 13968 29606 13977
rect 29472 10198 29500 13942
rect 29550 13903 29606 13912
rect 29460 10192 29512 10198
rect 29460 10134 29512 10140
rect 29460 9036 29512 9042
rect 29460 8978 29512 8984
rect 29472 5953 29500 8978
rect 29564 7546 29592 13903
rect 29656 13258 29684 14758
rect 29840 13938 29868 15438
rect 29932 13977 29960 15438
rect 30024 15065 30052 17070
rect 30010 15056 30066 15065
rect 30010 14991 30066 15000
rect 29918 13968 29974 13977
rect 29828 13932 29880 13938
rect 29918 13903 29974 13912
rect 29828 13874 29880 13880
rect 29920 13864 29972 13870
rect 29918 13832 29920 13841
rect 29972 13832 29974 13841
rect 29918 13767 29974 13776
rect 29736 13728 29788 13734
rect 29736 13670 29788 13676
rect 29748 13462 29776 13670
rect 29736 13456 29788 13462
rect 29736 13398 29788 13404
rect 29828 13456 29880 13462
rect 29828 13398 29880 13404
rect 29644 13252 29696 13258
rect 29644 13194 29696 13200
rect 29840 12918 29868 13398
rect 29828 12912 29880 12918
rect 29828 12854 29880 12860
rect 29644 12844 29696 12850
rect 29644 12786 29696 12792
rect 29656 11014 29684 12786
rect 30024 12434 30052 14991
rect 30196 14952 30248 14958
rect 30196 14894 30248 14900
rect 30104 14408 30156 14414
rect 30104 14350 30156 14356
rect 29932 12406 30052 12434
rect 29932 12238 29960 12406
rect 29920 12232 29972 12238
rect 30116 12186 30144 14350
rect 30208 13734 30236 14894
rect 30300 13818 30328 17274
rect 30748 16108 30800 16114
rect 30748 16050 30800 16056
rect 30300 13790 30604 13818
rect 30196 13728 30248 13734
rect 30196 13670 30248 13676
rect 30472 13728 30524 13734
rect 30472 13670 30524 13676
rect 29920 12174 29972 12180
rect 30024 12158 30144 12186
rect 29736 11824 29788 11830
rect 29734 11792 29736 11801
rect 29788 11792 29790 11801
rect 29734 11727 29790 11736
rect 29828 11756 29880 11762
rect 29828 11698 29880 11704
rect 29840 11234 29868 11698
rect 29920 11280 29972 11286
rect 29840 11228 29920 11234
rect 29840 11222 29972 11228
rect 29736 11212 29788 11218
rect 29736 11154 29788 11160
rect 29840 11206 29960 11222
rect 29644 11008 29696 11014
rect 29644 10950 29696 10956
rect 29656 10266 29684 10950
rect 29748 10742 29776 11154
rect 29840 10810 29868 11206
rect 29920 11144 29972 11150
rect 29920 11086 29972 11092
rect 29828 10804 29880 10810
rect 29828 10746 29880 10752
rect 29736 10736 29788 10742
rect 29736 10678 29788 10684
rect 29932 10538 29960 11086
rect 29920 10532 29972 10538
rect 29920 10474 29972 10480
rect 29644 10260 29696 10266
rect 29644 10202 29696 10208
rect 29644 10056 29696 10062
rect 29644 9998 29696 10004
rect 29552 7540 29604 7546
rect 29552 7482 29604 7488
rect 29564 7002 29592 7482
rect 29552 6996 29604 7002
rect 29552 6938 29604 6944
rect 29552 6656 29604 6662
rect 29552 6598 29604 6604
rect 29458 5944 29514 5953
rect 29458 5879 29514 5888
rect 29460 5160 29512 5166
rect 29460 5102 29512 5108
rect 29472 4865 29500 5102
rect 29458 4856 29514 4865
rect 29458 4791 29514 4800
rect 29564 4214 29592 6598
rect 29656 5846 29684 9998
rect 29736 9376 29788 9382
rect 29736 9318 29788 9324
rect 29748 8022 29776 9318
rect 29828 8832 29880 8838
rect 29828 8774 29880 8780
rect 29840 8566 29868 8774
rect 29828 8560 29880 8566
rect 29828 8502 29880 8508
rect 29920 8288 29972 8294
rect 29920 8230 29972 8236
rect 29736 8016 29788 8022
rect 29736 7958 29788 7964
rect 29828 7540 29880 7546
rect 29828 7482 29880 7488
rect 29736 7200 29788 7206
rect 29736 7142 29788 7148
rect 29748 6798 29776 7142
rect 29736 6792 29788 6798
rect 29736 6734 29788 6740
rect 29748 6458 29776 6734
rect 29736 6452 29788 6458
rect 29736 6394 29788 6400
rect 29840 6338 29868 7482
rect 29748 6310 29868 6338
rect 29644 5840 29696 5846
rect 29644 5782 29696 5788
rect 29642 5536 29698 5545
rect 29642 5471 29698 5480
rect 29656 5370 29684 5471
rect 29644 5364 29696 5370
rect 29644 5306 29696 5312
rect 29552 4208 29604 4214
rect 29552 4150 29604 4156
rect 29368 4072 29420 4078
rect 29368 4014 29420 4020
rect 29000 3936 29052 3942
rect 29000 3878 29052 3884
rect 29276 3936 29328 3942
rect 29276 3878 29328 3884
rect 29000 3528 29052 3534
rect 29000 3470 29052 3476
rect 28908 3120 28960 3126
rect 28908 3062 28960 3068
rect 27988 3052 28040 3058
rect 27988 2994 28040 3000
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 27436 2440 27488 2446
rect 27436 2382 27488 2388
rect 26792 2372 26844 2378
rect 26792 2314 26844 2320
rect 26804 2106 26832 2314
rect 26976 2304 27028 2310
rect 26976 2246 27028 2252
rect 26792 2100 26844 2106
rect 26792 2042 26844 2048
rect 26884 2100 26936 2106
rect 26884 2042 26936 2048
rect 26896 1970 26924 2042
rect 26988 1970 27016 2246
rect 26884 1964 26936 1970
rect 26884 1906 26936 1912
rect 26976 1964 27028 1970
rect 26976 1906 27028 1912
rect 27080 800 27108 2382
rect 27712 2372 27764 2378
rect 27712 2314 27764 2320
rect 27724 1766 27752 2314
rect 27712 1760 27764 1766
rect 27712 1702 27764 1708
rect 29012 800 29040 3470
rect 29288 3194 29316 3878
rect 29276 3188 29328 3194
rect 29276 3130 29328 3136
rect 29380 3126 29408 4014
rect 29644 3664 29696 3670
rect 29642 3632 29644 3641
rect 29696 3632 29698 3641
rect 29642 3567 29698 3576
rect 29748 3398 29776 6310
rect 29828 6248 29880 6254
rect 29828 6190 29880 6196
rect 29840 6089 29868 6190
rect 29826 6080 29882 6089
rect 29826 6015 29882 6024
rect 29932 5930 29960 8230
rect 30024 7410 30052 12158
rect 30104 12096 30156 12102
rect 30104 12038 30156 12044
rect 30116 11937 30144 12038
rect 30102 11928 30158 11937
rect 30102 11863 30158 11872
rect 30104 10804 30156 10810
rect 30104 10746 30156 10752
rect 30116 10470 30144 10746
rect 30104 10464 30156 10470
rect 30104 10406 30156 10412
rect 30208 10266 30236 13670
rect 30484 13530 30512 13670
rect 30576 13530 30604 13790
rect 30472 13524 30524 13530
rect 30472 13466 30524 13472
rect 30564 13524 30616 13530
rect 30564 13466 30616 13472
rect 30484 13326 30512 13466
rect 30472 13320 30524 13326
rect 30472 13262 30524 13268
rect 30288 13252 30340 13258
rect 30288 13194 30340 13200
rect 30300 12986 30328 13194
rect 30654 13016 30710 13025
rect 30288 12980 30340 12986
rect 30654 12951 30710 12960
rect 30288 12922 30340 12928
rect 30668 12782 30696 12951
rect 30656 12776 30708 12782
rect 30656 12718 30708 12724
rect 30380 12232 30432 12238
rect 30380 12174 30432 12180
rect 30288 11756 30340 11762
rect 30288 11698 30340 11704
rect 30300 11082 30328 11698
rect 30288 11076 30340 11082
rect 30288 11018 30340 11024
rect 30288 10464 30340 10470
rect 30288 10406 30340 10412
rect 30196 10260 30248 10266
rect 30196 10202 30248 10208
rect 30300 9994 30328 10406
rect 30288 9988 30340 9994
rect 30288 9930 30340 9936
rect 30196 9376 30248 9382
rect 30196 9318 30248 9324
rect 30288 9376 30340 9382
rect 30288 9318 30340 9324
rect 30104 8560 30156 8566
rect 30104 8502 30156 8508
rect 30116 8362 30144 8502
rect 30104 8356 30156 8362
rect 30104 8298 30156 8304
rect 30012 7404 30064 7410
rect 30012 7346 30064 7352
rect 29840 5902 29960 5930
rect 29840 3534 29868 5902
rect 29918 5808 29974 5817
rect 29918 5743 29974 5752
rect 29932 5642 29960 5743
rect 29920 5636 29972 5642
rect 29920 5578 29972 5584
rect 29918 5400 29974 5409
rect 29918 5335 29920 5344
rect 29972 5335 29974 5344
rect 29920 5306 29972 5312
rect 30024 4842 30052 7346
rect 30208 7274 30236 9318
rect 30300 9110 30328 9318
rect 30288 9104 30340 9110
rect 30288 9046 30340 9052
rect 30392 8129 30420 12174
rect 30472 12164 30524 12170
rect 30472 12106 30524 12112
rect 30484 12073 30512 12106
rect 30470 12064 30526 12073
rect 30470 11999 30526 12008
rect 30470 11520 30526 11529
rect 30470 11455 30526 11464
rect 30484 11354 30512 11455
rect 30472 11348 30524 11354
rect 30472 11290 30524 11296
rect 30472 11212 30524 11218
rect 30472 11154 30524 11160
rect 30378 8120 30434 8129
rect 30378 8055 30434 8064
rect 30380 7948 30432 7954
rect 30380 7890 30432 7896
rect 30288 7880 30340 7886
rect 30288 7822 30340 7828
rect 30196 7268 30248 7274
rect 30196 7210 30248 7216
rect 30300 7206 30328 7822
rect 30392 7750 30420 7890
rect 30380 7744 30432 7750
rect 30380 7686 30432 7692
rect 30288 7200 30340 7206
rect 30288 7142 30340 7148
rect 30484 6746 30512 11154
rect 30564 11144 30616 11150
rect 30562 11112 30564 11121
rect 30616 11112 30618 11121
rect 30562 11047 30618 11056
rect 30656 10668 30708 10674
rect 30656 10610 30708 10616
rect 30564 10464 30616 10470
rect 30564 10406 30616 10412
rect 30576 9722 30604 10406
rect 30668 10198 30696 10610
rect 30656 10192 30708 10198
rect 30656 10134 30708 10140
rect 30668 9926 30696 10134
rect 30656 9920 30708 9926
rect 30656 9862 30708 9868
rect 30564 9716 30616 9722
rect 30564 9658 30616 9664
rect 30576 8022 30604 9658
rect 30656 8424 30708 8430
rect 30656 8366 30708 8372
rect 30564 8016 30616 8022
rect 30564 7958 30616 7964
rect 30564 6860 30616 6866
rect 30564 6802 30616 6808
rect 30300 6730 30512 6746
rect 30288 6724 30512 6730
rect 30340 6718 30512 6724
rect 30288 6666 30340 6672
rect 30288 6384 30340 6390
rect 30288 6326 30340 6332
rect 30196 6248 30248 6254
rect 30196 6190 30248 6196
rect 30208 5846 30236 6190
rect 30196 5840 30248 5846
rect 30196 5782 30248 5788
rect 30300 5370 30328 6326
rect 30288 5364 30340 5370
rect 30288 5306 30340 5312
rect 30300 5234 30328 5306
rect 30288 5228 30340 5234
rect 30288 5170 30340 5176
rect 29932 4814 30052 4842
rect 29932 3670 29960 4814
rect 29920 3664 29972 3670
rect 29920 3606 29972 3612
rect 29828 3528 29880 3534
rect 29828 3470 29880 3476
rect 29736 3392 29788 3398
rect 29736 3334 29788 3340
rect 29368 3120 29420 3126
rect 29368 3062 29420 3068
rect 29736 3120 29788 3126
rect 29736 3062 29788 3068
rect 29748 2514 29776 3062
rect 30194 2952 30250 2961
rect 30194 2887 30250 2896
rect 30208 2854 30236 2887
rect 30196 2848 30248 2854
rect 30196 2790 30248 2796
rect 30288 2848 30340 2854
rect 30288 2790 30340 2796
rect 29736 2508 29788 2514
rect 29736 2450 29788 2456
rect 29920 2372 29972 2378
rect 29920 2314 29972 2320
rect 29932 1834 29960 2314
rect 29920 1828 29972 1834
rect 29920 1770 29972 1776
rect 30300 800 30328 2790
rect 30392 2650 30420 6718
rect 30576 6458 30604 6802
rect 30564 6452 30616 6458
rect 30564 6394 30616 6400
rect 30668 5778 30696 8366
rect 30760 7002 30788 16050
rect 33612 15706 33640 19314
rect 34428 18148 34480 18154
rect 34428 18090 34480 18096
rect 34440 16574 34468 18090
rect 34440 16546 34560 16574
rect 33600 15700 33652 15706
rect 33600 15642 33652 15648
rect 31668 15632 31720 15638
rect 31668 15574 31720 15580
rect 31392 15020 31444 15026
rect 31392 14962 31444 14968
rect 31300 14952 31352 14958
rect 31404 14929 31432 14962
rect 31300 14894 31352 14900
rect 31390 14920 31446 14929
rect 31208 14000 31260 14006
rect 31208 13942 31260 13948
rect 31116 13864 31168 13870
rect 31116 13806 31168 13812
rect 31024 13320 31076 13326
rect 31024 13262 31076 13268
rect 30840 11892 30892 11898
rect 30840 11834 30892 11840
rect 30852 9382 30880 11834
rect 30932 11008 30984 11014
rect 30932 10950 30984 10956
rect 30840 9376 30892 9382
rect 30840 9318 30892 9324
rect 30838 9208 30894 9217
rect 30838 9143 30894 9152
rect 30852 8566 30880 9143
rect 30840 8560 30892 8566
rect 30840 8502 30892 8508
rect 30748 6996 30800 7002
rect 30748 6938 30800 6944
rect 30656 5772 30708 5778
rect 30656 5714 30708 5720
rect 30760 4078 30788 6938
rect 30944 6746 30972 10950
rect 31036 9217 31064 13262
rect 31128 11626 31156 13806
rect 31220 11898 31248 13942
rect 31312 13802 31340 14894
rect 31390 14855 31446 14864
rect 31576 14340 31628 14346
rect 31576 14282 31628 14288
rect 31300 13796 31352 13802
rect 31300 13738 31352 13744
rect 31208 11892 31260 11898
rect 31208 11834 31260 11840
rect 31208 11756 31260 11762
rect 31208 11698 31260 11704
rect 31116 11620 31168 11626
rect 31116 11562 31168 11568
rect 31220 11558 31248 11698
rect 31208 11552 31260 11558
rect 31208 11494 31260 11500
rect 31116 9376 31168 9382
rect 31116 9318 31168 9324
rect 31022 9208 31078 9217
rect 31022 9143 31078 9152
rect 31024 9036 31076 9042
rect 31024 8978 31076 8984
rect 31036 8906 31064 8978
rect 31024 8900 31076 8906
rect 31024 8842 31076 8848
rect 31036 8430 31064 8842
rect 31024 8424 31076 8430
rect 31024 8366 31076 8372
rect 31128 7546 31156 9318
rect 31208 8628 31260 8634
rect 31208 8570 31260 8576
rect 31116 7540 31168 7546
rect 31116 7482 31168 7488
rect 31024 7336 31076 7342
rect 31024 7278 31076 7284
rect 31036 6769 31064 7278
rect 31220 6934 31248 8570
rect 31208 6928 31260 6934
rect 31208 6870 31260 6876
rect 30852 6718 30972 6746
rect 31022 6760 31078 6769
rect 30852 4078 30880 6718
rect 31022 6695 31078 6704
rect 30932 6656 30984 6662
rect 31024 6656 31076 6662
rect 30932 6598 30984 6604
rect 31022 6624 31024 6633
rect 31076 6624 31078 6633
rect 30944 6118 30972 6598
rect 31022 6559 31078 6568
rect 31114 6352 31170 6361
rect 31114 6287 31116 6296
rect 31168 6287 31170 6296
rect 31116 6258 31168 6264
rect 30932 6112 30984 6118
rect 30932 6054 30984 6060
rect 31312 5234 31340 13738
rect 31392 13184 31444 13190
rect 31392 13126 31444 13132
rect 31300 5228 31352 5234
rect 31300 5170 31352 5176
rect 31298 5128 31354 5137
rect 31298 5063 31354 5072
rect 31312 4826 31340 5063
rect 31404 4826 31432 13126
rect 31588 12850 31616 14282
rect 31680 13530 31708 15574
rect 33508 15496 33560 15502
rect 33508 15438 33560 15444
rect 31760 15088 31812 15094
rect 31760 15030 31812 15036
rect 31772 14618 31800 15030
rect 32310 14648 32366 14657
rect 31760 14612 31812 14618
rect 32310 14583 32312 14592
rect 31760 14554 31812 14560
rect 32364 14583 32366 14592
rect 32312 14554 32364 14560
rect 32036 14408 32088 14414
rect 32036 14350 32088 14356
rect 31760 13796 31812 13802
rect 31760 13738 31812 13744
rect 31772 13705 31800 13738
rect 31758 13696 31814 13705
rect 31758 13631 31814 13640
rect 31668 13524 31720 13530
rect 31668 13466 31720 13472
rect 31760 13456 31812 13462
rect 31760 13398 31812 13404
rect 31576 12844 31628 12850
rect 31576 12786 31628 12792
rect 31588 12374 31616 12786
rect 31772 12442 31800 13398
rect 31852 12776 31904 12782
rect 31852 12718 31904 12724
rect 31760 12436 31812 12442
rect 31864 12434 31892 12718
rect 31864 12406 31984 12434
rect 31760 12378 31812 12384
rect 31576 12368 31628 12374
rect 31576 12310 31628 12316
rect 31668 12232 31720 12238
rect 31668 12174 31720 12180
rect 31680 11218 31708 12174
rect 31852 11688 31904 11694
rect 31852 11630 31904 11636
rect 31864 11354 31892 11630
rect 31852 11348 31904 11354
rect 31852 11290 31904 11296
rect 31668 11212 31720 11218
rect 31668 11154 31720 11160
rect 31956 8906 31984 12406
rect 31944 8900 31996 8906
rect 31944 8842 31996 8848
rect 31956 8566 31984 8842
rect 31944 8560 31996 8566
rect 31944 8502 31996 8508
rect 31668 8084 31720 8090
rect 31668 8026 31720 8032
rect 31680 7546 31708 8026
rect 31668 7540 31720 7546
rect 31668 7482 31720 7488
rect 31680 7206 31708 7482
rect 31668 7200 31720 7206
rect 31668 7142 31720 7148
rect 31680 6730 31708 7142
rect 31760 6996 31812 7002
rect 31760 6938 31812 6944
rect 31668 6724 31720 6730
rect 31668 6666 31720 6672
rect 31482 6080 31538 6089
rect 31482 6015 31538 6024
rect 31496 5914 31524 6015
rect 31484 5908 31536 5914
rect 31484 5850 31536 5856
rect 31680 5778 31708 6666
rect 31668 5772 31720 5778
rect 31668 5714 31720 5720
rect 31574 5264 31630 5273
rect 31574 5199 31630 5208
rect 31588 5030 31616 5199
rect 31576 5024 31628 5030
rect 31576 4966 31628 4972
rect 31300 4820 31352 4826
rect 31300 4762 31352 4768
rect 31392 4820 31444 4826
rect 31392 4762 31444 4768
rect 31300 4684 31352 4690
rect 31300 4626 31352 4632
rect 31312 4214 31340 4626
rect 31300 4208 31352 4214
rect 31300 4150 31352 4156
rect 30748 4072 30800 4078
rect 30748 4014 30800 4020
rect 30840 4072 30892 4078
rect 30840 4014 30892 4020
rect 31116 4072 31168 4078
rect 31116 4014 31168 4020
rect 30930 3632 30986 3641
rect 30930 3567 30986 3576
rect 30944 3466 30972 3567
rect 30932 3460 30984 3466
rect 30932 3402 30984 3408
rect 30564 3392 30616 3398
rect 30564 3334 30616 3340
rect 30576 2854 30604 3334
rect 30564 2848 30616 2854
rect 30564 2790 30616 2796
rect 31128 2650 31156 4014
rect 31206 3768 31262 3777
rect 31206 3703 31262 3712
rect 31220 3602 31248 3703
rect 31208 3596 31260 3602
rect 31208 3538 31260 3544
rect 31300 3460 31352 3466
rect 31300 3402 31352 3408
rect 31312 2990 31340 3402
rect 31300 2984 31352 2990
rect 31300 2926 31352 2932
rect 30380 2644 30432 2650
rect 30380 2586 30432 2592
rect 31116 2644 31168 2650
rect 31116 2586 31168 2592
rect 31298 2544 31354 2553
rect 31404 2514 31432 4762
rect 31680 4622 31708 5714
rect 31668 4616 31720 4622
rect 31668 4558 31720 4564
rect 31680 4146 31708 4558
rect 31484 4140 31536 4146
rect 31484 4082 31536 4088
rect 31668 4140 31720 4146
rect 31668 4082 31720 4088
rect 31496 3602 31524 4082
rect 31668 3732 31720 3738
rect 31668 3674 31720 3680
rect 31576 3664 31628 3670
rect 31576 3606 31628 3612
rect 31484 3596 31536 3602
rect 31484 3538 31536 3544
rect 31496 3126 31524 3538
rect 31588 3466 31616 3606
rect 31576 3460 31628 3466
rect 31576 3402 31628 3408
rect 31680 3233 31708 3674
rect 31666 3224 31722 3233
rect 31666 3159 31722 3168
rect 31484 3120 31536 3126
rect 31484 3062 31536 3068
rect 31496 2990 31524 3062
rect 31772 3058 31800 6938
rect 32048 6066 32076 14350
rect 32588 13932 32640 13938
rect 32588 13874 32640 13880
rect 32128 13320 32180 13326
rect 32128 13262 32180 13268
rect 31956 6038 32076 6066
rect 31956 5409 31984 6038
rect 31942 5400 31998 5409
rect 31942 5335 31998 5344
rect 31956 3738 31984 5335
rect 32036 5296 32088 5302
rect 32036 5238 32088 5244
rect 32048 4593 32076 5238
rect 32034 4584 32090 4593
rect 32034 4519 32090 4528
rect 32140 4010 32168 13262
rect 32402 12336 32458 12345
rect 32402 12271 32404 12280
rect 32456 12271 32458 12280
rect 32404 12242 32456 12248
rect 32404 10464 32456 10470
rect 32404 10406 32456 10412
rect 32416 10062 32444 10406
rect 32312 10056 32364 10062
rect 32312 9998 32364 10004
rect 32404 10056 32456 10062
rect 32404 9998 32456 10004
rect 32324 8650 32352 9998
rect 32496 9716 32548 9722
rect 32496 9658 32548 9664
rect 32324 8622 32444 8650
rect 32220 8560 32272 8566
rect 32272 8508 32352 8514
rect 32220 8502 32352 8508
rect 32232 8486 32352 8502
rect 32324 5030 32352 8486
rect 32312 5024 32364 5030
rect 32312 4966 32364 4972
rect 32218 4856 32274 4865
rect 32218 4791 32220 4800
rect 32272 4791 32274 4800
rect 32220 4762 32272 4768
rect 32128 4004 32180 4010
rect 32128 3946 32180 3952
rect 31944 3732 31996 3738
rect 31944 3674 31996 3680
rect 32036 3732 32088 3738
rect 32036 3674 32088 3680
rect 32048 3641 32076 3674
rect 32312 3664 32364 3670
rect 32034 3632 32090 3641
rect 32034 3567 32090 3576
rect 32310 3632 32312 3641
rect 32364 3632 32366 3641
rect 32310 3567 32366 3576
rect 32416 3233 32444 8622
rect 32508 7449 32536 9658
rect 32494 7440 32550 7449
rect 32494 7375 32550 7384
rect 32600 6202 32628 13874
rect 33520 13734 33548 15438
rect 33508 13728 33560 13734
rect 33508 13670 33560 13676
rect 32864 13320 32916 13326
rect 32864 13262 32916 13268
rect 32876 11014 32904 13262
rect 32956 12912 33008 12918
rect 32954 12880 32956 12889
rect 33008 12880 33010 12889
rect 32954 12815 33010 12824
rect 33600 12844 33652 12850
rect 33600 12786 33652 12792
rect 33416 11756 33468 11762
rect 33416 11698 33468 11704
rect 32864 11008 32916 11014
rect 32864 10950 32916 10956
rect 32678 10024 32734 10033
rect 32678 9959 32734 9968
rect 32692 6458 32720 9959
rect 32956 9648 33008 9654
rect 32956 9590 33008 9596
rect 32772 9444 32824 9450
rect 32772 9386 32824 9392
rect 32784 8634 32812 9386
rect 32864 9376 32916 9382
rect 32864 9318 32916 9324
rect 32876 8974 32904 9318
rect 32864 8968 32916 8974
rect 32864 8910 32916 8916
rect 32876 8838 32904 8910
rect 32864 8832 32916 8838
rect 32864 8774 32916 8780
rect 32772 8628 32824 8634
rect 32772 8570 32824 8576
rect 32876 8498 32904 8774
rect 32864 8492 32916 8498
rect 32864 8434 32916 8440
rect 32876 8294 32904 8434
rect 32864 8288 32916 8294
rect 32864 8230 32916 8236
rect 32968 7478 32996 9590
rect 33048 7812 33100 7818
rect 33048 7754 33100 7760
rect 32956 7472 33008 7478
rect 32956 7414 33008 7420
rect 32864 7200 32916 7206
rect 32862 7168 32864 7177
rect 32916 7168 32918 7177
rect 32862 7103 32918 7112
rect 33060 6798 33088 7754
rect 33324 6928 33376 6934
rect 33324 6870 33376 6876
rect 33048 6792 33100 6798
rect 33048 6734 33100 6740
rect 33336 6458 33364 6870
rect 32680 6452 32732 6458
rect 32680 6394 32732 6400
rect 33324 6452 33376 6458
rect 33324 6394 33376 6400
rect 33140 6316 33192 6322
rect 33140 6258 33192 6264
rect 32600 6174 32720 6202
rect 32588 6112 32640 6118
rect 32588 6054 32640 6060
rect 32600 5778 32628 6054
rect 32588 5772 32640 5778
rect 32588 5714 32640 5720
rect 32496 5568 32548 5574
rect 32496 5510 32548 5516
rect 32508 4554 32536 5510
rect 32496 4548 32548 4554
rect 32496 4490 32548 4496
rect 32588 4072 32640 4078
rect 32588 4014 32640 4020
rect 32402 3224 32458 3233
rect 32220 3188 32272 3194
rect 32402 3159 32458 3168
rect 32220 3130 32272 3136
rect 31760 3052 31812 3058
rect 31760 2994 31812 3000
rect 31484 2984 31536 2990
rect 31484 2926 31536 2932
rect 31772 2922 31800 2994
rect 31760 2916 31812 2922
rect 31760 2858 31812 2864
rect 31298 2479 31354 2488
rect 31392 2508 31444 2514
rect 31312 2378 31340 2479
rect 31392 2450 31444 2456
rect 31300 2372 31352 2378
rect 31300 2314 31352 2320
rect 32232 800 32260 3130
rect 32600 2582 32628 4014
rect 32692 3126 32720 6174
rect 32956 6112 33008 6118
rect 32956 6054 33008 6060
rect 32968 5710 32996 6054
rect 33152 5710 33180 6258
rect 33324 5908 33376 5914
rect 33324 5850 33376 5856
rect 32956 5704 33008 5710
rect 32956 5646 33008 5652
rect 33140 5704 33192 5710
rect 33140 5646 33192 5652
rect 33152 5001 33180 5646
rect 33138 4992 33194 5001
rect 33138 4927 33194 4936
rect 33140 4072 33192 4078
rect 33140 4014 33192 4020
rect 32680 3120 32732 3126
rect 32680 3062 32732 3068
rect 33152 2774 33180 4014
rect 33232 3732 33284 3738
rect 33232 3674 33284 3680
rect 33244 3346 33272 3674
rect 33336 3466 33364 5850
rect 33428 3466 33456 11698
rect 33508 6792 33560 6798
rect 33508 6734 33560 6740
rect 33520 6458 33548 6734
rect 33508 6452 33560 6458
rect 33508 6394 33560 6400
rect 33508 4752 33560 4758
rect 33508 4694 33560 4700
rect 33324 3460 33376 3466
rect 33324 3402 33376 3408
rect 33416 3460 33468 3466
rect 33416 3402 33468 3408
rect 33520 3346 33548 4694
rect 33244 3318 33548 3346
rect 33612 2774 33640 12786
rect 34428 12232 34480 12238
rect 34428 12174 34480 12180
rect 33876 11076 33928 11082
rect 33876 11018 33928 11024
rect 33692 10668 33744 10674
rect 33692 10610 33744 10616
rect 33704 7002 33732 10610
rect 33888 10470 33916 11018
rect 34440 10674 34468 12174
rect 34532 11082 34560 16546
rect 34808 11354 34836 37062
rect 36280 36922 36308 37062
rect 36464 36922 36492 37130
rect 37384 37126 37412 39200
rect 38198 37496 38254 37505
rect 38198 37431 38254 37440
rect 37372 37120 37424 37126
rect 37372 37062 37424 37068
rect 38212 36922 38240 37431
rect 36268 36916 36320 36922
rect 36268 36858 36320 36864
rect 36452 36916 36504 36922
rect 36452 36858 36504 36864
rect 38200 36916 38252 36922
rect 38200 36858 38252 36864
rect 35532 36780 35584 36786
rect 35532 36722 35584 36728
rect 37280 36780 37332 36786
rect 37280 36722 37332 36728
rect 35544 36582 35572 36722
rect 35532 36576 35584 36582
rect 35532 36518 35584 36524
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35544 13802 35572 36518
rect 37292 30122 37320 36722
rect 38672 36378 38700 39200
rect 38660 36372 38712 36378
rect 38660 36314 38712 36320
rect 37372 36168 37424 36174
rect 37372 36110 37424 36116
rect 37384 35630 37412 36110
rect 37372 35624 37424 35630
rect 37372 35566 37424 35572
rect 38292 35624 38344 35630
rect 38292 35566 38344 35572
rect 37280 30116 37332 30122
rect 37280 30058 37332 30064
rect 37384 27470 37412 35566
rect 38304 35465 38332 35566
rect 38290 35456 38346 35465
rect 38290 35391 38346 35400
rect 38304 35290 38332 35391
rect 38292 35284 38344 35290
rect 38292 35226 38344 35232
rect 38198 33416 38254 33425
rect 38198 33351 38200 33360
rect 38252 33351 38254 33360
rect 38200 33322 38252 33328
rect 38292 32360 38344 32366
rect 38292 32302 38344 32308
rect 38304 32065 38332 32302
rect 38290 32056 38346 32065
rect 38290 31991 38292 32000
rect 38344 31991 38346 32000
rect 38292 31962 38344 31968
rect 38200 30252 38252 30258
rect 38200 30194 38252 30200
rect 38108 30048 38160 30054
rect 38212 30025 38240 30194
rect 38108 29990 38160 29996
rect 38198 30016 38254 30025
rect 37924 27940 37976 27946
rect 37924 27882 37976 27888
rect 37372 27464 37424 27470
rect 37372 27406 37424 27412
rect 37832 24744 37884 24750
rect 37832 24686 37884 24692
rect 35992 22636 36044 22642
rect 35992 22578 36044 22584
rect 36004 21690 36032 22578
rect 35992 21684 36044 21690
rect 35992 21626 36044 21632
rect 37844 15502 37872 24686
rect 37936 16522 37964 27882
rect 38016 21548 38068 21554
rect 38016 21490 38068 21496
rect 38028 20330 38056 21490
rect 38016 20324 38068 20330
rect 38016 20266 38068 20272
rect 37924 16516 37976 16522
rect 37924 16458 37976 16464
rect 38016 16108 38068 16114
rect 38016 16050 38068 16056
rect 38028 15706 38056 16050
rect 38016 15700 38068 15706
rect 38016 15642 38068 15648
rect 37832 15496 37884 15502
rect 37832 15438 37884 15444
rect 37740 15428 37792 15434
rect 37740 15370 37792 15376
rect 37372 14068 37424 14074
rect 37372 14010 37424 14016
rect 35532 13796 35584 13802
rect 35532 13738 35584 13744
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 37384 12434 37412 14010
rect 37648 12640 37700 12646
rect 37648 12582 37700 12588
rect 37292 12406 37412 12434
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34796 11348 34848 11354
rect 34796 11290 34848 11296
rect 34520 11076 34572 11082
rect 34520 11018 34572 11024
rect 35808 11076 35860 11082
rect 35808 11018 35860 11024
rect 36084 11076 36136 11082
rect 36084 11018 36136 11024
rect 36820 11076 36872 11082
rect 36820 11018 36872 11024
rect 36912 11076 36964 11082
rect 36912 11018 36964 11024
rect 35716 11008 35768 11014
rect 35716 10950 35768 10956
rect 34428 10668 34480 10674
rect 34428 10610 34480 10616
rect 33876 10464 33928 10470
rect 33876 10406 33928 10412
rect 33888 7970 33916 10406
rect 34060 10124 34112 10130
rect 34060 10066 34112 10072
rect 33888 7942 34008 7970
rect 33784 7744 33836 7750
rect 33784 7686 33836 7692
rect 33692 6996 33744 7002
rect 33692 6938 33744 6944
rect 33796 5302 33824 7686
rect 33784 5296 33836 5302
rect 33784 5238 33836 5244
rect 33692 5160 33744 5166
rect 33796 5137 33824 5238
rect 33692 5102 33744 5108
rect 33782 5128 33838 5137
rect 33152 2746 33364 2774
rect 32588 2576 32640 2582
rect 32588 2518 32640 2524
rect 33336 2378 33364 2746
rect 33520 2746 33640 2774
rect 33324 2372 33376 2378
rect 33324 2314 33376 2320
rect 32404 2032 32456 2038
rect 32404 1974 32456 1980
rect 32416 1698 32444 1974
rect 33520 1766 33548 2746
rect 33704 2378 33732 5102
rect 33782 5063 33838 5072
rect 33784 4480 33836 4486
rect 33784 4422 33836 4428
rect 33796 3942 33824 4422
rect 33876 4276 33928 4282
rect 33876 4218 33928 4224
rect 33888 4146 33916 4218
rect 33876 4140 33928 4146
rect 33876 4082 33928 4088
rect 33784 3936 33836 3942
rect 33784 3878 33836 3884
rect 33876 3936 33928 3942
rect 33876 3878 33928 3884
rect 33784 3664 33836 3670
rect 33782 3632 33784 3641
rect 33836 3632 33838 3641
rect 33782 3567 33838 3576
rect 33888 3466 33916 3878
rect 33876 3460 33928 3466
rect 33876 3402 33928 3408
rect 33980 2774 34008 7942
rect 34072 6798 34100 10066
rect 34440 9194 34468 10610
rect 34704 10600 34756 10606
rect 34704 10542 34756 10548
rect 34348 9166 34468 9194
rect 34060 6792 34112 6798
rect 34060 6734 34112 6740
rect 34244 6180 34296 6186
rect 34244 6122 34296 6128
rect 34150 5944 34206 5953
rect 34150 5879 34206 5888
rect 34164 5710 34192 5879
rect 34152 5704 34204 5710
rect 34152 5646 34204 5652
rect 34152 5228 34204 5234
rect 34152 5170 34204 5176
rect 34060 5160 34112 5166
rect 34060 5102 34112 5108
rect 34072 3602 34100 5102
rect 34164 4622 34192 5170
rect 34152 4616 34204 4622
rect 34152 4558 34204 4564
rect 34152 3936 34204 3942
rect 34152 3878 34204 3884
rect 34060 3596 34112 3602
rect 34060 3538 34112 3544
rect 33796 2746 34008 2774
rect 33796 2514 33824 2746
rect 34072 2514 34100 3538
rect 34164 3369 34192 3878
rect 34256 3738 34284 6122
rect 34348 5234 34376 9166
rect 34428 8832 34480 8838
rect 34428 8774 34480 8780
rect 34440 6390 34468 8774
rect 34612 8288 34664 8294
rect 34612 8230 34664 8236
rect 34624 8090 34652 8230
rect 34612 8084 34664 8090
rect 34612 8026 34664 8032
rect 34520 6656 34572 6662
rect 34520 6598 34572 6604
rect 34428 6384 34480 6390
rect 34428 6326 34480 6332
rect 34532 5522 34560 6598
rect 34610 6488 34666 6497
rect 34610 6423 34612 6432
rect 34664 6423 34666 6432
rect 34612 6394 34664 6400
rect 34612 6316 34664 6322
rect 34612 6258 34664 6264
rect 34624 6186 34652 6258
rect 34612 6180 34664 6186
rect 34612 6122 34664 6128
rect 34440 5494 34560 5522
rect 34336 5228 34388 5234
rect 34336 5170 34388 5176
rect 34440 5166 34468 5494
rect 34518 5264 34574 5273
rect 34518 5199 34520 5208
rect 34572 5199 34574 5208
rect 34520 5170 34572 5176
rect 34428 5160 34480 5166
rect 34428 5102 34480 5108
rect 34336 5092 34388 5098
rect 34336 5034 34388 5040
rect 34244 3732 34296 3738
rect 34244 3674 34296 3680
rect 34244 3528 34296 3534
rect 34244 3470 34296 3476
rect 34150 3360 34206 3369
rect 34150 3295 34206 3304
rect 34256 2961 34284 3470
rect 34242 2952 34298 2961
rect 34348 2922 34376 5034
rect 34624 4622 34652 6122
rect 34612 4616 34664 4622
rect 34612 4558 34664 4564
rect 34612 4140 34664 4146
rect 34612 4082 34664 4088
rect 34520 4004 34572 4010
rect 34520 3946 34572 3952
rect 34532 3505 34560 3946
rect 34518 3496 34574 3505
rect 34518 3431 34574 3440
rect 34426 3224 34482 3233
rect 34624 3210 34652 4082
rect 34716 3942 34744 10542
rect 35624 10532 35676 10538
rect 35624 10474 35676 10480
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34980 9920 35032 9926
rect 34980 9862 35032 9868
rect 35440 9920 35492 9926
rect 35440 9862 35492 9868
rect 34992 9450 35020 9862
rect 34980 9444 35032 9450
rect 34980 9386 35032 9392
rect 35348 9444 35400 9450
rect 35348 9386 35400 9392
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 35360 8906 35388 9386
rect 34796 8900 34848 8906
rect 34796 8842 34848 8848
rect 35348 8900 35400 8906
rect 35348 8842 35400 8848
rect 34808 6458 34836 8842
rect 35360 8362 35388 8842
rect 35348 8356 35400 8362
rect 35348 8298 35400 8304
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34888 6792 34940 6798
rect 34888 6734 34940 6740
rect 34796 6452 34848 6458
rect 34796 6394 34848 6400
rect 34900 6338 34928 6734
rect 35360 6730 35388 8298
rect 35348 6724 35400 6730
rect 35348 6666 35400 6672
rect 34808 6310 34928 6338
rect 34808 6118 34836 6310
rect 34796 6112 34848 6118
rect 34796 6054 34848 6060
rect 34808 5234 34836 6054
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35072 5704 35124 5710
rect 35072 5646 35124 5652
rect 35084 5234 35112 5646
rect 34796 5228 34848 5234
rect 34796 5170 34848 5176
rect 35072 5228 35124 5234
rect 35072 5170 35124 5176
rect 34808 4740 34836 5170
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34808 4712 34928 4740
rect 34900 4214 34928 4712
rect 34980 4480 35032 4486
rect 34978 4448 34980 4457
rect 35348 4480 35400 4486
rect 35032 4448 35034 4457
rect 35348 4422 35400 4428
rect 34978 4383 35034 4392
rect 34888 4208 34940 4214
rect 34888 4150 34940 4156
rect 34980 4140 35032 4146
rect 34980 4082 35032 4088
rect 34992 4026 35020 4082
rect 34808 3998 35020 4026
rect 34704 3936 34756 3942
rect 34704 3878 34756 3884
rect 34808 3777 34836 3998
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34794 3768 34850 3777
rect 34934 3771 35242 3780
rect 34794 3703 34850 3712
rect 34980 3392 35032 3398
rect 34980 3334 35032 3340
rect 34426 3159 34482 3168
rect 34532 3182 34652 3210
rect 34440 2922 34468 3159
rect 34242 2887 34298 2896
rect 34336 2916 34388 2922
rect 34336 2858 34388 2864
rect 34428 2916 34480 2922
rect 34428 2858 34480 2864
rect 34532 2854 34560 3182
rect 34992 3097 35020 3334
rect 34978 3088 35034 3097
rect 34612 3052 34664 3058
rect 34978 3023 35034 3032
rect 34612 2994 34664 3000
rect 34244 2848 34296 2854
rect 34244 2790 34296 2796
rect 34520 2848 34572 2854
rect 34520 2790 34572 2796
rect 33784 2508 33836 2514
rect 33784 2450 33836 2456
rect 34060 2508 34112 2514
rect 34060 2450 34112 2456
rect 33692 2372 33744 2378
rect 33692 2314 33744 2320
rect 34152 2304 34204 2310
rect 34152 2246 34204 2252
rect 33508 1760 33560 1766
rect 33508 1702 33560 1708
rect 32404 1692 32456 1698
rect 32404 1634 32456 1640
rect 34164 800 34192 2246
rect 34256 1766 34284 2790
rect 34244 1760 34296 1766
rect 34244 1702 34296 1708
rect 34624 1698 34652 2994
rect 34704 2848 34756 2854
rect 34704 2790 34756 2796
rect 34716 2650 34744 2790
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34704 2644 34756 2650
rect 34704 2586 34756 2592
rect 35360 1970 35388 4422
rect 35452 4146 35480 9862
rect 35636 9674 35664 10474
rect 35728 10470 35756 10950
rect 35716 10464 35768 10470
rect 35716 10406 35768 10412
rect 35728 9994 35756 10406
rect 35716 9988 35768 9994
rect 35716 9930 35768 9936
rect 35636 9646 35756 9674
rect 35728 9382 35756 9646
rect 35716 9376 35768 9382
rect 35716 9318 35768 9324
rect 35728 8838 35756 9318
rect 35716 8832 35768 8838
rect 35716 8774 35768 8780
rect 35716 8492 35768 8498
rect 35716 8434 35768 8440
rect 35624 7880 35676 7886
rect 35624 7822 35676 7828
rect 35532 6792 35584 6798
rect 35532 6734 35584 6740
rect 35544 6186 35572 6734
rect 35636 6390 35664 7822
rect 35728 7546 35756 8434
rect 35716 7540 35768 7546
rect 35716 7482 35768 7488
rect 35820 7426 35848 11018
rect 35728 7398 35848 7426
rect 35624 6384 35676 6390
rect 35624 6326 35676 6332
rect 35532 6180 35584 6186
rect 35532 6122 35584 6128
rect 35440 4140 35492 4146
rect 35440 4082 35492 4088
rect 35624 3392 35676 3398
rect 35624 3334 35676 3340
rect 35440 2304 35492 2310
rect 35440 2246 35492 2252
rect 35348 1964 35400 1970
rect 35348 1906 35400 1912
rect 34612 1692 34664 1698
rect 34612 1634 34664 1640
rect 35452 800 35480 2246
rect 35636 2106 35664 3334
rect 35728 2774 35756 7398
rect 35808 5704 35860 5710
rect 35808 5646 35860 5652
rect 35820 4622 35848 5646
rect 35900 5024 35952 5030
rect 35900 4966 35952 4972
rect 35912 4690 35940 4966
rect 35900 4684 35952 4690
rect 35900 4626 35952 4632
rect 35808 4616 35860 4622
rect 35808 4558 35860 4564
rect 35820 4146 35848 4558
rect 35992 4480 36044 4486
rect 35992 4422 36044 4428
rect 35808 4140 35860 4146
rect 35808 4082 35860 4088
rect 35820 3058 35848 4082
rect 35900 3936 35952 3942
rect 35900 3878 35952 3884
rect 35808 3052 35860 3058
rect 35808 2994 35860 3000
rect 35728 2746 35848 2774
rect 35820 2514 35848 2746
rect 35808 2508 35860 2514
rect 35808 2450 35860 2456
rect 35624 2100 35676 2106
rect 35624 2042 35676 2048
rect 35912 1902 35940 3878
rect 36004 3466 36032 4422
rect 35992 3460 36044 3466
rect 35992 3402 36044 3408
rect 36096 3194 36124 11018
rect 36268 9648 36320 9654
rect 36268 9590 36320 9596
rect 36280 9178 36308 9590
rect 36268 9172 36320 9178
rect 36268 9114 36320 9120
rect 36280 8090 36308 9114
rect 36268 8084 36320 8090
rect 36268 8026 36320 8032
rect 36280 6254 36308 8026
rect 36542 6760 36598 6769
rect 36542 6695 36598 6704
rect 36556 6458 36584 6695
rect 36636 6656 36688 6662
rect 36636 6598 36688 6604
rect 36544 6452 36596 6458
rect 36544 6394 36596 6400
rect 36648 6322 36676 6598
rect 36636 6316 36688 6322
rect 36636 6258 36688 6264
rect 36268 6248 36320 6254
rect 36268 6190 36320 6196
rect 36280 5710 36308 6190
rect 36268 5704 36320 5710
rect 36268 5646 36320 5652
rect 36280 5234 36308 5646
rect 36268 5228 36320 5234
rect 36268 5170 36320 5176
rect 36280 4604 36308 5170
rect 36544 5024 36596 5030
rect 36544 4966 36596 4972
rect 36360 4616 36412 4622
rect 36280 4576 36360 4604
rect 36360 4558 36412 4564
rect 36372 4214 36400 4558
rect 36556 4282 36584 4966
rect 36544 4276 36596 4282
rect 36544 4218 36596 4224
rect 36360 4208 36412 4214
rect 36360 4150 36412 4156
rect 36648 4010 36676 6258
rect 36636 4004 36688 4010
rect 36636 3946 36688 3952
rect 36176 3936 36228 3942
rect 36176 3878 36228 3884
rect 36084 3188 36136 3194
rect 36084 3130 36136 3136
rect 36096 3058 36124 3130
rect 36084 3052 36136 3058
rect 36084 2994 36136 3000
rect 36188 2553 36216 3878
rect 36648 3534 36676 3946
rect 36832 3670 36860 11018
rect 36924 10266 36952 11018
rect 36912 10260 36964 10266
rect 36912 10202 36964 10208
rect 36924 9654 36952 10202
rect 37292 9722 37320 12406
rect 37556 12164 37608 12170
rect 37556 12106 37608 12112
rect 37372 11552 37424 11558
rect 37372 11494 37424 11500
rect 37280 9716 37332 9722
rect 37280 9658 37332 9664
rect 36912 9648 36964 9654
rect 36912 9590 36964 9596
rect 37280 9512 37332 9518
rect 37280 9454 37332 9460
rect 37292 8838 37320 9454
rect 37280 8832 37332 8838
rect 37280 8774 37332 8780
rect 37292 8294 37320 8774
rect 37280 8288 37332 8294
rect 37280 8230 37332 8236
rect 37188 8084 37240 8090
rect 37188 8026 37240 8032
rect 37200 7546 37228 8026
rect 37292 7750 37320 8230
rect 37280 7744 37332 7750
rect 37280 7686 37332 7692
rect 37188 7540 37240 7546
rect 37188 7482 37240 7488
rect 37292 7410 37320 7686
rect 37280 7404 37332 7410
rect 37280 7346 37332 7352
rect 37292 6798 37320 7346
rect 37280 6792 37332 6798
rect 37280 6734 37332 6740
rect 37292 5710 37320 6734
rect 37280 5704 37332 5710
rect 37280 5646 37332 5652
rect 37280 5568 37332 5574
rect 37280 5510 37332 5516
rect 37004 4480 37056 4486
rect 37004 4422 37056 4428
rect 36820 3664 36872 3670
rect 36820 3606 36872 3612
rect 36832 3534 36860 3606
rect 36636 3528 36688 3534
rect 36636 3470 36688 3476
rect 36820 3528 36872 3534
rect 36820 3470 36872 3476
rect 36268 3392 36320 3398
rect 36268 3334 36320 3340
rect 36174 2544 36230 2553
rect 36174 2479 36230 2488
rect 36280 2417 36308 3334
rect 36636 2848 36688 2854
rect 36636 2790 36688 2796
rect 36648 2446 36676 2790
rect 36636 2440 36688 2446
rect 36266 2408 36322 2417
rect 36636 2382 36688 2388
rect 36266 2343 36322 2352
rect 35900 1896 35952 1902
rect 35900 1838 35952 1844
rect 37016 1834 37044 4422
rect 37292 3126 37320 5510
rect 37280 3120 37332 3126
rect 37280 3062 37332 3068
rect 37384 3058 37412 11494
rect 37568 6322 37596 12106
rect 37660 10266 37688 12582
rect 37648 10260 37700 10266
rect 37648 10202 37700 10208
rect 37660 9382 37688 10202
rect 37648 9376 37700 9382
rect 37648 9318 37700 9324
rect 37556 6316 37608 6322
rect 37556 6258 37608 6264
rect 37556 5024 37608 5030
rect 37556 4966 37608 4972
rect 37568 3602 37596 4966
rect 37648 4616 37700 4622
rect 37648 4558 37700 4564
rect 37660 4010 37688 4558
rect 37648 4004 37700 4010
rect 37648 3946 37700 3952
rect 37556 3596 37608 3602
rect 37556 3538 37608 3544
rect 37568 3398 37596 3538
rect 37556 3392 37608 3398
rect 37556 3334 37608 3340
rect 37568 3194 37596 3334
rect 37556 3188 37608 3194
rect 37556 3130 37608 3136
rect 37752 3126 37780 15370
rect 38120 14618 38148 29990
rect 38198 29951 38254 29960
rect 38200 28076 38252 28082
rect 38200 28018 38252 28024
rect 38212 27985 38240 28018
rect 38198 27976 38254 27985
rect 38198 27911 38254 27920
rect 38292 26920 38344 26926
rect 38292 26862 38344 26868
rect 38304 26625 38332 26862
rect 38290 26616 38346 26625
rect 38290 26551 38292 26560
rect 38344 26551 38346 26560
rect 38292 26522 38344 26528
rect 38292 24744 38344 24750
rect 38292 24686 38344 24692
rect 38304 24585 38332 24686
rect 38290 24576 38346 24585
rect 38290 24511 38346 24520
rect 38304 24410 38332 24511
rect 38292 24404 38344 24410
rect 38292 24346 38344 24352
rect 38198 22536 38254 22545
rect 38198 22471 38200 22480
rect 38252 22471 38254 22480
rect 38200 22442 38252 22448
rect 38200 21344 38252 21350
rect 38200 21286 38252 21292
rect 38212 21185 38240 21286
rect 38198 21176 38254 21185
rect 38198 21111 38254 21120
rect 38200 19168 38252 19174
rect 38198 19136 38200 19145
rect 38252 19136 38254 19145
rect 38198 19071 38254 19080
rect 38292 17128 38344 17134
rect 38290 17096 38292 17105
rect 38344 17096 38346 17105
rect 38290 17031 38346 17040
rect 38304 16794 38332 17031
rect 38292 16788 38344 16794
rect 38292 16730 38344 16736
rect 38200 15904 38252 15910
rect 38200 15846 38252 15852
rect 38212 15745 38240 15846
rect 38198 15736 38254 15745
rect 38198 15671 38254 15680
rect 38108 14612 38160 14618
rect 38108 14554 38160 14560
rect 38292 13932 38344 13938
rect 38292 13874 38344 13880
rect 38304 13705 38332 13874
rect 38290 13696 38346 13705
rect 38290 13631 38346 13640
rect 37832 12096 37884 12102
rect 37832 12038 37884 12044
rect 37924 12096 37976 12102
rect 37924 12038 37976 12044
rect 37740 3120 37792 3126
rect 37740 3062 37792 3068
rect 37372 3052 37424 3058
rect 37372 2994 37424 3000
rect 37188 2304 37240 2310
rect 37188 2246 37240 2252
rect 37004 1828 37056 1834
rect 37004 1770 37056 1776
rect 37200 1465 37228 2246
rect 37186 1456 37242 1465
rect 37186 1391 37242 1400
rect 37384 800 37412 2994
rect 37844 2774 37872 12038
rect 37936 9518 37964 12038
rect 38200 11756 38252 11762
rect 38200 11698 38252 11704
rect 38212 11665 38240 11698
rect 38384 11688 38436 11694
rect 38198 11656 38254 11665
rect 38016 11620 38068 11626
rect 38384 11630 38436 11636
rect 38198 11591 38254 11600
rect 38016 11562 38068 11568
rect 37924 9512 37976 9518
rect 37924 9454 37976 9460
rect 38028 9081 38056 11562
rect 38108 11076 38160 11082
rect 38108 11018 38160 11024
rect 38014 9072 38070 9081
rect 38014 9007 38070 9016
rect 38016 7200 38068 7206
rect 38016 7142 38068 7148
rect 38028 6662 38056 7142
rect 38016 6656 38068 6662
rect 38016 6598 38068 6604
rect 38016 5704 38068 5710
rect 38016 5646 38068 5652
rect 37922 5536 37978 5545
rect 37922 5471 37978 5480
rect 37936 5302 37964 5471
rect 37924 5296 37976 5302
rect 37924 5238 37976 5244
rect 38028 4622 38056 5646
rect 38120 5302 38148 11018
rect 38292 10600 38344 10606
rect 38292 10542 38344 10548
rect 38304 10305 38332 10542
rect 38290 10296 38346 10305
rect 38290 10231 38292 10240
rect 38344 10231 38346 10240
rect 38292 10202 38344 10208
rect 38200 9376 38252 9382
rect 38200 9318 38252 9324
rect 38212 6322 38240 9318
rect 38292 8492 38344 8498
rect 38292 8434 38344 8440
rect 38304 8265 38332 8434
rect 38290 8256 38346 8265
rect 38290 8191 38346 8200
rect 38200 6316 38252 6322
rect 38200 6258 38252 6264
rect 38212 6225 38240 6258
rect 38198 6216 38254 6225
rect 38198 6151 38254 6160
rect 38108 5296 38160 5302
rect 38108 5238 38160 5244
rect 38120 4865 38148 5238
rect 38106 4856 38162 4865
rect 38106 4791 38162 4800
rect 38016 4616 38068 4622
rect 38016 4558 38068 4564
rect 38200 3392 38252 3398
rect 38200 3334 38252 3340
rect 38212 2825 38240 3334
rect 37660 2746 37872 2774
rect 38198 2816 38254 2825
rect 38198 2751 38254 2760
rect 37660 2514 37688 2746
rect 38396 2514 38424 11630
rect 37648 2508 37700 2514
rect 37648 2450 37700 2456
rect 38384 2508 38436 2514
rect 38384 2450 38436 2456
rect 39304 2440 39356 2446
rect 39304 2382 39356 2388
rect 39316 800 39344 2382
rect 18 200 74 800
rect 1306 200 1362 800
rect 3238 200 3294 800
rect 4526 200 4582 800
rect 6458 200 6514 800
rect 8390 200 8446 800
rect 9678 200 9734 800
rect 11610 200 11666 800
rect 13542 200 13598 800
rect 14830 200 14886 800
rect 16762 200 16818 800
rect 18694 200 18750 800
rect 19982 200 20038 800
rect 21914 200 21970 800
rect 23846 200 23902 800
rect 25134 200 25190 800
rect 27066 200 27122 800
rect 28998 200 29054 800
rect 30286 200 30342 800
rect 32218 200 32274 800
rect 34150 200 34206 800
rect 35438 200 35494 800
rect 37370 200 37426 800
rect 39302 200 39358 800
<< via2 >>
rect 2870 39480 2926 39536
rect 1674 37440 1730 37496
rect 1674 36080 1730 36136
rect 1674 34040 1730 34096
rect 1674 32000 1730 32056
rect 1674 30660 1730 30696
rect 1674 30640 1676 30660
rect 1676 30640 1728 30660
rect 1728 30640 1730 30660
rect 1582 28636 1584 28656
rect 1584 28636 1636 28656
rect 1636 28636 1638 28656
rect 1582 28600 1638 28636
rect 1674 26560 1730 26616
rect 1582 25236 1584 25256
rect 1584 25236 1636 25256
rect 1636 25236 1638 25256
rect 1582 25200 1638 25236
rect 1582 23196 1584 23216
rect 1584 23196 1636 23216
rect 1636 23196 1638 23216
rect 1582 23160 1638 23196
rect 1674 21120 1730 21176
rect 1674 19780 1730 19816
rect 1674 19760 1676 19780
rect 1676 19760 1728 19780
rect 1728 19760 1730 19780
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 1674 17720 1730 17776
rect 1674 15680 1730 15736
rect 1582 14356 1584 14376
rect 1584 14356 1636 14376
rect 1636 14356 1638 14376
rect 1582 14320 1638 14356
rect 1674 12280 1730 12336
rect 1674 10240 1730 10296
rect 1674 8900 1730 8936
rect 1674 8880 1676 8900
rect 1676 8880 1728 8900
rect 1728 8880 1730 8900
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 1674 6840 1730 6896
rect 1674 4800 1730 4856
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 1674 3440 1730 3496
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 7838 7384 7894 7440
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4066 2508 4122 2544
rect 4066 2488 4068 2508
rect 4068 2488 4120 2508
rect 4120 2488 4122 2508
rect 12438 5092 12494 5128
rect 12438 5072 12440 5092
rect 12440 5072 12492 5092
rect 12492 5072 12494 5092
rect 12346 4820 12402 4856
rect 12346 4800 12348 4820
rect 12348 4800 12400 4820
rect 12400 4800 12402 4820
rect 12254 4120 12310 4176
rect 2778 1400 2834 1456
rect 16210 15428 16266 15464
rect 16210 15408 16212 15428
rect 16212 15408 16264 15428
rect 16264 15408 16266 15428
rect 14738 13368 14794 13424
rect 14830 10512 14886 10568
rect 14278 9016 14334 9072
rect 14370 5344 14426 5400
rect 15842 12180 15844 12200
rect 15844 12180 15896 12200
rect 15896 12180 15898 12200
rect 15842 12144 15898 12180
rect 15290 9424 15346 9480
rect 16302 11872 16358 11928
rect 15658 10124 15714 10160
rect 15658 10104 15660 10124
rect 15660 10104 15712 10124
rect 15712 10104 15714 10124
rect 15658 9696 15714 9752
rect 15014 5616 15070 5672
rect 16670 12144 16726 12200
rect 16854 12144 16910 12200
rect 16854 10104 16910 10160
rect 16302 9424 16358 9480
rect 16394 8236 16396 8256
rect 16396 8236 16448 8256
rect 16448 8236 16450 8256
rect 16394 8200 16450 8236
rect 16670 9288 16726 9344
rect 17222 13232 17278 13288
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 17222 12824 17278 12880
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19890 18164 19892 18184
rect 19892 18164 19944 18184
rect 19944 18164 19946 18184
rect 19890 18128 19946 18164
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 16578 6568 16634 6624
rect 15842 4564 15844 4584
rect 15844 4564 15896 4584
rect 15896 4564 15898 4584
rect 15842 4528 15898 4564
rect 13726 3476 13728 3496
rect 13728 3476 13780 3496
rect 13780 3476 13782 3496
rect 13726 3440 13782 3476
rect 16670 4564 16672 4584
rect 16672 4564 16724 4584
rect 16724 4564 16726 4584
rect 16670 4528 16726 4564
rect 16118 3984 16174 4040
rect 17774 9832 17830 9888
rect 19062 13232 19118 13288
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 20442 17856 20498 17912
rect 20534 15952 20590 16008
rect 22098 17856 22154 17912
rect 21454 16496 21510 16552
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19982 14068 20038 14104
rect 19982 14048 19984 14068
rect 19984 14048 20036 14068
rect 20036 14048 20038 14068
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 21270 15308 21272 15328
rect 21272 15308 21324 15328
rect 21324 15308 21326 15328
rect 20626 14492 20628 14512
rect 20628 14492 20680 14512
rect 20680 14492 20682 14512
rect 20626 14456 20682 14492
rect 17222 4548 17278 4584
rect 17222 4528 17224 4548
rect 17224 4528 17276 4548
rect 17276 4528 17278 4548
rect 17958 8336 18014 8392
rect 18234 9696 18290 9752
rect 17774 6724 17830 6760
rect 17774 6704 17776 6724
rect 17776 6704 17828 6724
rect 17828 6704 17830 6724
rect 17958 6296 18014 6352
rect 17682 5752 17738 5808
rect 17866 3984 17922 4040
rect 18418 9832 18474 9888
rect 18142 6840 18198 6896
rect 19246 11192 19302 11248
rect 18602 9696 18658 9752
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19798 11756 19854 11792
rect 19798 11736 19800 11756
rect 19800 11736 19852 11756
rect 19852 11736 19854 11756
rect 20626 12416 20682 12472
rect 21270 15272 21326 15308
rect 21086 12144 21142 12200
rect 21638 14048 21694 14104
rect 22282 14456 22338 14512
rect 22006 14356 22008 14376
rect 22008 14356 22060 14376
rect 22060 14356 22062 14376
rect 22006 14320 22062 14356
rect 20994 11464 21050 11520
rect 19798 11056 19854 11112
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 18510 6568 18566 6624
rect 18970 8336 19026 8392
rect 18878 2624 18934 2680
rect 19430 10240 19486 10296
rect 20350 10376 20406 10432
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19982 9596 19984 9616
rect 19984 9596 20036 9616
rect 20036 9596 20038 9616
rect 19982 9560 20038 9596
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19062 7404 19118 7440
rect 19062 7384 19064 7404
rect 19064 7384 19116 7404
rect 19116 7384 19118 7404
rect 19246 6740 19248 6760
rect 19248 6740 19300 6760
rect 19300 6740 19302 6760
rect 19246 6704 19302 6740
rect 20166 8880 20222 8936
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19246 5208 19302 5264
rect 19154 4800 19210 4856
rect 20258 7692 20260 7712
rect 20260 7692 20312 7712
rect 20312 7692 20314 7712
rect 20258 7656 20314 7692
rect 20994 11192 21050 11248
rect 20626 10104 20682 10160
rect 20534 9832 20590 9888
rect 20350 6840 20406 6896
rect 20258 6704 20314 6760
rect 19522 6024 19578 6080
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19430 4664 19486 4720
rect 19062 3984 19118 4040
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19982 3460 20038 3496
rect 19982 3440 19984 3460
rect 19984 3440 20036 3460
rect 20036 3440 20038 3460
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19982 3032 20038 3088
rect 20718 8472 20774 8528
rect 20442 5616 20498 5672
rect 20626 5344 20682 5400
rect 20902 7656 20958 7712
rect 20810 5480 20866 5536
rect 21546 10648 21602 10704
rect 21270 8472 21326 8528
rect 21362 8200 21418 8256
rect 21178 8064 21234 8120
rect 20902 3168 20958 3224
rect 21086 4392 21142 4448
rect 21178 3576 21234 3632
rect 22282 13776 22338 13832
rect 22098 10920 22154 10976
rect 21914 10240 21970 10296
rect 22190 10648 22246 10704
rect 21914 10004 21916 10024
rect 21916 10004 21968 10024
rect 21968 10004 21970 10024
rect 21914 9968 21970 10004
rect 21822 9696 21878 9752
rect 23570 17312 23626 17368
rect 23294 13932 23350 13968
rect 23294 13912 23296 13932
rect 23296 13912 23348 13932
rect 23348 13912 23350 13932
rect 21914 9288 21970 9344
rect 22098 9152 22154 9208
rect 22098 8608 22154 8664
rect 22006 8472 22062 8528
rect 21822 8356 21878 8392
rect 21822 8336 21824 8356
rect 21824 8336 21876 8356
rect 21876 8336 21878 8356
rect 22558 9560 22614 9616
rect 21730 7112 21786 7168
rect 21730 6160 21786 6216
rect 22098 7148 22100 7168
rect 22100 7148 22152 7168
rect 22152 7148 22154 7168
rect 22098 7112 22154 7148
rect 21914 6976 21970 7032
rect 22374 6976 22430 7032
rect 22834 11228 22836 11248
rect 22836 11228 22888 11248
rect 22888 11228 22890 11248
rect 22834 11192 22890 11228
rect 22834 10512 22890 10568
rect 23478 11056 23534 11112
rect 22926 9832 22982 9888
rect 22742 9696 22798 9752
rect 23110 8744 23166 8800
rect 22926 8064 22982 8120
rect 22374 6024 22430 6080
rect 21914 5888 21970 5944
rect 22098 5908 22154 5944
rect 22098 5888 22100 5908
rect 22100 5888 22152 5908
rect 22152 5888 22154 5908
rect 22190 5344 22246 5400
rect 21638 5208 21694 5264
rect 23386 8064 23442 8120
rect 21362 2896 21418 2952
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20626 2372 20682 2408
rect 20626 2352 20628 2372
rect 20628 2352 20680 2372
rect 20680 2352 20682 2372
rect 22374 4020 22376 4040
rect 22376 4020 22428 4040
rect 22428 4020 22430 4040
rect 22374 3984 22430 4020
rect 22098 3884 22100 3904
rect 22100 3884 22152 3904
rect 22152 3884 22154 3904
rect 22098 3848 22154 3884
rect 22098 3576 22154 3632
rect 22926 4936 22982 4992
rect 23202 3984 23258 4040
rect 22190 3304 22246 3360
rect 22190 3188 22246 3224
rect 22190 3168 22192 3188
rect 22192 3168 22244 3188
rect 22244 3168 22246 3188
rect 23754 11600 23810 11656
rect 24122 14048 24178 14104
rect 24030 13368 24086 13424
rect 23570 9424 23626 9480
rect 24214 11056 24270 11112
rect 23754 8608 23810 8664
rect 23478 4800 23534 4856
rect 23386 3052 23442 3088
rect 23386 3032 23388 3052
rect 23388 3032 23440 3052
rect 23440 3032 23442 3052
rect 24122 7248 24178 7304
rect 24306 8880 24362 8936
rect 24582 10920 24638 10976
rect 24490 9696 24546 9752
rect 25134 14320 25190 14376
rect 26054 17620 26056 17640
rect 26056 17620 26108 17640
rect 26108 17620 26110 17640
rect 26054 17584 26110 17620
rect 25778 16516 25834 16552
rect 25778 16496 25780 16516
rect 25780 16496 25832 16516
rect 25832 16496 25834 16516
rect 25502 14356 25504 14376
rect 25504 14356 25556 14376
rect 25556 14356 25558 14376
rect 25502 14320 25558 14356
rect 25134 12008 25190 12064
rect 25134 11328 25190 11384
rect 25686 13252 25742 13288
rect 25686 13232 25688 13252
rect 25688 13232 25740 13252
rect 25740 13232 25742 13252
rect 25410 11192 25466 11248
rect 25226 8472 25282 8528
rect 24858 7792 24914 7848
rect 24766 7656 24822 7712
rect 24582 5516 24584 5536
rect 24584 5516 24636 5536
rect 24636 5516 24638 5536
rect 24582 5480 24638 5516
rect 24306 5208 24362 5264
rect 26514 17312 26570 17368
rect 26698 15020 26754 15056
rect 26698 15000 26700 15020
rect 26700 15000 26752 15020
rect 26752 15000 26754 15020
rect 26514 11192 26570 11248
rect 26422 10376 26478 10432
rect 26146 10260 26202 10296
rect 26146 10240 26148 10260
rect 26148 10240 26200 10260
rect 26200 10240 26202 10260
rect 25778 6704 25834 6760
rect 26790 11056 26846 11112
rect 27158 18128 27214 18184
rect 27250 17856 27306 17912
rect 27526 15988 27528 16008
rect 27528 15988 27580 16008
rect 27580 15988 27582 16008
rect 27250 14456 27306 14512
rect 27250 11464 27306 11520
rect 26514 6160 26570 6216
rect 25134 5208 25190 5264
rect 24766 5072 24822 5128
rect 24950 4156 24952 4176
rect 24952 4156 25004 4176
rect 25004 4156 25006 4176
rect 24950 4120 25006 4156
rect 26698 4820 26754 4856
rect 26698 4800 26700 4820
rect 26700 4800 26752 4820
rect 26752 4800 26754 4820
rect 27250 9696 27306 9752
rect 27526 15952 27582 15988
rect 27526 13640 27582 13696
rect 27618 13232 27674 13288
rect 27802 11872 27858 11928
rect 27342 7248 27398 7304
rect 26790 4664 26846 4720
rect 26606 3848 26662 3904
rect 27526 8744 27582 8800
rect 27526 8064 27582 8120
rect 27434 6432 27490 6488
rect 27618 7692 27620 7712
rect 27620 7692 27672 7712
rect 27672 7692 27674 7712
rect 27618 7656 27674 7692
rect 26514 3168 26570 3224
rect 26790 2932 26792 2952
rect 26792 2932 26844 2952
rect 26844 2932 26846 2952
rect 26790 2896 26846 2932
rect 27986 12416 28042 12472
rect 27986 11056 28042 11112
rect 27802 3440 27858 3496
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 36818 38800 36874 38856
rect 28262 15272 28318 15328
rect 28538 15136 28594 15192
rect 28446 14592 28502 14648
rect 28814 15272 28870 15328
rect 28998 15272 29054 15328
rect 28906 15136 28962 15192
rect 29182 15408 29238 15464
rect 28630 14864 28686 14920
rect 28262 14068 28318 14104
rect 28262 14048 28264 14068
rect 28264 14048 28316 14068
rect 28316 14048 28318 14068
rect 28170 11620 28226 11656
rect 28170 11600 28172 11620
rect 28172 11600 28224 11620
rect 28224 11600 28226 11620
rect 28538 12008 28594 12064
rect 28446 10920 28502 10976
rect 28906 14612 28962 14648
rect 28906 14592 28908 14612
rect 28908 14592 28960 14612
rect 28960 14592 28962 14612
rect 28906 14476 28962 14512
rect 28906 14456 28908 14476
rect 28908 14456 28960 14476
rect 28960 14456 28962 14476
rect 29182 14592 29238 14648
rect 28998 13796 29054 13832
rect 28998 13776 29000 13796
rect 29000 13776 29052 13796
rect 29052 13776 29054 13796
rect 29182 13812 29184 13832
rect 29184 13812 29236 13832
rect 29236 13812 29238 13832
rect 29182 13776 29238 13812
rect 29182 13640 29238 13696
rect 28998 12960 29054 13016
rect 28998 12844 29054 12880
rect 28998 12824 29000 12844
rect 29000 12824 29052 12844
rect 29052 12824 29054 12844
rect 28998 12300 29054 12336
rect 28998 12280 29000 12300
rect 29000 12280 29052 12300
rect 29052 12280 29054 12300
rect 29090 12044 29092 12064
rect 29092 12044 29144 12064
rect 29144 12044 29146 12064
rect 29090 12008 29146 12044
rect 29090 11756 29146 11792
rect 29090 11736 29092 11756
rect 29092 11736 29144 11756
rect 29144 11736 29146 11756
rect 28998 11464 29054 11520
rect 29182 11328 29238 11384
rect 29090 11192 29146 11248
rect 28814 6604 28816 6624
rect 28816 6604 28868 6624
rect 28868 6604 28870 6624
rect 28814 6568 28870 6604
rect 29090 6332 29092 6352
rect 29092 6332 29144 6352
rect 29144 6332 29146 6352
rect 29090 6296 29146 6332
rect 29458 15272 29514 15328
rect 29366 14356 29368 14376
rect 29368 14356 29420 14376
rect 29420 14356 29422 14376
rect 29366 14320 29422 14356
rect 29274 7148 29276 7168
rect 29276 7148 29328 7168
rect 29328 7148 29330 7168
rect 29274 7112 29330 7148
rect 29274 6316 29330 6352
rect 29274 6296 29276 6316
rect 29276 6296 29328 6316
rect 29328 6296 29330 6316
rect 29550 13912 29606 13968
rect 30010 15000 30066 15056
rect 29918 13912 29974 13968
rect 29918 13812 29920 13832
rect 29920 13812 29972 13832
rect 29972 13812 29974 13832
rect 29918 13776 29974 13812
rect 29734 11772 29736 11792
rect 29736 11772 29788 11792
rect 29788 11772 29790 11792
rect 29734 11736 29790 11772
rect 29458 5888 29514 5944
rect 29458 4800 29514 4856
rect 29642 5480 29698 5536
rect 29642 3612 29644 3632
rect 29644 3612 29696 3632
rect 29696 3612 29698 3632
rect 29642 3576 29698 3612
rect 29826 6024 29882 6080
rect 30102 11872 30158 11928
rect 30654 12960 30710 13016
rect 29918 5752 29974 5808
rect 29918 5364 29974 5400
rect 29918 5344 29920 5364
rect 29920 5344 29972 5364
rect 29972 5344 29974 5364
rect 30470 12008 30526 12064
rect 30470 11464 30526 11520
rect 30378 8064 30434 8120
rect 30562 11092 30564 11112
rect 30564 11092 30616 11112
rect 30616 11092 30618 11112
rect 30562 11056 30618 11092
rect 30194 2896 30250 2952
rect 30838 9152 30894 9208
rect 31390 14864 31446 14920
rect 31022 9152 31078 9208
rect 31022 6704 31078 6760
rect 31022 6604 31024 6624
rect 31024 6604 31076 6624
rect 31076 6604 31078 6624
rect 31022 6568 31078 6604
rect 31114 6316 31170 6352
rect 31114 6296 31116 6316
rect 31116 6296 31168 6316
rect 31168 6296 31170 6316
rect 31298 5072 31354 5128
rect 32310 14612 32366 14648
rect 32310 14592 32312 14612
rect 32312 14592 32364 14612
rect 32364 14592 32366 14612
rect 31758 13640 31814 13696
rect 31482 6024 31538 6080
rect 31574 5208 31630 5264
rect 30930 3576 30986 3632
rect 31206 3712 31262 3768
rect 31298 2488 31354 2544
rect 31666 3168 31722 3224
rect 31942 5344 31998 5400
rect 32034 4528 32090 4584
rect 32402 12300 32458 12336
rect 32402 12280 32404 12300
rect 32404 12280 32456 12300
rect 32456 12280 32458 12300
rect 32218 4820 32274 4856
rect 32218 4800 32220 4820
rect 32220 4800 32272 4820
rect 32272 4800 32274 4820
rect 32034 3576 32090 3632
rect 32310 3612 32312 3632
rect 32312 3612 32364 3632
rect 32364 3612 32366 3632
rect 32310 3576 32366 3612
rect 32494 7384 32550 7440
rect 32954 12860 32956 12880
rect 32956 12860 33008 12880
rect 33008 12860 33010 12880
rect 32954 12824 33010 12860
rect 32678 9968 32734 10024
rect 32862 7148 32864 7168
rect 32864 7148 32916 7168
rect 32916 7148 32918 7168
rect 32862 7112 32918 7148
rect 32402 3168 32458 3224
rect 33138 4936 33194 4992
rect 38198 37440 38254 37496
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 38290 35400 38346 35456
rect 38198 33380 38254 33416
rect 38198 33360 38200 33380
rect 38200 33360 38252 33380
rect 38252 33360 38254 33380
rect 38290 32020 38346 32056
rect 38290 32000 38292 32020
rect 38292 32000 38344 32020
rect 38344 32000 38346 32020
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 33782 5072 33838 5128
rect 33782 3612 33784 3632
rect 33784 3612 33836 3632
rect 33836 3612 33838 3632
rect 33782 3576 33838 3612
rect 34150 5888 34206 5944
rect 34610 6452 34666 6488
rect 34610 6432 34612 6452
rect 34612 6432 34664 6452
rect 34664 6432 34666 6452
rect 34518 5228 34574 5264
rect 34518 5208 34520 5228
rect 34520 5208 34572 5228
rect 34572 5208 34574 5228
rect 34150 3304 34206 3360
rect 34242 2896 34298 2952
rect 34518 3440 34574 3496
rect 34426 3168 34482 3224
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34978 4428 34980 4448
rect 34980 4428 35032 4448
rect 35032 4428 35034 4448
rect 34978 4392 35034 4428
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34794 3712 34850 3768
rect 34978 3032 35034 3088
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 36542 6704 36598 6760
rect 36174 2488 36230 2544
rect 36266 2352 36322 2408
rect 38198 29960 38254 30016
rect 38198 27920 38254 27976
rect 38290 26580 38346 26616
rect 38290 26560 38292 26580
rect 38292 26560 38344 26580
rect 38344 26560 38346 26580
rect 38290 24520 38346 24576
rect 38198 22500 38254 22536
rect 38198 22480 38200 22500
rect 38200 22480 38252 22500
rect 38252 22480 38254 22500
rect 38198 21120 38254 21176
rect 38198 19116 38200 19136
rect 38200 19116 38252 19136
rect 38252 19116 38254 19136
rect 38198 19080 38254 19116
rect 38290 17076 38292 17096
rect 38292 17076 38344 17096
rect 38344 17076 38346 17096
rect 38290 17040 38346 17076
rect 38198 15680 38254 15736
rect 38290 13640 38346 13696
rect 37186 1400 37242 1456
rect 38198 11600 38254 11656
rect 38014 9016 38070 9072
rect 37922 5480 37978 5536
rect 38290 10260 38346 10296
rect 38290 10240 38292 10260
rect 38292 10240 38344 10260
rect 38344 10240 38346 10260
rect 38290 8200 38346 8256
rect 38198 6160 38254 6216
rect 38106 4800 38162 4856
rect 38198 2760 38254 2816
<< metal3 >>
rect 200 39538 800 39568
rect 2865 39538 2931 39541
rect 200 39536 2931 39538
rect 200 39480 2870 39536
rect 2926 39480 2931 39536
rect 200 39478 2931 39480
rect 200 39448 800 39478
rect 2865 39475 2931 39478
rect 36813 38858 36879 38861
rect 39200 38858 39800 38888
rect 36813 38856 39800 38858
rect 36813 38800 36818 38856
rect 36874 38800 39800 38856
rect 36813 38798 39800 38800
rect 36813 38795 36879 38798
rect 39200 38768 39800 38798
rect 4210 37568 4526 37569
rect 200 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 1669 37498 1735 37501
rect 200 37496 1735 37498
rect 200 37440 1674 37496
rect 1730 37440 1735 37496
rect 200 37438 1735 37440
rect 200 37408 800 37438
rect 1669 37435 1735 37438
rect 38193 37498 38259 37501
rect 39200 37498 39800 37528
rect 38193 37496 39800 37498
rect 38193 37440 38198 37496
rect 38254 37440 39800 37496
rect 38193 37438 39800 37440
rect 38193 37435 38259 37438
rect 39200 37408 39800 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 200 36138 800 36168
rect 1669 36138 1735 36141
rect 200 36136 1735 36138
rect 200 36080 1674 36136
rect 1730 36080 1735 36136
rect 200 36078 1735 36080
rect 200 36048 800 36078
rect 1669 36075 1735 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 38285 35458 38351 35461
rect 39200 35458 39800 35488
rect 38285 35456 39800 35458
rect 38285 35400 38290 35456
rect 38346 35400 39800 35456
rect 38285 35398 39800 35400
rect 38285 35395 38351 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 39200 35368 39800 35398
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 200 34098 800 34128
rect 1669 34098 1735 34101
rect 200 34096 1735 34098
rect 200 34040 1674 34096
rect 1730 34040 1735 34096
rect 200 34038 1735 34040
rect 200 34008 800 34038
rect 1669 34035 1735 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 38193 33418 38259 33421
rect 39200 33418 39800 33448
rect 38193 33416 39800 33418
rect 38193 33360 38198 33416
rect 38254 33360 39800 33416
rect 38193 33358 39800 33360
rect 38193 33355 38259 33358
rect 39200 33328 39800 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 200 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1669 32058 1735 32061
rect 200 32056 1735 32058
rect 200 32000 1674 32056
rect 1730 32000 1735 32056
rect 200 31998 1735 32000
rect 200 31968 800 31998
rect 1669 31995 1735 31998
rect 38285 32058 38351 32061
rect 39200 32058 39800 32088
rect 38285 32056 39800 32058
rect 38285 32000 38290 32056
rect 38346 32000 39800 32056
rect 38285 31998 39800 32000
rect 38285 31995 38351 31998
rect 39200 31968 39800 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30698 800 30728
rect 1669 30698 1735 30701
rect 200 30696 1735 30698
rect 200 30640 1674 30696
rect 1730 30640 1735 30696
rect 200 30638 1735 30640
rect 200 30608 800 30638
rect 1669 30635 1735 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 38193 30018 38259 30021
rect 39200 30018 39800 30048
rect 38193 30016 39800 30018
rect 38193 29960 38198 30016
rect 38254 29960 39800 30016
rect 38193 29958 39800 29960
rect 38193 29955 38259 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 39200 29928 39800 29958
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 200 28658 800 28688
rect 1577 28658 1643 28661
rect 200 28656 1643 28658
rect 200 28600 1582 28656
rect 1638 28600 1643 28656
rect 200 28598 1643 28600
rect 200 28568 800 28598
rect 1577 28595 1643 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 38193 27978 38259 27981
rect 39200 27978 39800 28008
rect 38193 27976 39800 27978
rect 38193 27920 38198 27976
rect 38254 27920 39800 27976
rect 38193 27918 39800 27920
rect 38193 27915 38259 27918
rect 39200 27888 39800 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 200 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 1669 26618 1735 26621
rect 200 26616 1735 26618
rect 200 26560 1674 26616
rect 1730 26560 1735 26616
rect 200 26558 1735 26560
rect 200 26528 800 26558
rect 1669 26555 1735 26558
rect 38285 26618 38351 26621
rect 39200 26618 39800 26648
rect 38285 26616 39800 26618
rect 38285 26560 38290 26616
rect 38346 26560 39800 26616
rect 38285 26558 39800 26560
rect 38285 26555 38351 26558
rect 39200 26528 39800 26558
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 200 25258 800 25288
rect 1577 25258 1643 25261
rect 200 25256 1643 25258
rect 200 25200 1582 25256
rect 1638 25200 1643 25256
rect 200 25198 1643 25200
rect 200 25168 800 25198
rect 1577 25195 1643 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 38285 24578 38351 24581
rect 39200 24578 39800 24608
rect 38285 24576 39800 24578
rect 38285 24520 38290 24576
rect 38346 24520 39800 24576
rect 38285 24518 39800 24520
rect 38285 24515 38351 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 39200 24488 39800 24518
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 200 23218 800 23248
rect 1577 23218 1643 23221
rect 200 23216 1643 23218
rect 200 23160 1582 23216
rect 1638 23160 1643 23216
rect 200 23158 1643 23160
rect 200 23128 800 23158
rect 1577 23155 1643 23158
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 38193 22538 38259 22541
rect 39200 22538 39800 22568
rect 38193 22536 39800 22538
rect 38193 22480 38198 22536
rect 38254 22480 39800 22536
rect 38193 22478 39800 22480
rect 38193 22475 38259 22478
rect 39200 22448 39800 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 200 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 1669 21178 1735 21181
rect 200 21176 1735 21178
rect 200 21120 1674 21176
rect 1730 21120 1735 21176
rect 200 21118 1735 21120
rect 200 21088 800 21118
rect 1669 21115 1735 21118
rect 38193 21178 38259 21181
rect 39200 21178 39800 21208
rect 38193 21176 39800 21178
rect 38193 21120 38198 21176
rect 38254 21120 39800 21176
rect 38193 21118 39800 21120
rect 38193 21115 38259 21118
rect 39200 21088 39800 21118
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 200 19818 800 19848
rect 1669 19818 1735 19821
rect 200 19816 1735 19818
rect 200 19760 1674 19816
rect 1730 19760 1735 19816
rect 200 19758 1735 19760
rect 200 19728 800 19758
rect 1669 19755 1735 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 38193 19138 38259 19141
rect 39200 19138 39800 19168
rect 38193 19136 39800 19138
rect 38193 19080 38198 19136
rect 38254 19080 39800 19136
rect 38193 19078 39800 19080
rect 38193 19075 38259 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 39800 19078
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 19885 18186 19951 18189
rect 27153 18186 27219 18189
rect 19885 18184 27219 18186
rect 19885 18128 19890 18184
rect 19946 18128 27158 18184
rect 27214 18128 27219 18184
rect 19885 18126 27219 18128
rect 19885 18123 19951 18126
rect 27153 18123 27219 18126
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 20437 17914 20503 17917
rect 22093 17914 22159 17917
rect 27245 17914 27311 17917
rect 20437 17912 27311 17914
rect 20437 17856 20442 17912
rect 20498 17856 22098 17912
rect 22154 17856 27250 17912
rect 27306 17856 27311 17912
rect 20437 17854 27311 17856
rect 20437 17851 20503 17854
rect 22093 17851 22159 17854
rect 27245 17851 27311 17854
rect 200 17778 800 17808
rect 1669 17778 1735 17781
rect 200 17776 1735 17778
rect 200 17720 1674 17776
rect 1730 17720 1735 17776
rect 200 17718 1735 17720
rect 200 17688 800 17718
rect 1669 17715 1735 17718
rect 23238 17580 23244 17644
rect 23308 17642 23314 17644
rect 26049 17642 26115 17645
rect 23308 17640 26115 17642
rect 23308 17584 26054 17640
rect 26110 17584 26115 17640
rect 23308 17582 26115 17584
rect 23308 17580 23314 17582
rect 26049 17579 26115 17582
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 23565 17370 23631 17373
rect 26509 17370 26575 17373
rect 23565 17368 26575 17370
rect 23565 17312 23570 17368
rect 23626 17312 26514 17368
rect 26570 17312 26575 17368
rect 23565 17310 26575 17312
rect 23565 17307 23631 17310
rect 26509 17307 26575 17310
rect 38285 17098 38351 17101
rect 39200 17098 39800 17128
rect 38285 17096 39800 17098
rect 38285 17040 38290 17096
rect 38346 17040 39800 17096
rect 38285 17038 39800 17040
rect 38285 17035 38351 17038
rect 39200 17008 39800 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 21449 16554 21515 16557
rect 25773 16554 25839 16557
rect 21449 16552 25839 16554
rect 21449 16496 21454 16552
rect 21510 16496 25778 16552
rect 25834 16496 25839 16552
rect 21449 16494 25839 16496
rect 21449 16491 21515 16494
rect 25773 16491 25839 16494
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 20529 16010 20595 16013
rect 27521 16010 27587 16013
rect 20529 16008 27587 16010
rect 20529 15952 20534 16008
rect 20590 15952 27526 16008
rect 27582 15952 27587 16008
rect 20529 15950 27587 15952
rect 20529 15947 20595 15950
rect 27521 15947 27587 15950
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1669 15738 1735 15741
rect 200 15736 1735 15738
rect 200 15680 1674 15736
rect 1730 15680 1735 15736
rect 200 15678 1735 15680
rect 200 15648 800 15678
rect 1669 15675 1735 15678
rect 38193 15738 38259 15741
rect 39200 15738 39800 15768
rect 38193 15736 39800 15738
rect 38193 15680 38198 15736
rect 38254 15680 39800 15736
rect 38193 15678 39800 15680
rect 38193 15675 38259 15678
rect 39200 15648 39800 15678
rect 16205 15466 16271 15469
rect 29177 15466 29243 15469
rect 16205 15464 29243 15466
rect 16205 15408 16210 15464
rect 16266 15408 29182 15464
rect 29238 15408 29243 15464
rect 16205 15406 29243 15408
rect 16205 15403 16271 15406
rect 29177 15403 29243 15406
rect 21265 15330 21331 15333
rect 21398 15330 21404 15332
rect 21265 15328 21404 15330
rect 21265 15272 21270 15328
rect 21326 15272 21404 15328
rect 21265 15270 21404 15272
rect 21265 15267 21331 15270
rect 21398 15268 21404 15270
rect 21468 15268 21474 15332
rect 28257 15330 28323 15333
rect 28809 15330 28875 15333
rect 28257 15328 28875 15330
rect 28257 15272 28262 15328
rect 28318 15272 28814 15328
rect 28870 15272 28875 15328
rect 28257 15270 28875 15272
rect 28257 15267 28323 15270
rect 28809 15267 28875 15270
rect 28993 15330 29059 15333
rect 29453 15330 29519 15333
rect 28993 15328 29519 15330
rect 28993 15272 28998 15328
rect 29054 15272 29458 15328
rect 29514 15272 29519 15328
rect 28993 15270 29519 15272
rect 28993 15267 29059 15270
rect 29453 15267 29519 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 28533 15194 28599 15197
rect 28901 15194 28967 15197
rect 28533 15192 28967 15194
rect 28533 15136 28538 15192
rect 28594 15136 28906 15192
rect 28962 15136 28967 15192
rect 28533 15134 28967 15136
rect 28533 15131 28599 15134
rect 28901 15131 28967 15134
rect 26693 15058 26759 15061
rect 30005 15058 30071 15061
rect 26693 15056 30071 15058
rect 26693 15000 26698 15056
rect 26754 15000 30010 15056
rect 30066 15000 30071 15056
rect 26693 14998 30071 15000
rect 26693 14995 26759 14998
rect 30005 14995 30071 14998
rect 28625 14922 28691 14925
rect 31385 14922 31451 14925
rect 28625 14920 31451 14922
rect 28625 14864 28630 14920
rect 28686 14864 31390 14920
rect 31446 14864 31451 14920
rect 28625 14862 31451 14864
rect 28625 14859 28691 14862
rect 31385 14859 31451 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 28441 14650 28507 14653
rect 28901 14650 28967 14653
rect 28441 14648 28967 14650
rect 28441 14592 28446 14648
rect 28502 14592 28906 14648
rect 28962 14592 28967 14648
rect 28441 14590 28967 14592
rect 28441 14587 28507 14590
rect 28901 14587 28967 14590
rect 29177 14650 29243 14653
rect 32305 14650 32371 14653
rect 29177 14648 32371 14650
rect 29177 14592 29182 14648
rect 29238 14592 32310 14648
rect 32366 14592 32371 14648
rect 29177 14590 32371 14592
rect 29177 14587 29243 14590
rect 32305 14587 32371 14590
rect 20621 14514 20687 14517
rect 22277 14514 22343 14517
rect 20621 14512 22343 14514
rect 20621 14456 20626 14512
rect 20682 14456 22282 14512
rect 22338 14456 22343 14512
rect 20621 14454 22343 14456
rect 20621 14451 20687 14454
rect 22277 14451 22343 14454
rect 27245 14514 27311 14517
rect 28901 14514 28967 14517
rect 27245 14512 28967 14514
rect 27245 14456 27250 14512
rect 27306 14456 28906 14512
rect 28962 14456 28967 14512
rect 27245 14454 28967 14456
rect 27245 14451 27311 14454
rect 28901 14451 28967 14454
rect 200 14378 800 14408
rect 1577 14378 1643 14381
rect 200 14376 1643 14378
rect 200 14320 1582 14376
rect 1638 14320 1643 14376
rect 200 14318 1643 14320
rect 200 14288 800 14318
rect 1577 14315 1643 14318
rect 22001 14378 22067 14381
rect 25129 14378 25195 14381
rect 25497 14378 25563 14381
rect 29361 14378 29427 14381
rect 22001 14376 29427 14378
rect 22001 14320 22006 14376
rect 22062 14320 25134 14376
rect 25190 14320 25502 14376
rect 25558 14320 29366 14376
rect 29422 14320 29427 14376
rect 22001 14318 29427 14320
rect 22001 14315 22067 14318
rect 25129 14315 25195 14318
rect 25497 14315 25563 14318
rect 29361 14315 29427 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 19977 14106 20043 14109
rect 21633 14106 21699 14109
rect 19977 14104 21699 14106
rect 19977 14048 19982 14104
rect 20038 14048 21638 14104
rect 21694 14048 21699 14104
rect 19977 14046 21699 14048
rect 19977 14043 20043 14046
rect 21633 14043 21699 14046
rect 24117 14106 24183 14109
rect 28257 14106 28323 14109
rect 24117 14104 28323 14106
rect 24117 14048 24122 14104
rect 24178 14048 28262 14104
rect 28318 14048 28323 14104
rect 24117 14046 28323 14048
rect 24117 14043 24183 14046
rect 28257 14043 28323 14046
rect 23289 13970 23355 13973
rect 29545 13970 29611 13973
rect 29913 13970 29979 13973
rect 23289 13968 29979 13970
rect 23289 13912 23294 13968
rect 23350 13912 29550 13968
rect 29606 13912 29918 13968
rect 29974 13912 29979 13968
rect 23289 13910 29979 13912
rect 23289 13907 23355 13910
rect 29545 13907 29611 13910
rect 29913 13907 29979 13910
rect 22277 13834 22343 13837
rect 28993 13834 29059 13837
rect 22277 13832 29059 13834
rect 22277 13776 22282 13832
rect 22338 13776 28998 13832
rect 29054 13776 29059 13832
rect 22277 13774 29059 13776
rect 22277 13771 22343 13774
rect 28993 13771 29059 13774
rect 29177 13834 29243 13837
rect 29913 13834 29979 13837
rect 29177 13832 29979 13834
rect 29177 13776 29182 13832
rect 29238 13776 29918 13832
rect 29974 13776 29979 13832
rect 29177 13774 29979 13776
rect 29177 13771 29243 13774
rect 29913 13771 29979 13774
rect 27521 13698 27587 13701
rect 29177 13698 29243 13701
rect 31753 13698 31819 13701
rect 27521 13696 31819 13698
rect 27521 13640 27526 13696
rect 27582 13640 29182 13696
rect 29238 13640 31758 13696
rect 31814 13640 31819 13696
rect 27521 13638 31819 13640
rect 27521 13635 27587 13638
rect 29177 13635 29243 13638
rect 31753 13635 31819 13638
rect 38285 13698 38351 13701
rect 39200 13698 39800 13728
rect 38285 13696 39800 13698
rect 38285 13640 38290 13696
rect 38346 13640 39800 13696
rect 38285 13638 39800 13640
rect 38285 13635 38351 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 39200 13608 39800 13638
rect 34930 13567 35246 13568
rect 14733 13426 14799 13429
rect 24025 13426 24091 13429
rect 14733 13424 24091 13426
rect 14733 13368 14738 13424
rect 14794 13368 24030 13424
rect 24086 13368 24091 13424
rect 14733 13366 24091 13368
rect 14733 13363 14799 13366
rect 24025 13363 24091 13366
rect 17217 13290 17283 13293
rect 19057 13290 19123 13293
rect 17217 13288 19123 13290
rect 17217 13232 17222 13288
rect 17278 13232 19062 13288
rect 19118 13232 19123 13288
rect 17217 13230 19123 13232
rect 17217 13227 17283 13230
rect 19057 13227 19123 13230
rect 25681 13290 25747 13293
rect 27613 13290 27679 13293
rect 25681 13288 27679 13290
rect 25681 13232 25686 13288
rect 25742 13232 27618 13288
rect 27674 13232 27679 13288
rect 25681 13230 27679 13232
rect 25681 13227 25747 13230
rect 27613 13227 27679 13230
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 28993 13018 29059 13021
rect 30649 13018 30715 13021
rect 28993 13016 30715 13018
rect 28993 12960 28998 13016
rect 29054 12960 30654 13016
rect 30710 12960 30715 13016
rect 28993 12958 30715 12960
rect 28993 12955 29059 12958
rect 30649 12955 30715 12958
rect 17217 12882 17283 12885
rect 17350 12882 17356 12884
rect 17217 12880 17356 12882
rect 17217 12824 17222 12880
rect 17278 12824 17356 12880
rect 17217 12822 17356 12824
rect 17217 12819 17283 12822
rect 17350 12820 17356 12822
rect 17420 12820 17426 12884
rect 28993 12882 29059 12885
rect 32949 12882 33015 12885
rect 28993 12880 33015 12882
rect 28993 12824 28998 12880
rect 29054 12824 32954 12880
rect 33010 12824 33015 12880
rect 28993 12822 33015 12824
rect 28993 12819 29059 12822
rect 32949 12819 33015 12822
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 20621 12474 20687 12477
rect 27981 12474 28047 12477
rect 20621 12472 28047 12474
rect 20621 12416 20626 12472
rect 20682 12416 27986 12472
rect 28042 12416 28047 12472
rect 20621 12414 28047 12416
rect 20621 12411 20687 12414
rect 27981 12411 28047 12414
rect 200 12338 800 12368
rect 1669 12338 1735 12341
rect 200 12336 1735 12338
rect 200 12280 1674 12336
rect 1730 12280 1735 12336
rect 200 12278 1735 12280
rect 200 12248 800 12278
rect 1669 12275 1735 12278
rect 28993 12338 29059 12341
rect 32397 12338 32463 12341
rect 28993 12336 32463 12338
rect 28993 12280 28998 12336
rect 29054 12280 32402 12336
rect 32458 12280 32463 12336
rect 28993 12278 32463 12280
rect 28993 12275 29059 12278
rect 32397 12275 32463 12278
rect 15837 12202 15903 12205
rect 16665 12202 16731 12205
rect 15837 12200 16731 12202
rect 15837 12144 15842 12200
rect 15898 12144 16670 12200
rect 16726 12144 16731 12200
rect 15837 12142 16731 12144
rect 15837 12139 15903 12142
rect 16665 12139 16731 12142
rect 16849 12202 16915 12205
rect 21081 12202 21147 12205
rect 16849 12200 21147 12202
rect 16849 12144 16854 12200
rect 16910 12144 21086 12200
rect 21142 12144 21147 12200
rect 16849 12142 21147 12144
rect 16849 12139 16915 12142
rect 21081 12139 21147 12142
rect 25129 12066 25195 12069
rect 28533 12066 28599 12069
rect 25129 12064 28599 12066
rect 25129 12008 25134 12064
rect 25190 12008 28538 12064
rect 28594 12008 28599 12064
rect 25129 12006 28599 12008
rect 25129 12003 25195 12006
rect 28533 12003 28599 12006
rect 29085 12066 29151 12069
rect 30465 12066 30531 12069
rect 29085 12064 30531 12066
rect 29085 12008 29090 12064
rect 29146 12008 30470 12064
rect 30526 12008 30531 12064
rect 29085 12006 30531 12008
rect 29085 12003 29151 12006
rect 30465 12003 30531 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 16297 11930 16363 11933
rect 27797 11930 27863 11933
rect 30097 11930 30163 11933
rect 16297 11928 19350 11930
rect 16297 11872 16302 11928
rect 16358 11872 19350 11928
rect 16297 11870 19350 11872
rect 16297 11867 16363 11870
rect 19290 11794 19350 11870
rect 27797 11928 30163 11930
rect 27797 11872 27802 11928
rect 27858 11872 30102 11928
rect 30158 11872 30163 11928
rect 27797 11870 30163 11872
rect 27797 11867 27863 11870
rect 30097 11867 30163 11870
rect 19793 11794 19859 11797
rect 19290 11792 19859 11794
rect 19290 11736 19798 11792
rect 19854 11736 19859 11792
rect 19290 11734 19859 11736
rect 19793 11731 19859 11734
rect 29085 11794 29151 11797
rect 29729 11794 29795 11797
rect 29085 11792 29795 11794
rect 29085 11736 29090 11792
rect 29146 11736 29734 11792
rect 29790 11736 29795 11792
rect 29085 11734 29795 11736
rect 29085 11731 29151 11734
rect 29729 11731 29795 11734
rect 23749 11658 23815 11661
rect 28165 11658 28231 11661
rect 23749 11656 28231 11658
rect 23749 11600 23754 11656
rect 23810 11600 28170 11656
rect 28226 11600 28231 11656
rect 23749 11598 28231 11600
rect 23749 11595 23815 11598
rect 28165 11595 28231 11598
rect 38193 11658 38259 11661
rect 39200 11658 39800 11688
rect 38193 11656 39800 11658
rect 38193 11600 38198 11656
rect 38254 11600 39800 11656
rect 38193 11598 39800 11600
rect 38193 11595 38259 11598
rect 39200 11568 39800 11598
rect 20989 11522 21055 11525
rect 27245 11522 27311 11525
rect 20989 11520 27311 11522
rect 20989 11464 20994 11520
rect 21050 11464 27250 11520
rect 27306 11464 27311 11520
rect 20989 11462 27311 11464
rect 20989 11459 21055 11462
rect 27245 11459 27311 11462
rect 28993 11522 29059 11525
rect 30465 11522 30531 11525
rect 28993 11520 30531 11522
rect 28993 11464 28998 11520
rect 29054 11464 30470 11520
rect 30526 11464 30531 11520
rect 28993 11462 30531 11464
rect 28993 11459 29059 11462
rect 30465 11459 30531 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 25129 11386 25195 11389
rect 29177 11386 29243 11389
rect 25129 11384 29243 11386
rect 25129 11328 25134 11384
rect 25190 11328 29182 11384
rect 29238 11328 29243 11384
rect 25129 11326 29243 11328
rect 25129 11323 25195 11326
rect 29177 11323 29243 11326
rect 19241 11250 19307 11253
rect 20989 11250 21055 11253
rect 19241 11248 21055 11250
rect 19241 11192 19246 11248
rect 19302 11192 20994 11248
rect 21050 11192 21055 11248
rect 19241 11190 21055 11192
rect 19241 11187 19307 11190
rect 20989 11187 21055 11190
rect 22829 11250 22895 11253
rect 25405 11250 25471 11253
rect 22829 11248 25471 11250
rect 22829 11192 22834 11248
rect 22890 11192 25410 11248
rect 25466 11192 25471 11248
rect 22829 11190 25471 11192
rect 22829 11187 22895 11190
rect 25405 11187 25471 11190
rect 26509 11250 26575 11253
rect 29085 11250 29151 11253
rect 26509 11248 29151 11250
rect 26509 11192 26514 11248
rect 26570 11192 29090 11248
rect 29146 11192 29151 11248
rect 26509 11190 29151 11192
rect 26509 11187 26575 11190
rect 29085 11187 29151 11190
rect 19793 11114 19859 11117
rect 23473 11114 23539 11117
rect 19793 11112 23539 11114
rect 19793 11056 19798 11112
rect 19854 11056 23478 11112
rect 23534 11056 23539 11112
rect 19793 11054 23539 11056
rect 19793 11051 19859 11054
rect 23473 11051 23539 11054
rect 24209 11114 24275 11117
rect 26785 11114 26851 11117
rect 24209 11112 26851 11114
rect 24209 11056 24214 11112
rect 24270 11056 26790 11112
rect 26846 11056 26851 11112
rect 24209 11054 26851 11056
rect 24209 11051 24275 11054
rect 26785 11051 26851 11054
rect 27981 11114 28047 11117
rect 30557 11114 30623 11117
rect 27981 11112 30623 11114
rect 27981 11056 27986 11112
rect 28042 11056 30562 11112
rect 30618 11056 30623 11112
rect 27981 11054 30623 11056
rect 27981 11051 28047 11054
rect 30557 11051 30623 11054
rect 22093 10978 22159 10981
rect 24577 10978 24643 10981
rect 28441 10978 28507 10981
rect 22093 10976 28507 10978
rect 22093 10920 22098 10976
rect 22154 10920 24582 10976
rect 24638 10920 28446 10976
rect 28502 10920 28507 10976
rect 22093 10918 28507 10920
rect 22093 10915 22159 10918
rect 24577 10915 24643 10918
rect 28441 10915 28507 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 21541 10706 21607 10709
rect 22185 10706 22251 10709
rect 21541 10704 22251 10706
rect 21541 10648 21546 10704
rect 21602 10648 22190 10704
rect 22246 10648 22251 10704
rect 21541 10646 22251 10648
rect 21541 10643 21607 10646
rect 22185 10643 22251 10646
rect 14825 10570 14891 10573
rect 22829 10570 22895 10573
rect 14825 10568 22895 10570
rect 14825 10512 14830 10568
rect 14886 10512 22834 10568
rect 22890 10512 22895 10568
rect 14825 10510 22895 10512
rect 14825 10507 14891 10510
rect 22829 10507 22895 10510
rect 20345 10434 20411 10437
rect 26417 10434 26483 10437
rect 20345 10432 26483 10434
rect 20345 10376 20350 10432
rect 20406 10376 26422 10432
rect 26478 10376 26483 10432
rect 20345 10374 26483 10376
rect 20345 10371 20411 10374
rect 26417 10371 26483 10374
rect 4210 10368 4526 10369
rect 200 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 1669 10298 1735 10301
rect 200 10296 1735 10298
rect 200 10240 1674 10296
rect 1730 10240 1735 10296
rect 200 10238 1735 10240
rect 200 10208 800 10238
rect 1669 10235 1735 10238
rect 19425 10298 19491 10301
rect 21909 10298 21975 10301
rect 26141 10298 26207 10301
rect 19425 10296 26207 10298
rect 19425 10240 19430 10296
rect 19486 10240 21914 10296
rect 21970 10240 26146 10296
rect 26202 10240 26207 10296
rect 19425 10238 26207 10240
rect 19425 10235 19491 10238
rect 21909 10235 21975 10238
rect 26141 10235 26207 10238
rect 38285 10298 38351 10301
rect 39200 10298 39800 10328
rect 38285 10296 39800 10298
rect 38285 10240 38290 10296
rect 38346 10240 39800 10296
rect 38285 10238 39800 10240
rect 38285 10235 38351 10238
rect 39200 10208 39800 10238
rect 15653 10162 15719 10165
rect 16849 10162 16915 10165
rect 20621 10162 20687 10165
rect 15653 10160 20687 10162
rect 15653 10104 15658 10160
rect 15714 10104 16854 10160
rect 16910 10104 20626 10160
rect 20682 10104 20687 10160
rect 15653 10102 20687 10104
rect 15653 10099 15719 10102
rect 16849 10099 16915 10102
rect 20621 10099 20687 10102
rect 21909 10026 21975 10029
rect 32673 10026 32739 10029
rect 21909 10024 32739 10026
rect 21909 9968 21914 10024
rect 21970 9968 32678 10024
rect 32734 9968 32739 10024
rect 21909 9966 32739 9968
rect 21909 9963 21975 9966
rect 32673 9963 32739 9966
rect 17769 9890 17835 9893
rect 18413 9890 18479 9893
rect 17769 9888 18479 9890
rect 17769 9832 17774 9888
rect 17830 9832 18418 9888
rect 18474 9832 18479 9888
rect 17769 9830 18479 9832
rect 17769 9827 17835 9830
rect 18413 9827 18479 9830
rect 20529 9890 20595 9893
rect 22921 9890 22987 9893
rect 20529 9888 22987 9890
rect 20529 9832 20534 9888
rect 20590 9832 22926 9888
rect 22982 9832 22987 9888
rect 20529 9830 22987 9832
rect 20529 9827 20595 9830
rect 22921 9827 22987 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 15653 9754 15719 9757
rect 18229 9754 18295 9757
rect 18597 9754 18663 9757
rect 15653 9752 18663 9754
rect 15653 9696 15658 9752
rect 15714 9696 18234 9752
rect 18290 9696 18602 9752
rect 18658 9696 18663 9752
rect 15653 9694 18663 9696
rect 15653 9691 15719 9694
rect 18229 9691 18295 9694
rect 18597 9691 18663 9694
rect 21817 9754 21883 9757
rect 22737 9754 22803 9757
rect 21817 9752 22803 9754
rect 21817 9696 21822 9752
rect 21878 9696 22742 9752
rect 22798 9696 22803 9752
rect 21817 9694 22803 9696
rect 21817 9691 21883 9694
rect 22737 9691 22803 9694
rect 24485 9754 24551 9757
rect 27245 9754 27311 9757
rect 24485 9752 27311 9754
rect 24485 9696 24490 9752
rect 24546 9696 27250 9752
rect 27306 9696 27311 9752
rect 24485 9694 27311 9696
rect 24485 9691 24551 9694
rect 27245 9691 27311 9694
rect 19977 9618 20043 9621
rect 22553 9618 22619 9621
rect 19977 9616 22619 9618
rect 19977 9560 19982 9616
rect 20038 9560 22558 9616
rect 22614 9560 22619 9616
rect 19977 9558 22619 9560
rect 19977 9555 20043 9558
rect 22553 9555 22619 9558
rect 15285 9482 15351 9485
rect 16297 9482 16363 9485
rect 23565 9482 23631 9485
rect 15285 9480 23631 9482
rect 15285 9424 15290 9480
rect 15346 9424 16302 9480
rect 16358 9424 23570 9480
rect 23626 9424 23631 9480
rect 15285 9422 23631 9424
rect 15285 9419 15351 9422
rect 16297 9419 16363 9422
rect 23565 9419 23631 9422
rect 16665 9346 16731 9349
rect 21909 9346 21975 9349
rect 16665 9344 21975 9346
rect 16665 9288 16670 9344
rect 16726 9288 21914 9344
rect 21970 9288 21975 9344
rect 16665 9286 21975 9288
rect 16665 9283 16731 9286
rect 21909 9283 21975 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 22093 9210 22159 9213
rect 30833 9210 30899 9213
rect 31017 9210 31083 9213
rect 22093 9208 31083 9210
rect 22093 9152 22098 9208
rect 22154 9152 30838 9208
rect 30894 9152 31022 9208
rect 31078 9152 31083 9208
rect 22093 9150 31083 9152
rect 22093 9147 22159 9150
rect 30833 9147 30899 9150
rect 31017 9147 31083 9150
rect 14273 9074 14339 9077
rect 38009 9074 38075 9077
rect 14273 9072 38075 9074
rect 14273 9016 14278 9072
rect 14334 9016 38014 9072
rect 38070 9016 38075 9072
rect 14273 9014 38075 9016
rect 14273 9011 14339 9014
rect 38009 9011 38075 9014
rect 200 8938 800 8968
rect 1669 8938 1735 8941
rect 200 8936 1735 8938
rect 200 8880 1674 8936
rect 1730 8880 1735 8936
rect 200 8878 1735 8880
rect 200 8848 800 8878
rect 1669 8875 1735 8878
rect 20161 8938 20227 8941
rect 24301 8938 24367 8941
rect 20161 8936 24367 8938
rect 20161 8880 20166 8936
rect 20222 8880 24306 8936
rect 24362 8880 24367 8936
rect 20161 8878 24367 8880
rect 20161 8875 20227 8878
rect 24301 8875 24367 8878
rect 23105 8802 23171 8805
rect 27521 8802 27587 8805
rect 23105 8800 27587 8802
rect 23105 8744 23110 8800
rect 23166 8744 27526 8800
rect 27582 8744 27587 8800
rect 23105 8742 27587 8744
rect 23105 8739 23171 8742
rect 27521 8739 27587 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 22093 8666 22159 8669
rect 23749 8666 23815 8669
rect 22093 8664 23815 8666
rect 22093 8608 22098 8664
rect 22154 8608 23754 8664
rect 23810 8608 23815 8664
rect 22093 8606 23815 8608
rect 22093 8603 22159 8606
rect 23749 8603 23815 8606
rect 20713 8530 20779 8533
rect 21265 8530 21331 8533
rect 22001 8530 22067 8533
rect 25221 8530 25287 8533
rect 20713 8528 25287 8530
rect 20713 8472 20718 8528
rect 20774 8472 21270 8528
rect 21326 8472 22006 8528
rect 22062 8472 25226 8528
rect 25282 8472 25287 8528
rect 20713 8470 25287 8472
rect 20713 8467 20779 8470
rect 21265 8467 21331 8470
rect 22001 8467 22067 8470
rect 25221 8467 25287 8470
rect 17953 8394 18019 8397
rect 18965 8394 19031 8397
rect 21817 8394 21883 8397
rect 17953 8392 21883 8394
rect 17953 8336 17958 8392
rect 18014 8336 18970 8392
rect 19026 8336 21822 8392
rect 21878 8336 21883 8392
rect 17953 8334 21883 8336
rect 17953 8331 18019 8334
rect 18965 8331 19031 8334
rect 21817 8331 21883 8334
rect 16389 8258 16455 8261
rect 21357 8258 21423 8261
rect 16389 8256 21423 8258
rect 16389 8200 16394 8256
rect 16450 8200 21362 8256
rect 21418 8200 21423 8256
rect 16389 8198 21423 8200
rect 16389 8195 16455 8198
rect 21357 8195 21423 8198
rect 38285 8258 38351 8261
rect 39200 8258 39800 8288
rect 38285 8256 39800 8258
rect 38285 8200 38290 8256
rect 38346 8200 39800 8256
rect 38285 8198 39800 8200
rect 38285 8195 38351 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 39200 8168 39800 8198
rect 34930 8127 35246 8128
rect 21173 8122 21239 8125
rect 22921 8122 22987 8125
rect 21173 8120 22987 8122
rect 21173 8064 21178 8120
rect 21234 8064 22926 8120
rect 22982 8064 22987 8120
rect 21173 8062 22987 8064
rect 21173 8059 21239 8062
rect 22921 8059 22987 8062
rect 23381 8122 23447 8125
rect 27521 8122 27587 8125
rect 30373 8122 30439 8125
rect 23381 8120 30439 8122
rect 23381 8064 23386 8120
rect 23442 8064 27526 8120
rect 27582 8064 30378 8120
rect 30434 8064 30439 8120
rect 23381 8062 30439 8064
rect 23381 8059 23447 8062
rect 27521 8059 27587 8062
rect 30373 8059 30439 8062
rect 16614 7788 16620 7852
rect 16684 7850 16690 7852
rect 24853 7850 24919 7853
rect 16684 7848 24919 7850
rect 16684 7792 24858 7848
rect 24914 7792 24919 7848
rect 16684 7790 24919 7792
rect 16684 7788 16690 7790
rect 24853 7787 24919 7790
rect 20253 7714 20319 7717
rect 20897 7714 20963 7717
rect 20253 7712 20963 7714
rect 20253 7656 20258 7712
rect 20314 7656 20902 7712
rect 20958 7656 20963 7712
rect 20253 7654 20963 7656
rect 20253 7651 20319 7654
rect 20897 7651 20963 7654
rect 24761 7714 24827 7717
rect 27613 7714 27679 7717
rect 24761 7712 27679 7714
rect 24761 7656 24766 7712
rect 24822 7656 27618 7712
rect 27674 7656 27679 7712
rect 24761 7654 27679 7656
rect 24761 7651 24827 7654
rect 27613 7651 27679 7654
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 7833 7442 7899 7445
rect 19057 7442 19123 7445
rect 32489 7442 32555 7445
rect 7833 7440 32555 7442
rect 7833 7384 7838 7440
rect 7894 7384 19062 7440
rect 19118 7384 32494 7440
rect 32550 7384 32555 7440
rect 7833 7382 32555 7384
rect 7833 7379 7899 7382
rect 19057 7379 19123 7382
rect 32489 7379 32555 7382
rect 24117 7306 24183 7309
rect 27337 7306 27403 7309
rect 24117 7304 27403 7306
rect 24117 7248 24122 7304
rect 24178 7248 27342 7304
rect 27398 7248 27403 7304
rect 24117 7246 27403 7248
rect 24117 7243 24183 7246
rect 27337 7243 27403 7246
rect 21725 7170 21791 7173
rect 22093 7170 22159 7173
rect 21725 7168 22159 7170
rect 21725 7112 21730 7168
rect 21786 7112 22098 7168
rect 22154 7112 22159 7168
rect 21725 7110 22159 7112
rect 21725 7107 21791 7110
rect 22093 7107 22159 7110
rect 29269 7170 29335 7173
rect 32857 7170 32923 7173
rect 29269 7168 32923 7170
rect 29269 7112 29274 7168
rect 29330 7112 32862 7168
rect 32918 7112 32923 7168
rect 29269 7110 32923 7112
rect 29269 7107 29335 7110
rect 32857 7107 32923 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 21909 7034 21975 7037
rect 22369 7034 22435 7037
rect 21909 7032 22435 7034
rect 21909 6976 21914 7032
rect 21970 6976 22374 7032
rect 22430 6976 22435 7032
rect 21909 6974 22435 6976
rect 21909 6971 21975 6974
rect 22369 6971 22435 6974
rect 200 6898 800 6928
rect 1669 6898 1735 6901
rect 200 6896 1735 6898
rect 200 6840 1674 6896
rect 1730 6840 1735 6896
rect 200 6838 1735 6840
rect 200 6808 800 6838
rect 1669 6835 1735 6838
rect 18137 6898 18203 6901
rect 20345 6898 20411 6901
rect 18137 6896 20411 6898
rect 18137 6840 18142 6896
rect 18198 6840 20350 6896
rect 20406 6840 20411 6896
rect 18137 6838 20411 6840
rect 18137 6835 18203 6838
rect 20345 6835 20411 6838
rect 17769 6762 17835 6765
rect 19241 6762 19307 6765
rect 17769 6760 19307 6762
rect 17769 6704 17774 6760
rect 17830 6704 19246 6760
rect 19302 6704 19307 6760
rect 17769 6702 19307 6704
rect 17769 6699 17835 6702
rect 19241 6699 19307 6702
rect 20253 6762 20319 6765
rect 25773 6762 25839 6765
rect 20253 6760 25839 6762
rect 20253 6704 20258 6760
rect 20314 6704 25778 6760
rect 25834 6704 25839 6760
rect 20253 6702 25839 6704
rect 20253 6699 20319 6702
rect 25773 6699 25839 6702
rect 31017 6762 31083 6765
rect 36537 6762 36603 6765
rect 31017 6760 36603 6762
rect 31017 6704 31022 6760
rect 31078 6704 36542 6760
rect 36598 6704 36603 6760
rect 31017 6702 36603 6704
rect 31017 6699 31083 6702
rect 36537 6699 36603 6702
rect 16573 6626 16639 6629
rect 18505 6626 18571 6629
rect 16573 6624 18571 6626
rect 16573 6568 16578 6624
rect 16634 6568 18510 6624
rect 18566 6568 18571 6624
rect 16573 6566 18571 6568
rect 16573 6563 16639 6566
rect 18505 6563 18571 6566
rect 28809 6626 28875 6629
rect 31017 6626 31083 6629
rect 28809 6624 31083 6626
rect 28809 6568 28814 6624
rect 28870 6568 31022 6624
rect 31078 6568 31083 6624
rect 28809 6566 31083 6568
rect 28809 6563 28875 6566
rect 31017 6563 31083 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 27429 6490 27495 6493
rect 34605 6490 34671 6493
rect 27429 6488 34671 6490
rect 27429 6432 27434 6488
rect 27490 6432 34610 6488
rect 34666 6432 34671 6488
rect 27429 6430 34671 6432
rect 27429 6427 27495 6430
rect 34605 6427 34671 6430
rect 17953 6354 18019 6357
rect 29085 6354 29151 6357
rect 17953 6352 29151 6354
rect 17953 6296 17958 6352
rect 18014 6296 29090 6352
rect 29146 6296 29151 6352
rect 17953 6294 29151 6296
rect 17953 6291 18019 6294
rect 29085 6291 29151 6294
rect 29269 6354 29335 6357
rect 31109 6354 31175 6357
rect 29269 6352 31175 6354
rect 29269 6296 29274 6352
rect 29330 6296 31114 6352
rect 31170 6296 31175 6352
rect 29269 6294 31175 6296
rect 29269 6291 29335 6294
rect 31109 6291 31175 6294
rect 21725 6218 21791 6221
rect 26509 6218 26575 6221
rect 21725 6216 26575 6218
rect 21725 6160 21730 6216
rect 21786 6160 26514 6216
rect 26570 6160 26575 6216
rect 21725 6158 26575 6160
rect 21725 6155 21791 6158
rect 26509 6155 26575 6158
rect 38193 6218 38259 6221
rect 39200 6218 39800 6248
rect 38193 6216 39800 6218
rect 38193 6160 38198 6216
rect 38254 6160 39800 6216
rect 38193 6158 39800 6160
rect 38193 6155 38259 6158
rect 39200 6128 39800 6158
rect 19517 6082 19583 6085
rect 22369 6082 22435 6085
rect 19517 6080 22435 6082
rect 19517 6024 19522 6080
rect 19578 6024 22374 6080
rect 22430 6024 22435 6080
rect 19517 6022 22435 6024
rect 19517 6019 19583 6022
rect 22369 6019 22435 6022
rect 29821 6082 29887 6085
rect 31477 6082 31543 6085
rect 29821 6080 31543 6082
rect 29821 6024 29826 6080
rect 29882 6024 31482 6080
rect 31538 6024 31543 6080
rect 29821 6022 31543 6024
rect 29821 6019 29887 6022
rect 31477 6019 31543 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 21909 5946 21975 5949
rect 22093 5946 22159 5949
rect 21909 5944 22159 5946
rect 21909 5888 21914 5944
rect 21970 5888 22098 5944
rect 22154 5888 22159 5944
rect 21909 5886 22159 5888
rect 21909 5883 21975 5886
rect 22093 5883 22159 5886
rect 29453 5946 29519 5949
rect 34145 5946 34211 5949
rect 29453 5944 34211 5946
rect 29453 5888 29458 5944
rect 29514 5888 34150 5944
rect 34206 5888 34211 5944
rect 29453 5886 34211 5888
rect 29453 5883 29519 5886
rect 34145 5883 34211 5886
rect 17677 5810 17743 5813
rect 29913 5810 29979 5813
rect 17677 5808 29979 5810
rect 17677 5752 17682 5808
rect 17738 5752 29918 5808
rect 29974 5752 29979 5808
rect 17677 5750 29979 5752
rect 17677 5747 17743 5750
rect 29913 5747 29979 5750
rect 15009 5674 15075 5677
rect 20437 5674 20503 5677
rect 15009 5672 20503 5674
rect 15009 5616 15014 5672
rect 15070 5616 20442 5672
rect 20498 5616 20503 5672
rect 15009 5614 20503 5616
rect 15009 5611 15075 5614
rect 20437 5611 20503 5614
rect 20805 5538 20871 5541
rect 24577 5538 24643 5541
rect 20805 5536 24643 5538
rect 20805 5480 20810 5536
rect 20866 5480 24582 5536
rect 24638 5480 24643 5536
rect 20805 5478 24643 5480
rect 20805 5475 20871 5478
rect 24577 5475 24643 5478
rect 29637 5538 29703 5541
rect 37917 5538 37983 5541
rect 29637 5536 37983 5538
rect 29637 5480 29642 5536
rect 29698 5480 37922 5536
rect 37978 5480 37983 5536
rect 29637 5478 37983 5480
rect 29637 5475 29703 5478
rect 37917 5475 37983 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 14365 5402 14431 5405
rect 16614 5402 16620 5404
rect 14365 5400 16620 5402
rect 14365 5344 14370 5400
rect 14426 5344 16620 5400
rect 14365 5342 16620 5344
rect 14365 5339 14431 5342
rect 16614 5340 16620 5342
rect 16684 5340 16690 5404
rect 20621 5402 20687 5405
rect 22185 5402 22251 5405
rect 20621 5400 22251 5402
rect 20621 5344 20626 5400
rect 20682 5344 22190 5400
rect 22246 5344 22251 5400
rect 20621 5342 22251 5344
rect 20621 5339 20687 5342
rect 22185 5339 22251 5342
rect 29913 5402 29979 5405
rect 31937 5402 32003 5405
rect 29913 5400 32003 5402
rect 29913 5344 29918 5400
rect 29974 5344 31942 5400
rect 31998 5344 32003 5400
rect 29913 5342 32003 5344
rect 29913 5339 29979 5342
rect 31937 5339 32003 5342
rect 19241 5266 19307 5269
rect 21633 5266 21699 5269
rect 19241 5264 21699 5266
rect 19241 5208 19246 5264
rect 19302 5208 21638 5264
rect 21694 5208 21699 5264
rect 19241 5206 21699 5208
rect 19241 5203 19307 5206
rect 21633 5203 21699 5206
rect 24301 5266 24367 5269
rect 25129 5266 25195 5269
rect 24301 5264 25195 5266
rect 24301 5208 24306 5264
rect 24362 5208 25134 5264
rect 25190 5208 25195 5264
rect 24301 5206 25195 5208
rect 24301 5203 24367 5206
rect 25129 5203 25195 5206
rect 31569 5266 31635 5269
rect 34513 5266 34579 5269
rect 31569 5264 34579 5266
rect 31569 5208 31574 5264
rect 31630 5208 34518 5264
rect 34574 5208 34579 5264
rect 31569 5206 34579 5208
rect 31569 5203 31635 5206
rect 34513 5203 34579 5206
rect 12433 5130 12499 5133
rect 24761 5130 24827 5133
rect 12433 5128 24827 5130
rect 12433 5072 12438 5128
rect 12494 5072 24766 5128
rect 24822 5072 24827 5128
rect 12433 5070 24827 5072
rect 12433 5067 12499 5070
rect 24761 5067 24827 5070
rect 31293 5130 31359 5133
rect 33777 5130 33843 5133
rect 31293 5128 33843 5130
rect 31293 5072 31298 5128
rect 31354 5072 33782 5128
rect 33838 5072 33843 5128
rect 31293 5070 33843 5072
rect 31293 5067 31359 5070
rect 33777 5067 33843 5070
rect 22921 4994 22987 4997
rect 33133 4994 33199 4997
rect 22921 4992 33199 4994
rect 22921 4936 22926 4992
rect 22982 4936 33138 4992
rect 33194 4936 33199 4992
rect 22921 4934 33199 4936
rect 22921 4931 22987 4934
rect 33133 4931 33199 4934
rect 4210 4928 4526 4929
rect 200 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 1669 4858 1735 4861
rect 200 4856 1735 4858
rect 200 4800 1674 4856
rect 1730 4800 1735 4856
rect 200 4798 1735 4800
rect 200 4768 800 4798
rect 1669 4795 1735 4798
rect 12341 4858 12407 4861
rect 19149 4858 19215 4861
rect 12341 4856 19215 4858
rect 12341 4800 12346 4856
rect 12402 4800 19154 4856
rect 19210 4800 19215 4856
rect 12341 4798 19215 4800
rect 12341 4795 12407 4798
rect 19149 4795 19215 4798
rect 23473 4858 23539 4861
rect 26693 4858 26759 4861
rect 23473 4856 26759 4858
rect 23473 4800 23478 4856
rect 23534 4800 26698 4856
rect 26754 4800 26759 4856
rect 23473 4798 26759 4800
rect 23473 4795 23539 4798
rect 26693 4795 26759 4798
rect 29453 4858 29519 4861
rect 32213 4858 32279 4861
rect 29453 4856 32279 4858
rect 29453 4800 29458 4856
rect 29514 4800 32218 4856
rect 32274 4800 32279 4856
rect 29453 4798 32279 4800
rect 29453 4795 29519 4798
rect 32213 4795 32279 4798
rect 38101 4858 38167 4861
rect 39200 4858 39800 4888
rect 38101 4856 39800 4858
rect 38101 4800 38106 4856
rect 38162 4800 39800 4856
rect 38101 4798 39800 4800
rect 38101 4795 38167 4798
rect 39200 4768 39800 4798
rect 19425 4722 19491 4725
rect 26785 4722 26851 4725
rect 19425 4720 26851 4722
rect 19425 4664 19430 4720
rect 19486 4664 26790 4720
rect 26846 4664 26851 4720
rect 19425 4662 26851 4664
rect 19425 4659 19491 4662
rect 26785 4659 26851 4662
rect 15837 4586 15903 4589
rect 16665 4586 16731 4589
rect 15837 4584 16731 4586
rect 15837 4528 15842 4584
rect 15898 4528 16670 4584
rect 16726 4528 16731 4584
rect 15837 4526 16731 4528
rect 15837 4523 15903 4526
rect 16665 4523 16731 4526
rect 17217 4586 17283 4589
rect 32029 4586 32095 4589
rect 17217 4584 32095 4586
rect 17217 4528 17222 4584
rect 17278 4528 32034 4584
rect 32090 4528 32095 4584
rect 17217 4526 32095 4528
rect 17217 4523 17283 4526
rect 32029 4523 32095 4526
rect 21081 4450 21147 4453
rect 34973 4450 35039 4453
rect 21081 4448 35039 4450
rect 21081 4392 21086 4448
rect 21142 4392 34978 4448
rect 35034 4392 35039 4448
rect 21081 4390 35039 4392
rect 21081 4387 21147 4390
rect 34973 4387 35039 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 12249 4178 12315 4181
rect 24945 4178 25011 4181
rect 12249 4176 25011 4178
rect 12249 4120 12254 4176
rect 12310 4120 24950 4176
rect 25006 4120 25011 4176
rect 12249 4118 25011 4120
rect 12249 4115 12315 4118
rect 24945 4115 25011 4118
rect 16113 4042 16179 4045
rect 17861 4042 17927 4045
rect 16113 4040 17927 4042
rect 16113 3984 16118 4040
rect 16174 3984 17866 4040
rect 17922 3984 17927 4040
rect 16113 3982 17927 3984
rect 16113 3979 16179 3982
rect 17861 3979 17927 3982
rect 19057 4042 19123 4045
rect 22369 4042 22435 4045
rect 23197 4044 23263 4045
rect 23197 4042 23244 4044
rect 19057 4040 22435 4042
rect 19057 3984 19062 4040
rect 19118 3984 22374 4040
rect 22430 3984 22435 4040
rect 19057 3982 22435 3984
rect 23152 4040 23244 4042
rect 23152 3984 23202 4040
rect 23152 3982 23244 3984
rect 19057 3979 19123 3982
rect 22369 3979 22435 3982
rect 23197 3980 23244 3982
rect 23308 3980 23314 4044
rect 23197 3979 23263 3980
rect 22093 3906 22159 3909
rect 26601 3906 26667 3909
rect 22093 3904 26667 3906
rect 22093 3848 22098 3904
rect 22154 3848 26606 3904
rect 26662 3848 26667 3904
rect 22093 3846 26667 3848
rect 22093 3843 22159 3846
rect 26601 3843 26667 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 31201 3770 31267 3773
rect 34789 3770 34855 3773
rect 31201 3768 34855 3770
rect 31201 3712 31206 3768
rect 31262 3712 34794 3768
rect 34850 3712 34855 3768
rect 31201 3710 34855 3712
rect 31201 3707 31267 3710
rect 34789 3707 34855 3710
rect 21173 3634 21239 3637
rect 22093 3634 22159 3637
rect 21173 3632 22159 3634
rect 21173 3576 21178 3632
rect 21234 3576 22098 3632
rect 22154 3576 22159 3632
rect 21173 3574 22159 3576
rect 21173 3571 21239 3574
rect 22093 3571 22159 3574
rect 29637 3634 29703 3637
rect 30925 3634 30991 3637
rect 32029 3634 32095 3637
rect 29637 3632 32095 3634
rect 29637 3576 29642 3632
rect 29698 3576 30930 3632
rect 30986 3576 32034 3632
rect 32090 3576 32095 3632
rect 29637 3574 32095 3576
rect 29637 3571 29703 3574
rect 30925 3571 30991 3574
rect 32029 3571 32095 3574
rect 32305 3634 32371 3637
rect 33777 3634 33843 3637
rect 32305 3632 33843 3634
rect 32305 3576 32310 3632
rect 32366 3576 33782 3632
rect 33838 3576 33843 3632
rect 32305 3574 33843 3576
rect 32305 3571 32371 3574
rect 33777 3571 33843 3574
rect 200 3498 800 3528
rect 1669 3498 1735 3501
rect 200 3496 1735 3498
rect 200 3440 1674 3496
rect 1730 3440 1735 3496
rect 200 3438 1735 3440
rect 200 3408 800 3438
rect 1669 3435 1735 3438
rect 13721 3498 13787 3501
rect 19977 3498 20043 3501
rect 13721 3496 20043 3498
rect 13721 3440 13726 3496
rect 13782 3440 19982 3496
rect 20038 3440 20043 3496
rect 13721 3438 20043 3440
rect 13721 3435 13787 3438
rect 19977 3435 20043 3438
rect 27797 3498 27863 3501
rect 34513 3498 34579 3501
rect 27797 3496 34579 3498
rect 27797 3440 27802 3496
rect 27858 3440 34518 3496
rect 34574 3440 34579 3496
rect 27797 3438 34579 3440
rect 27797 3435 27863 3438
rect 34513 3435 34579 3438
rect 22185 3362 22251 3365
rect 34145 3362 34211 3365
rect 22185 3360 34211 3362
rect 22185 3304 22190 3360
rect 22246 3304 34150 3360
rect 34206 3304 34211 3360
rect 22185 3302 34211 3304
rect 22185 3299 22251 3302
rect 34145 3299 34211 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 20897 3226 20963 3229
rect 22185 3226 22251 3229
rect 26509 3226 26575 3229
rect 20897 3224 22251 3226
rect 20897 3168 20902 3224
rect 20958 3168 22190 3224
rect 22246 3168 22251 3224
rect 20897 3166 22251 3168
rect 20897 3163 20963 3166
rect 22185 3163 22251 3166
rect 22326 3224 26575 3226
rect 22326 3168 26514 3224
rect 26570 3168 26575 3224
rect 22326 3166 26575 3168
rect 19977 3090 20043 3093
rect 22326 3090 22386 3166
rect 26509 3163 26575 3166
rect 31661 3226 31727 3229
rect 32397 3226 32463 3229
rect 34421 3226 34487 3229
rect 31661 3224 34487 3226
rect 31661 3168 31666 3224
rect 31722 3168 32402 3224
rect 32458 3168 34426 3224
rect 34482 3168 34487 3224
rect 31661 3166 34487 3168
rect 31661 3163 31727 3166
rect 32397 3163 32463 3166
rect 34421 3163 34487 3166
rect 19977 3088 22386 3090
rect 19977 3032 19982 3088
rect 20038 3032 22386 3088
rect 19977 3030 22386 3032
rect 23381 3090 23447 3093
rect 34973 3090 35039 3093
rect 23381 3088 35039 3090
rect 23381 3032 23386 3088
rect 23442 3032 34978 3088
rect 35034 3032 35039 3088
rect 23381 3030 35039 3032
rect 19977 3027 20043 3030
rect 23381 3027 23447 3030
rect 34973 3027 35039 3030
rect 21357 2954 21423 2957
rect 26785 2954 26851 2957
rect 21357 2952 26851 2954
rect 21357 2896 21362 2952
rect 21418 2896 26790 2952
rect 26846 2896 26851 2952
rect 21357 2894 26851 2896
rect 21357 2891 21423 2894
rect 26785 2891 26851 2894
rect 30189 2954 30255 2957
rect 34237 2954 34303 2957
rect 30189 2952 34303 2954
rect 30189 2896 30194 2952
rect 30250 2896 34242 2952
rect 34298 2896 34303 2952
rect 30189 2894 34303 2896
rect 30189 2891 30255 2894
rect 34237 2891 34303 2894
rect 38193 2818 38259 2821
rect 39200 2818 39800 2848
rect 38193 2816 39800 2818
rect 38193 2760 38198 2816
rect 38254 2760 39800 2816
rect 38193 2758 39800 2760
rect 38193 2755 38259 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 39200 2728 39800 2758
rect 34930 2687 35246 2688
rect 18873 2682 18939 2685
rect 21398 2682 21404 2684
rect 18873 2680 21404 2682
rect 18873 2624 18878 2680
rect 18934 2624 21404 2680
rect 18873 2622 21404 2624
rect 18873 2619 18939 2622
rect 21398 2620 21404 2622
rect 21468 2620 21474 2684
rect 4061 2546 4127 2549
rect 17350 2546 17356 2548
rect 4061 2544 17356 2546
rect 4061 2488 4066 2544
rect 4122 2488 17356 2544
rect 4061 2486 17356 2488
rect 4061 2483 4127 2486
rect 17350 2484 17356 2486
rect 17420 2484 17426 2548
rect 31293 2546 31359 2549
rect 36169 2546 36235 2549
rect 31293 2544 36235 2546
rect 31293 2488 31298 2544
rect 31354 2488 36174 2544
rect 36230 2488 36235 2544
rect 31293 2486 36235 2488
rect 31293 2483 31359 2486
rect 36169 2483 36235 2486
rect 20621 2410 20687 2413
rect 36261 2410 36327 2413
rect 20621 2408 36327 2410
rect 20621 2352 20626 2408
rect 20682 2352 36266 2408
rect 36322 2352 36327 2408
rect 20621 2350 36327 2352
rect 20621 2347 20687 2350
rect 36261 2347 36327 2350
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 200 1458 800 1488
rect 2773 1458 2839 1461
rect 200 1456 2839 1458
rect 200 1400 2778 1456
rect 2834 1400 2839 1456
rect 200 1398 2839 1400
rect 200 1368 800 1398
rect 2773 1395 2839 1398
rect 37181 1458 37247 1461
rect 37181 1456 39314 1458
rect 37181 1400 37186 1456
rect 37242 1400 39314 1456
rect 37181 1398 39314 1400
rect 37181 1395 37247 1398
rect 39254 1050 39314 1398
rect 39070 990 39314 1050
rect 39070 778 39130 990
rect 39200 778 39800 808
rect 39070 718 39800 778
rect 39200 688 39800 718
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 23244 17580 23308 17644
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 21404 15268 21468 15332
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 17356 12820 17420 12884
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 16620 7788 16684 7852
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 16620 5340 16684 5404
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 23244 4040 23308 4044
rect 23244 3984 23258 4040
rect 23258 3984 23308 4040
rect 23244 3980 23308 3984
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 21404 2620 21468 2684
rect 17356 2484 17420 2548
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 23243 17644 23309 17645
rect 23243 17580 23244 17644
rect 23308 17580 23309 17644
rect 23243 17579 23309 17580
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 21403 15332 21469 15333
rect 21403 15268 21404 15332
rect 21468 15268 21469 15332
rect 21403 15267 21469 15268
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 17355 12884 17421 12885
rect 17355 12820 17356 12884
rect 17420 12820 17421 12884
rect 17355 12819 17421 12820
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 16619 7852 16685 7853
rect 16619 7788 16620 7852
rect 16684 7788 16685 7852
rect 16619 7787 16685 7788
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 16622 5405 16682 7787
rect 16619 5404 16685 5405
rect 16619 5340 16620 5404
rect 16684 5340 16685 5404
rect 16619 5339 16685 5340
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 17358 2549 17418 12819
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 17355 2548 17421 2549
rect 17355 2484 17356 2548
rect 17420 2484 17421 2548
rect 17355 2483 17421 2484
rect 19568 2208 19888 3232
rect 21406 2685 21466 15267
rect 23246 4045 23306 17579
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 23243 4044 23309 4045
rect 23243 3980 23244 4044
rect 23308 3980 23309 4044
rect 23243 3979 23309 3980
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 21403 2684 21469 2685
rect 21403 2620 21404 2684
rect 21468 2620 21469 2684
rect 21403 2619 21469 2620
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 19688 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__A
timestamp 1667941163
transform -1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A
timestamp 1667941163
transform 1 0 32108 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A
timestamp 1667941163
transform 1 0 23920 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__A
timestamp 1667941163
transform -1 0 18492 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__A
timestamp 1667941163
transform -1 0 12696 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__232__A
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A
timestamp 1667941163
transform -1 0 12696 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1667941163
transform -1 0 23000 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A
timestamp 1667941163
transform -1 0 33028 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A
timestamp 1667941163
transform -1 0 31188 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1667941163
transform -1 0 33120 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A
timestamp 1667941163
transform -1 0 33120 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A
timestamp 1667941163
transform -1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A
timestamp 1667941163
transform -1 0 17940 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1667941163
transform -1 0 14628 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A
timestamp 1667941163
transform -1 0 25944 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__A
timestamp 1667941163
transform -1 0 27876 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__A
timestamp 1667941163
transform -1 0 30452 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A
timestamp 1667941163
transform -1 0 22264 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A
timestamp 1667941163
transform 1 0 27140 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A
timestamp 1667941163
transform 1 0 20700 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A
timestamp 1667941163
transform -1 0 21712 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A
timestamp 1667941163
transform 1 0 19872 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A
timestamp 1667941163
transform 1 0 18768 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A
timestamp 1667941163
transform -1 0 14076 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__A
timestamp 1667941163
transform -1 0 26864 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A
timestamp 1667941163
transform -1 0 28980 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A
timestamp 1667941163
transform -1 0 29900 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__A
timestamp 1667941163
transform -1 0 13984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A
timestamp 1667941163
transform -1 0 15732 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__A
timestamp 1667941163
transform 1 0 14996 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A
timestamp 1667941163
transform -1 0 29808 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__A
timestamp 1667941163
transform -1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__A
timestamp 1667941163
transform -1 0 12972 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A
timestamp 1667941163
transform -1 0 29072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A
timestamp 1667941163
transform -1 0 14628 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__A
timestamp 1667941163
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__A
timestamp 1667941163
transform -1 0 18584 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__A
timestamp 1667941163
transform 1 0 32660 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__A
timestamp 1667941163
transform -1 0 31188 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__A
timestamp 1667941163
transform 1 0 19596 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A
timestamp 1667941163
transform -1 0 33120 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__A
timestamp 1667941163
transform -1 0 13248 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__A
timestamp 1667941163
transform -1 0 11224 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__A
timestamp 1667941163
transform 1 0 17848 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A
timestamp 1667941163
transform -1 0 31556 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__A
timestamp 1667941163
transform -1 0 13156 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__A
timestamp 1667941163
transform 1 0 17756 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__A
timestamp 1667941163
transform 1 0 14996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A
timestamp 1667941163
transform -1 0 29624 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__A
timestamp 1667941163
transform 1 0 29072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__A
timestamp 1667941163
transform 1 0 18952 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__A
timestamp 1667941163
transform -1 0 13340 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__A
timestamp 1667941163
transform -1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__A
timestamp 1667941163
transform 1 0 32292 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__A
timestamp 1667941163
transform -1 0 30360 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A
timestamp 1667941163
transform 1 0 13708 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__A
timestamp 1667941163
transform -1 0 33580 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__A
timestamp 1667941163
transform 1 0 13248 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__A
timestamp 1667941163
transform -1 0 13248 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__A
timestamp 1667941163
transform -1 0 13524 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__A
timestamp 1667941163
transform 1 0 19320 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__A
timestamp 1667941163
transform -1 0 15732 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__A
timestamp 1667941163
transform -1 0 13156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__A
timestamp 1667941163
transform 1 0 21528 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__A
timestamp 1667941163
transform -1 0 17848 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__A
timestamp 1667941163
transform -1 0 31740 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__A
timestamp 1667941163
transform -1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A
timestamp 1667941163
transform 1 0 23828 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__344__A
timestamp 1667941163
transform 1 0 2944 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A
timestamp 1667941163
transform 1 0 18216 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A
timestamp 1667941163
transform 1 0 28244 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__A
timestamp 1667941163
transform 1 0 32292 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__A
timestamp 1667941163
transform -1 0 27876 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__A
timestamp 1667941163
transform -1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__A
timestamp 1667941163
transform 1 0 20148 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__A
timestamp 1667941163
transform -1 0 12144 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__A
timestamp 1667941163
transform -1 0 10948 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__A
timestamp 1667941163
transform 1 0 18860 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__A
timestamp 1667941163
transform 1 0 32844 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__365__A
timestamp 1667941163
transform -1 0 35696 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__A
timestamp 1667941163
transform 1 0 23460 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__A
timestamp 1667941163
transform 1 0 13156 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__A
timestamp 1667941163
transform -1 0 12420 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1667941163
transform -1 0 15180 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__371__A
timestamp 1667941163
transform 1 0 19412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__373__A
timestamp 1667941163
transform 1 0 10488 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A
timestamp 1667941163
transform 1 0 16192 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__375__A
timestamp 1667941163
transform 1 0 29716 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__A
timestamp 1667941163
transform 1 0 18584 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__A
timestamp 1667941163
transform 1 0 19688 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__383__A
timestamp 1667941163
transform -1 0 27968 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1667941163
transform -1 0 20700 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__A
timestamp 1667941163
transform 1 0 5244 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__387__A
timestamp 1667941163
transform 1 0 13616 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__389__A
timestamp 1667941163
transform 1 0 11776 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__A
timestamp 1667941163
transform -1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__391__A
timestamp 1667941163
transform 1 0 11592 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__393__A
timestamp 1667941163
transform 1 0 35052 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__A
timestamp 1667941163
transform 1 0 37076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__395__A
timestamp 1667941163
transform 1 0 33948 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A
timestamp 1667941163
transform -1 0 38364 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__A
timestamp 1667941163
transform 1 0 33396 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__A
timestamp 1667941163
transform 1 0 37076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__A
timestamp 1667941163
transform -1 0 38088 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__A
timestamp 1667941163
transform 1 0 37444 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__A
timestamp 1667941163
transform 1 0 37628 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__402__A
timestamp 1667941163
transform 1 0 36708 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__A
timestamp 1667941163
transform 1 0 36524 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__A
timestamp 1667941163
transform 1 0 37996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__A
timestamp 1667941163
transform 1 0 35328 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__407__A
timestamp 1667941163
transform 1 0 35604 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__A
timestamp 1667941163
transform 1 0 36800 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__A
timestamp 1667941163
transform 1 0 34868 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__A
timestamp 1667941163
transform 1 0 37076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__A
timestamp 1667941163
transform 1 0 34684 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__A
timestamp 1667941163
transform 1 0 37628 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__413__A
timestamp 1667941163
transform -1 0 38088 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__415__A
timestamp 1667941163
transform 1 0 35972 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A
timestamp 1667941163
transform 1 0 37628 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__A
timestamp 1667941163
transform 1 0 35052 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__A
timestamp 1667941163
transform 1 0 36248 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__419__A
timestamp 1667941163
transform 1 0 35972 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__A
timestamp 1667941163
transform -1 0 35144 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__421__A
timestamp 1667941163
transform -1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__A
timestamp 1667941163
transform 1 0 34500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__A
timestamp 1667941163
transform 1 0 34868 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__A
timestamp 1667941163
transform 1 0 37076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__A
timestamp 1667941163
transform -1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__A
timestamp 1667941163
transform 1 0 36708 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__A
timestamp 1667941163
transform -1 0 37444 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__429__A
timestamp 1667941163
transform 1 0 36524 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__A
timestamp 1667941163
transform 1 0 35420 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__A
timestamp 1667941163
transform 1 0 37628 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__A
timestamp 1667941163
transform 1 0 36524 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__A
timestamp 1667941163
transform 1 0 36156 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__A
timestamp 1667941163
transform 1 0 35420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__435__A
timestamp 1667941163
transform 1 0 37444 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__A
timestamp 1667941163
transform 1 0 11040 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__A
timestamp 1667941163
transform 1 0 12880 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__A
timestamp 1667941163
transform 1 0 14536 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__449__A
timestamp 1667941163
transform 1 0 13800 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__A
timestamp 1667941163
transform 1 0 13616 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__A
timestamp 1667941163
transform 1 0 12328 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__452__A
timestamp 1667941163
transform -1 0 35604 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__453__A
timestamp 1667941163
transform 1 0 11776 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__A
timestamp 1667941163
transform 1 0 13156 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__455__A
timestamp 1667941163
transform 1 0 13064 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__456__A
timestamp 1667941163
transform -1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__457__A
timestamp 1667941163
transform 1 0 15088 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__464__CLK
timestamp 1667941163
transform 1 0 18584 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__CLK
timestamp 1667941163
transform 1 0 11040 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__CLK
timestamp 1667941163
transform 1 0 18216 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__D
timestamp 1667941163
transform -1 0 27324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__CLK
timestamp 1667941163
transform 1 0 29624 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__CLK
timestamp 1667941163
transform 1 0 27692 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__D
timestamp 1667941163
transform -1 0 29900 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__CLK
timestamp 1667941163
transform 1 0 31280 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__CLK
timestamp 1667941163
transform 1 0 33304 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__471__CLK
timestamp 1667941163
transform 1 0 33672 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__472__CLK
timestamp 1667941163
transform 1 0 35420 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__473__CLK
timestamp 1667941163
transform 1 0 34500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__CLK
timestamp 1667941163
transform 1 0 32292 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__CLK
timestamp 1667941163
transform 1 0 31096 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__D
timestamp 1667941163
transform -1 0 32108 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__476__CLK
timestamp 1667941163
transform 1 0 19504 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__477__CLK
timestamp 1667941163
transform 1 0 22816 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__CLK
timestamp 1667941163
transform 1 0 18768 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__D
timestamp 1667941163
transform -1 0 17020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__479__CLK
timestamp 1667941163
transform 1 0 30268 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__479__D
timestamp 1667941163
transform 1 0 30728 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__CLK
timestamp 1667941163
transform 1 0 31372 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__D
timestamp 1667941163
transform 1 0 29440 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__481__CLK
timestamp 1667941163
transform 1 0 12880 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__CLK
timestamp 1667941163
transform 1 0 32844 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__483__CLK
timestamp 1667941163
transform 1 0 33120 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__CLK
timestamp 1667941163
transform 1 0 35604 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__485__CLK
timestamp 1667941163
transform 1 0 30820 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__CLK
timestamp 1667941163
transform 1 0 28888 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__D
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__487__CLK
timestamp 1667941163
transform 1 0 33396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__488__CLK
timestamp 1667941163
transform 1 0 30544 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__489__CLK
timestamp 1667941163
transform 1 0 19136 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__CLK
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__D
timestamp 1667941163
transform 1 0 17480 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__RESET_B
timestamp 1667941163
transform -1 0 13156 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__491__CLK
timestamp 1667941163
transform 1 0 33028 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__491__D
timestamp 1667941163
transform 1 0 18584 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__CLK
timestamp 1667941163
transform 1 0 18216 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__D
timestamp 1667941163
transform 1 0 28060 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__CLK
timestamp 1667941163
transform 1 0 34868 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__CLK
timestamp 1667941163
transform 1 0 36156 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__495__CLK
timestamp 1667941163
transform 1 0 35604 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__CLK
timestamp 1667941163
transform 1 0 34224 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__D
timestamp 1667941163
transform -1 0 34040 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__CLK
timestamp 1667941163
transform 1 0 32200 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__D
timestamp 1667941163
transform 1 0 29716 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__CLK
timestamp 1667941163
transform 1 0 28980 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__D
timestamp 1667941163
transform 1 0 23920 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__499__CLK
timestamp 1667941163
transform 1 0 38180 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__500__CLK
timestamp 1667941163
transform 1 0 33856 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__501__CLK
timestamp 1667941163
transform 1 0 32292 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__502__CLK
timestamp 1667941163
transform 1 0 32476 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__502__D
timestamp 1667941163
transform -1 0 33028 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__503__CLK
timestamp 1667941163
transform 1 0 30820 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__503__D
timestamp 1667941163
transform -1 0 30728 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__504__CLK
timestamp 1667941163
transform 1 0 32568 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__504__D
timestamp 1667941163
transform -1 0 32200 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__505__CLK
timestamp 1667941163
transform 1 0 37444 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__506__CLK
timestamp 1667941163
transform 1 0 34132 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__507__CLK
timestamp 1667941163
transform 1 0 32844 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__508__CLK
timestamp 1667941163
transform 1 0 23368 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__508__D
timestamp 1667941163
transform -1 0 23000 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__509__CLK
timestamp 1667941163
transform 1 0 21988 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__509__D
timestamp 1667941163
transform -1 0 21068 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__510__CLK
timestamp 1667941163
transform 1 0 31648 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__511__CLK
timestamp 1667941163
transform 1 0 31924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__512__CLK
timestamp 1667941163
transform 1 0 32568 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__512__D
timestamp 1667941163
transform -1 0 36156 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__513__CLK
timestamp 1667941163
transform 1 0 33948 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__514__CLK
timestamp 1667941163
transform 1 0 28336 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__514__D
timestamp 1667941163
transform 1 0 23460 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__515__CLK
timestamp 1667941163
transform 1 0 20056 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__515__D
timestamp 1667941163
transform -1 0 26956 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__516__CLK
timestamp 1667941163
transform 1 0 29992 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__516__D
timestamp 1667941163
transform 1 0 30268 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__517__CLK
timestamp 1667941163
transform 1 0 34868 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__518__CLK
timestamp 1667941163
transform 1 0 30452 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__519__CLK
timestamp 1667941163
transform 1 0 19136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__520__CLK
timestamp 1667941163
transform 1 0 33396 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__520__D
timestamp 1667941163
transform -1 0 27692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__521__CLK
timestamp 1667941163
transform 1 0 28244 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__522__CLK
timestamp 1667941163
transform 1 0 27140 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__522__D
timestamp 1667941163
transform -1 0 23276 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__523__CLK
timestamp 1667941163
transform 1 0 32752 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__523__RESET_B
timestamp 1667941163
transform -1 0 32476 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__524__CLK
timestamp 1667941163
transform 1 0 35052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__525__CLK
timestamp 1667941163
transform 1 0 37444 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__CLK
timestamp 1667941163
transform 1 0 33580 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__527__CLK
timestamp 1667941163
transform 1 0 31280 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__528__CLK
timestamp 1667941163
transform 1 0 22540 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__529__CLK
timestamp 1667941163
transform 1 0 33948 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__541__A
timestamp 1667941163
transform -1 0 10580 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__542__A
timestamp 1667941163
transform 1 0 7544 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__543__A
timestamp 1667941163
transform -1 0 3128 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__544__A
timestamp 1667941163
transform -1 0 27968 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__545__A
timestamp 1667941163
transform -1 0 15640 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__546__A
timestamp 1667941163
transform 1 0 18124 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__547__A
timestamp 1667941163
transform -1 0 33396 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__548__A
timestamp 1667941163
transform 1 0 24564 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__549__A
timestamp 1667941163
transform -1 0 17756 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__550__A
timestamp 1667941163
transform 1 0 6992 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__551__A
timestamp 1667941163
transform 1 0 23552 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__555__A
timestamp 1667941163
transform 1 0 24932 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__556__A
timestamp 1667941163
transform 1 0 31556 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__557__A
timestamp 1667941163
transform -1 0 28520 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__558__A
timestamp 1667941163
transform 1 0 27784 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__560__A
timestamp 1667941163
transform -1 0 8004 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__562__A
timestamp 1667941163
transform 1 0 14352 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__564__A
timestamp 1667941163
transform -1 0 31004 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__566__A
timestamp 1667941163
transform -1 0 9936 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__567__A
timestamp 1667941163
transform -1 0 6716 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__572__A
timestamp 1667941163
transform -1 0 23828 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__573__A
timestamp 1667941163
transform -1 0 36800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__574__A
timestamp 1667941163
transform 1 0 25576 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__575__A
timestamp 1667941163
transform -1 0 15824 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__613__A
timestamp 1667941163
transform -1 0 12880 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__621__A
timestamp 1667941163
transform 1 0 15548 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__628__A
timestamp 1667941163
transform -1 0 13708 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__668__A
timestamp 1667941163
transform 1 0 20240 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__685__A
timestamp 1667941163
transform 1 0 17020 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__693__A
timestamp 1667941163
transform 1 0 14628 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1667941163
transform -1 0 37720 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1667941163
transform -1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1667941163
transform -1 0 10672 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1667941163
transform -1 0 37628 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1667941163
transform -1 0 38364 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1667941163
transform -1 0 38364 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1667941163
transform -1 0 38364 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1667941163
transform -1 0 38364 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1667941163
transform -1 0 1748 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1667941163
transform -1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1667941163
transform -1 0 38364 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1667941163
transform -1 0 1748 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1667941163
transform -1 0 1748 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1667941163
transform -1 0 37628 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1667941163
transform -1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1667941163
transform -1 0 24840 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1667941163
transform -1 0 4140 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1667941163
transform -1 0 37628 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1667941163
transform -1 0 1748 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1667941163
transform -1 0 1748 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1667941163
transform -1 0 9844 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1667941163
transform -1 0 36248 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1667941163
transform -1 0 37628 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1667941163
transform -1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1667941163
transform -1 0 32476 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1667941163
transform -1 0 3220 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1667941163
transform -1 0 37536 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1667941163
transform -1 0 1748 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1667941163
transform -1 0 38364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1667941163
transform -1 0 1748 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1667941163
transform -1 0 34684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1667941163
transform -1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1667941163
transform -1 0 11684 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1667941163
transform -1 0 6072 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1667941163
transform -1 0 18216 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1667941163
transform -1 0 3220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1667941163
transform -1 0 29164 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1667941163
transform -1 0 14444 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1667941163
transform -1 0 23276 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1667941163
transform -1 0 9384 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output49_A
timestamp 1667941163
transform -1 0 35144 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output53_A
timestamp 1667941163
transform -1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output55_A
timestamp 1667941163
transform -1 0 35696 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output56_A
timestamp 1667941163
transform -1 0 20976 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output57_A
timestamp 1667941163
transform 1 0 37444 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output68_A
timestamp 1667941163
transform 1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output72_A
timestamp 1667941163
transform 1 0 2300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output76_A
timestamp 1667941163
transform 1 0 36432 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output78_A
timestamp 1667941163
transform -1 0 5520 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output81_A
timestamp 1667941163
transform -1 0 10672 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output82_A
timestamp 1667941163
transform -1 0 2484 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output85_A
timestamp 1667941163
transform -1 0 2484 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2484 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3036 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37
timestamp 1667941163
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4968 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1667941163
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63
timestamp 1667941163
transform 1 0 6900 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1667941163
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79
timestamp 1667941163
transform 1 0 8372 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91
timestamp 1667941163
transform 1 0 9476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_98
timestamp 1667941163
transform 1 0 10120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104
timestamp 1667941163
transform 1 0 10672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1667941163
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12052 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_127
timestamp 1667941163
transform 1 0 12788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_130
timestamp 1667941163
transform 1 0 13064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_149
timestamp 1667941163
transform 1 0 14812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_157
timestamp 1667941163
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_161
timestamp 1667941163
transform 1 0 15916 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1667941163
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_173
timestamp 1667941163
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_183
timestamp 1667941163
transform 1 0 17940 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_189
timestamp 1667941163
transform 1 0 18492 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1667941163
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_201
timestamp 1667941163
transform 1 0 19596 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1667941163
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1667941163
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1667941163
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_275
timestamp 1667941163
transform 1 0 26404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1667941163
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_285
timestamp 1667941163
transform 1 0 27324 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1667941163
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_331
timestamp 1667941163
transform 1 0 31556 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1667941163
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_359
timestamp 1667941163
transform 1 0 34132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1667941163
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_371
timestamp 1667941163
transform 1 0 35236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_379
timestamp 1667941163
transform 1 0 35972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_385
timestamp 1667941163
transform 1 0 36524 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1667941163
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_17
timestamp 1667941163
transform 1 0 2668 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_23
timestamp 1667941163
transform 1 0 3220 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_35
timestamp 1667941163
transform 1 0 4324 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_46
timestamp 1667941163
transform 1 0 5336 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1667941163
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1667941163
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_95
timestamp 1667941163
transform 1 0 9844 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_101
timestamp 1667941163
transform 1 0 10396 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_104
timestamp 1667941163
transform 1 0 10672 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1667941163
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_119
timestamp 1667941163
transform 1 0 12052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_126
timestamp 1667941163
transform 1 0 12696 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_136
timestamp 1667941163
transform 1 0 13616 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_146
timestamp 1667941163
transform 1 0 14536 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_152
timestamp 1667941163
transform 1 0 15088 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_156
timestamp 1667941163
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1667941163
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_174
timestamp 1667941163
transform 1 0 17112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_198
timestamp 1667941163
transform 1 0 19320 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1667941163
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_248
timestamp 1667941163
transform 1 0 23920 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_254
timestamp 1667941163
transform 1 0 24472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1667941163
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_287
timestamp 1667941163
transform 1 0 27508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_314
timestamp 1667941163
transform 1 0 29992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_322
timestamp 1667941163
transform 1 0 30728 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_330
timestamp 1667941163
transform 1 0 31464 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1667941163
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_359
timestamp 1667941163
transform 1 0 34132 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_366
timestamp 1667941163
transform 1 0 34776 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_373
timestamp 1667941163
transform 1 0 35420 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_380
timestamp 1667941163
transform 1 0 36064 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_387
timestamp 1667941163
transform 1 0 36708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1667941163
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_399
timestamp 1667941163
transform 1 0 37812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_9
timestamp 1667941163
transform 1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1667941163
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1667941163
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1667941163
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1667941163
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_101
timestamp 1667941163
transform 1 0 10396 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_104
timestamp 1667941163
transform 1 0 10672 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_110
timestamp 1667941163
transform 1 0 11224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_116
timestamp 1667941163
transform 1 0 11776 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_123
timestamp 1667941163
transform 1 0 12420 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_131
timestamp 1667941163
transform 1 0 13156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1667941163
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1667941163
transform 1 0 14812 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_155
timestamp 1667941163
transform 1 0 15364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_162
timestamp 1667941163
transform 1 0 16008 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_175
timestamp 1667941163
transform 1 0 17204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_185
timestamp 1667941163
transform 1 0 18124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1667941163
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_203
timestamp 1667941163
transform 1 0 19780 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_234
timestamp 1667941163
transform 1 0 22632 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_242
timestamp 1667941163
transform 1 0 23368 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1667941163
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_259
timestamp 1667941163
transform 1 0 24932 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_283
timestamp 1667941163
transform 1 0 27140 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_295
timestamp 1667941163
transform 1 0 28244 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1667941163
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_331
timestamp 1667941163
transform 1 0 31556 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_355
timestamp 1667941163
transform 1 0 33764 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp 1667941163
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_370
timestamp 1667941163
transform 1 0 35144 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_384
timestamp 1667941163
transform 1 0 36432 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_391
timestamp 1667941163
transform 1 0 37076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_397
timestamp 1667941163
transform 1 0 37628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1667941163
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1667941163
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1667941163
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1667941163
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1667941163
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_118
timestamp 1667941163
transform 1 0 11960 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_124
timestamp 1667941163
transform 1 0 12512 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_130
timestamp 1667941163
transform 1 0 13064 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_137
timestamp 1667941163
transform 1 0 13708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_150
timestamp 1667941163
transform 1 0 14904 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_157
timestamp 1667941163
transform 1 0 15548 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1667941163
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_175
timestamp 1667941163
transform 1 0 17204 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_182
timestamp 1667941163
transform 1 0 17848 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_192
timestamp 1667941163
transform 1 0 18768 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_198
timestamp 1667941163
transform 1 0 19320 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1667941163
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_247
timestamp 1667941163
transform 1 0 23828 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_271
timestamp 1667941163
transform 1 0 26036 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1667941163
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_307
timestamp 1667941163
transform 1 0 29348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_331
timestamp 1667941163
transform 1 0 31556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_359
timestamp 1667941163
transform 1 0 34132 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_366
timestamp 1667941163
transform 1 0 34776 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_380
timestamp 1667941163
transform 1 0 36064 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_387
timestamp 1667941163
transform 1 0 36708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_398
timestamp 1667941163
transform 1 0 37720 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1667941163
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_113
timestamp 1667941163
transform 1 0 11500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_117
timestamp 1667941163
transform 1 0 11868 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_124
timestamp 1667941163
transform 1 0 12512 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_131
timestamp 1667941163
transform 1 0 13156 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1667941163
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_145
timestamp 1667941163
transform 1 0 14444 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1667941163
transform 1 0 14812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_156
timestamp 1667941163
transform 1 0 15456 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_163
timestamp 1667941163
transform 1 0 16100 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_170
timestamp 1667941163
transform 1 0 16744 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_185
timestamp 1667941163
transform 1 0 18124 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_188
timestamp 1667941163
transform 1 0 18400 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1667941163
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_202
timestamp 1667941163
transform 1 0 19688 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_208
timestamp 1667941163
transform 1 0 20240 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_232
timestamp 1667941163
transform 1 0 22448 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_238
timestamp 1667941163
transform 1 0 23000 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_246
timestamp 1667941163
transform 1 0 23736 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1667941163
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_275
timestamp 1667941163
transform 1 0 26404 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_299
timestamp 1667941163
transform 1 0 28612 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_305
timestamp 1667941163
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_331
timestamp 1667941163
transform 1 0 31556 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_355
timestamp 1667941163
transform 1 0 33764 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp 1667941163
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_370
timestamp 1667941163
transform 1 0 35144 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_384
timestamp 1667941163
transform 1 0 36432 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_391
timestamp 1667941163
transform 1 0 37076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_398
timestamp 1667941163
transform 1 0 37720 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1667941163
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_9
timestamp 1667941163
transform 1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1667941163
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1667941163
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1667941163
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1667941163
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1667941163
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_97
timestamp 1667941163
transform 1 0 10028 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_103
timestamp 1667941163
transform 1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1667941163
transform 1 0 11960 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_132
timestamp 1667941163
transform 1 0 13248 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_139
timestamp 1667941163
transform 1 0 13892 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_146
timestamp 1667941163
transform 1 0 14536 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_153
timestamp 1667941163
transform 1 0 15180 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_162
timestamp 1667941163
transform 1 0 16008 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_174
timestamp 1667941163
transform 1 0 17112 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_180
timestamp 1667941163
transform 1 0 17664 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_186
timestamp 1667941163
transform 1 0 18216 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_192
timestamp 1667941163
transform 1 0 18768 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_198
timestamp 1667941163
transform 1 0 19320 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1667941163
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_229
timestamp 1667941163
transform 1 0 22172 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_235
timestamp 1667941163
transform 1 0 22724 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_241
timestamp 1667941163
transform 1 0 23276 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_285
timestamp 1667941163
transform 1 0 27324 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_316
timestamp 1667941163
transform 1 0 30176 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_322
timestamp 1667941163
transform 1 0 30728 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_330
timestamp 1667941163
transform 1 0 31464 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_334
timestamp 1667941163
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_359
timestamp 1667941163
transform 1 0 34132 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_366
timestamp 1667941163
transform 1 0 34776 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_380
timestamp 1667941163
transform 1 0 36064 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_387
timestamp 1667941163
transform 1 0 36708 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_397
timestamp 1667941163
transform 1 0 37628 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_15
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_20
timestamp 1667941163
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1667941163
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1667941163
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1667941163
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_129
timestamp 1667941163
transform 1 0 12972 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_132
timestamp 1667941163
transform 1 0 13248 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1667941163
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_148
timestamp 1667941163
transform 1 0 14720 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_154
timestamp 1667941163
transform 1 0 15272 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_164
timestamp 1667941163
transform 1 0 16192 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_171
timestamp 1667941163
transform 1 0 16836 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_178
timestamp 1667941163
transform 1 0 17480 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_188
timestamp 1667941163
transform 1 0 18400 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1667941163
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_203
timestamp 1667941163
transform 1 0 19780 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_217
timestamp 1667941163
transform 1 0 21068 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_241
timestamp 1667941163
transform 1 0 23276 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_247
timestamp 1667941163
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_275
timestamp 1667941163
transform 1 0 26404 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_281
timestamp 1667941163
transform 1 0 26956 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1667941163
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_331
timestamp 1667941163
transform 1 0 31556 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_337
timestamp 1667941163
transform 1 0 32108 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_343
timestamp 1667941163
transform 1 0 32660 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_347
timestamp 1667941163
transform 1 0 33028 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_354
timestamp 1667941163
transform 1 0 33672 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_361
timestamp 1667941163
transform 1 0 34316 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_370
timestamp 1667941163
transform 1 0 35144 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_384
timestamp 1667941163
transform 1 0 36432 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_393
timestamp 1667941163
transform 1 0 37260 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_400
timestamp 1667941163
transform 1 0 37904 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_406
timestamp 1667941163
transform 1 0 38456 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1667941163
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1667941163
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1667941163
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_133
timestamp 1667941163
transform 1 0 13340 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_140
timestamp 1667941163
transform 1 0 13984 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_148
timestamp 1667941163
transform 1 0 14720 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_154
timestamp 1667941163
transform 1 0 15272 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_160
timestamp 1667941163
transform 1 0 15824 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1667941163
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_173
timestamp 1667941163
transform 1 0 17020 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_177
timestamp 1667941163
transform 1 0 17388 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_184
timestamp 1667941163
transform 1 0 18032 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_190
timestamp 1667941163
transform 1 0 18584 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_196
timestamp 1667941163
transform 1 0 19136 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1667941163
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_231
timestamp 1667941163
transform 1 0 22356 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_252
timestamp 1667941163
transform 1 0 24288 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1667941163
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_285
timestamp 1667941163
transform 1 0 27324 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_291
timestamp 1667941163
transform 1 0 27876 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_297
timestamp 1667941163
transform 1 0 28428 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_324
timestamp 1667941163
transform 1 0 30912 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_330
timestamp 1667941163
transform 1 0 31464 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_341
timestamp 1667941163
transform 1 0 32476 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_345
timestamp 1667941163
transform 1 0 32844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_352
timestamp 1667941163
transform 1 0 33488 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_359
timestamp 1667941163
transform 1 0 34132 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_366
timestamp 1667941163
transform 1 0 34776 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_377
timestamp 1667941163
transform 1 0 35788 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_381
timestamp 1667941163
transform 1 0 36156 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_388
timestamp 1667941163
transform 1 0 36800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1667941163
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_60
timestamp 1667941163
transform 1 0 6624 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_66
timestamp 1667941163
transform 1 0 7176 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_78
timestamp 1667941163
transform 1 0 8280 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1667941163
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_156
timestamp 1667941163
transform 1 0 15456 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_163
timestamp 1667941163
transform 1 0 16100 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_170
timestamp 1667941163
transform 1 0 16744 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_183
timestamp 1667941163
transform 1 0 17940 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_190
timestamp 1667941163
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_202
timestamp 1667941163
transform 1 0 19688 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_208
timestamp 1667941163
transform 1 0 20240 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_232
timestamp 1667941163
transform 1 0 22448 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_238
timestamp 1667941163
transform 1 0 23000 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_244
timestamp 1667941163
transform 1 0 23552 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1667941163
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_277
timestamp 1667941163
transform 1 0 26588 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_304
timestamp 1667941163
transform 1 0 29072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_332
timestamp 1667941163
transform 1 0 31648 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_338
timestamp 1667941163
transform 1 0 32200 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_344
timestamp 1667941163
transform 1 0 32752 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_353
timestamp 1667941163
transform 1 0 33580 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_360
timestamp 1667941163
transform 1 0 34224 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_369
timestamp 1667941163
transform 1 0 35052 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_375
timestamp 1667941163
transform 1 0 35604 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_383
timestamp 1667941163
transform 1 0 36340 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_387
timestamp 1667941163
transform 1 0 36708 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_393
timestamp 1667941163
transform 1 0 37260 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_399
timestamp 1667941163
transform 1 0 37812 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_405
timestamp 1667941163
transform 1 0 38364 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_9
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_16
timestamp 1667941163
transform 1 0 2576 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_28
timestamp 1667941163
transform 1 0 3680 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_40
timestamp 1667941163
transform 1 0 4784 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1667941163
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_133
timestamp 1667941163
transform 1 0 13340 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_139
timestamp 1667941163
transform 1 0 13892 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_153
timestamp 1667941163
transform 1 0 15180 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1667941163
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_180
timestamp 1667941163
transform 1 0 17664 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_191
timestamp 1667941163
transform 1 0 18676 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_198
timestamp 1667941163
transform 1 0 19320 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1667941163
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_248
timestamp 1667941163
transform 1 0 23920 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_252
timestamp 1667941163
transform 1 0 24288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_274
timestamp 1667941163
transform 1 0 26312 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_304
timestamp 1667941163
transform 1 0 29072 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_310
timestamp 1667941163
transform 1 0 29624 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_316
timestamp 1667941163
transform 1 0 30176 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_322
timestamp 1667941163
transform 1 0 30728 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_328
timestamp 1667941163
transform 1 0 31280 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp 1667941163
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_341
timestamp 1667941163
transform 1 0 32476 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_347
timestamp 1667941163
transform 1 0 33028 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_353
timestamp 1667941163
transform 1 0 33580 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_359
timestamp 1667941163
transform 1 0 34132 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_365
timestamp 1667941163
transform 1 0 34684 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_371
timestamp 1667941163
transform 1 0 35236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_377
timestamp 1667941163
transform 1 0 35788 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_389
timestamp 1667941163
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_397
timestamp 1667941163
transform 1 0 37628 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_403
timestamp 1667941163
transform 1 0 38180 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1667941163
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1667941163
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1667941163
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1667941163
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_159
timestamp 1667941163
transform 1 0 15732 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_166
timestamp 1667941163
transform 1 0 16376 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_173
timestamp 1667941163
transform 1 0 17020 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_180
timestamp 1667941163
transform 1 0 17664 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_187
timestamp 1667941163
transform 1 0 18308 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1667941163
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_201
timestamp 1667941163
transform 1 0 19596 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_205
timestamp 1667941163
transform 1 0 19964 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_212
timestamp 1667941163
transform 1 0 20608 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_239
timestamp 1667941163
transform 1 0 23092 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_276
timestamp 1667941163
transform 1 0 26496 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_282
timestamp 1667941163
transform 1 0 27048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1667941163
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_313
timestamp 1667941163
transform 1 0 29900 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_319
timestamp 1667941163
transform 1 0 30452 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_325
timestamp 1667941163
transform 1 0 31004 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_331
timestamp 1667941163
transform 1 0 31556 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_337
timestamp 1667941163
transform 1 0 32108 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_343
timestamp 1667941163
transform 1 0 32660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_349
timestamp 1667941163
transform 1 0 33212 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_355
timestamp 1667941163
transform 1 0 33764 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_361
timestamp 1667941163
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_369
timestamp 1667941163
transform 1 0 35052 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_375
timestamp 1667941163
transform 1 0 35604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_381
timestamp 1667941163
transform 1 0 36156 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_387
timestamp 1667941163
transform 1 0 36708 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_393
timestamp 1667941163
transform 1 0 37260 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_399
timestamp 1667941163
transform 1 0 37812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1667941163
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_7
timestamp 1667941163
transform 1 0 1748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_19
timestamp 1667941163
transform 1 0 2852 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_31
timestamp 1667941163
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_43
timestamp 1667941163
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1667941163
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_133
timestamp 1667941163
transform 1 0 13340 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_137
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_150
timestamp 1667941163
transform 1 0 14904 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_163
timestamp 1667941163
transform 1 0 16100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1667941163
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_180
timestamp 1667941163
transform 1 0 17664 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1667941163
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_274
timestamp 1667941163
transform 1 0 26312 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_306
timestamp 1667941163
transform 1 0 29256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_330
timestamp 1667941163
transform 1 0 31464 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_341
timestamp 1667941163
transform 1 0 32476 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_347
timestamp 1667941163
transform 1 0 33028 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_353
timestamp 1667941163
transform 1 0 33580 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_359
timestamp 1667941163
transform 1 0 34132 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_365
timestamp 1667941163
transform 1 0 34684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_371
timestamp 1667941163
transform 1 0 35236 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_377
timestamp 1667941163
transform 1 0 35788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_383
timestamp 1667941163
transform 1 0 36340 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp 1667941163
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_398
timestamp 1667941163
transform 1 0 37720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_9
timestamp 1667941163
transform 1 0 1932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1667941163
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1667941163
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_146
timestamp 1667941163
transform 1 0 14536 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_153
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_166
timestamp 1667941163
transform 1 0 16376 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_170
timestamp 1667941163
transform 1 0 16744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_174
timestamp 1667941163
transform 1 0 17112 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_181
timestamp 1667941163
transform 1 0 17756 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1667941163
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_208
timestamp 1667941163
transform 1 0 20240 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_214
timestamp 1667941163
transform 1 0 20792 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_238
timestamp 1667941163
transform 1 0 23000 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_258
timestamp 1667941163
transform 1 0 24840 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_292
timestamp 1667941163
transform 1 0 27968 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_298
timestamp 1667941163
transform 1 0 28520 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1667941163
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_334
timestamp 1667941163
transform 1 0 31832 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_340
timestamp 1667941163
transform 1 0 32384 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_346
timestamp 1667941163
transform 1 0 32936 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_352
timestamp 1667941163
transform 1 0 33488 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_358
timestamp 1667941163
transform 1 0 34040 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_369
timestamp 1667941163
transform 1 0 35052 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_375
timestamp 1667941163
transform 1 0 35604 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_381
timestamp 1667941163
transform 1 0 36156 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_387
timestamp 1667941163
transform 1 0 36708 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_393
timestamp 1667941163
transform 1 0 37260 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_399
timestamp 1667941163
transform 1 0 37812 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1667941163
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1667941163
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_27
timestamp 1667941163
transform 1 0 3588 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_35
timestamp 1667941163
transform 1 0 4324 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_41
timestamp 1667941163
transform 1 0 4876 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_47
timestamp 1667941163
transform 1 0 5428 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1667941163
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_133
timestamp 1667941163
transform 1 0 13340 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_139
timestamp 1667941163
transform 1 0 13892 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_146
timestamp 1667941163
transform 1 0 14536 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_153
timestamp 1667941163
transform 1 0 15180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1667941163
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_180
timestamp 1667941163
transform 1 0 17664 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_188
timestamp 1667941163
transform 1 0 18400 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_198
timestamp 1667941163
transform 1 0 19320 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1667941163
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_250
timestamp 1667941163
transform 1 0 24104 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1667941163
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_306
timestamp 1667941163
transform 1 0 29256 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_312
timestamp 1667941163
transform 1 0 29808 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_318
timestamp 1667941163
transform 1 0 30360 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_324
timestamp 1667941163
transform 1 0 30912 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_330
timestamp 1667941163
transform 1 0 31464 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_341
timestamp 1667941163
transform 1 0 32476 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_347
timestamp 1667941163
transform 1 0 33028 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_353
timestamp 1667941163
transform 1 0 33580 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_359
timestamp 1667941163
transform 1 0 34132 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_365
timestamp 1667941163
transform 1 0 34684 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_371
timestamp 1667941163
transform 1 0 35236 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_377
timestamp 1667941163
transform 1 0 35788 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_383
timestamp 1667941163
transform 1 0 36340 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_389
timestamp 1667941163
transform 1 0 36892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_397
timestamp 1667941163
transform 1 0 37628 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1667941163
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1667941163
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1667941163
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1667941163
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_131
timestamp 1667941163
transform 1 0 13156 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1667941163
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1667941163
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1667941163
transform 1 0 14812 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_162
timestamp 1667941163
transform 1 0 16008 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_171
timestamp 1667941163
transform 1 0 16836 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_184
timestamp 1667941163
transform 1 0 18032 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_190
timestamp 1667941163
transform 1 0 18584 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1667941163
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_203
timestamp 1667941163
transform 1 0 19780 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_207
timestamp 1667941163
transform 1 0 20148 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_232
timestamp 1667941163
transform 1 0 22448 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1667941163
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1667941163
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_258
timestamp 1667941163
transform 1 0 24840 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_285
timestamp 1667941163
transform 1 0 27324 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_292
timestamp 1667941163
transform 1 0 27968 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_299
timestamp 1667941163
transform 1 0 28612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_305
timestamp 1667941163
transform 1 0 29164 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_313
timestamp 1667941163
transform 1 0 29900 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_319
timestamp 1667941163
transform 1 0 30452 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_325
timestamp 1667941163
transform 1 0 31004 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_331
timestamp 1667941163
transform 1 0 31556 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_338
timestamp 1667941163
transform 1 0 32200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_344
timestamp 1667941163
transform 1 0 32752 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_350
timestamp 1667941163
transform 1 0 33304 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_356
timestamp 1667941163
transform 1 0 33856 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_362
timestamp 1667941163
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_369
timestamp 1667941163
transform 1 0 35052 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_375
timestamp 1667941163
transform 1 0 35604 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_381
timestamp 1667941163
transform 1 0 36156 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_387
timestamp 1667941163
transform 1 0 36708 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_393
timestamp 1667941163
transform 1 0 37260 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_399
timestamp 1667941163
transform 1 0 37812 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_405
timestamp 1667941163
transform 1 0 38364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_9
timestamp 1667941163
transform 1 0 1932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_21
timestamp 1667941163
transform 1 0 3036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_33
timestamp 1667941163
transform 1 0 4140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp 1667941163
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1667941163
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1667941163
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_125
timestamp 1667941163
transform 1 0 12604 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_133
timestamp 1667941163
transform 1 0 13340 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_139
timestamp 1667941163
transform 1 0 13892 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_146
timestamp 1667941163
transform 1 0 14536 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_159
timestamp 1667941163
transform 1 0 15732 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1667941163
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_173
timestamp 1667941163
transform 1 0 17020 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_183
timestamp 1667941163
transform 1 0 17940 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1667941163
transform 1 0 19136 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1667941163
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1667941163
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_247
timestamp 1667941163
transform 1 0 23828 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_260
timestamp 1667941163
transform 1 0 25024 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1667941163
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1667941163
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_308
timestamp 1667941163
transform 1 0 29440 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_315
timestamp 1667941163
transform 1 0 30084 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_321
timestamp 1667941163
transform 1 0 30636 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_327
timestamp 1667941163
transform 1 0 31188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_333
timestamp 1667941163
transform 1 0 31740 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_341
timestamp 1667941163
transform 1 0 32476 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_352
timestamp 1667941163
transform 1 0 33488 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_358
timestamp 1667941163
transform 1 0 34040 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_364
timestamp 1667941163
transform 1 0 34592 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_367
timestamp 1667941163
transform 1 0 34868 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_371
timestamp 1667941163
transform 1 0 35236 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_374
timestamp 1667941163
transform 1 0 35512 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_384
timestamp 1667941163
transform 1 0 36432 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_390
timestamp 1667941163
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1667941163
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1667941163
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1667941163
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1667941163
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_109
timestamp 1667941163
transform 1 0 11132 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_115
timestamp 1667941163
transform 1 0 11684 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_118
timestamp 1667941163
transform 1 0 11960 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_125
timestamp 1667941163
transform 1 0 12604 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_131
timestamp 1667941163
transform 1 0 13156 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1667941163
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_146
timestamp 1667941163
transform 1 0 14536 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_159
timestamp 1667941163
transform 1 0 15732 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_174
timestamp 1667941163
transform 1 0 17112 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_181
timestamp 1667941163
transform 1 0 17756 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1667941163
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_203
timestamp 1667941163
transform 1 0 19780 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_217
timestamp 1667941163
transform 1 0 21068 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_230
timestamp 1667941163
transform 1 0 22264 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_243
timestamp 1667941163
transform 1 0 23460 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1667941163
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_264
timestamp 1667941163
transform 1 0 25392 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_277
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_285
timestamp 1667941163
transform 1 0 27324 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_293
timestamp 1667941163
transform 1 0 28060 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_300
timestamp 1667941163
transform 1 0 28704 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1667941163
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_314
timestamp 1667941163
transform 1 0 29992 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_327
timestamp 1667941163
transform 1 0 31188 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_339
timestamp 1667941163
transform 1 0 32292 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_370
timestamp 1667941163
transform 1 0 35144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_376
timestamp 1667941163
transform 1 0 35696 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_382
timestamp 1667941163
transform 1 0 36248 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_388
timestamp 1667941163
transform 1 0 36800 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_392
timestamp 1667941163
transform 1 0 37168 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_395
timestamp 1667941163
transform 1 0 37444 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_405
timestamp 1667941163
transform 1 0 38364 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_47
timestamp 1667941163
transform 1 0 5428 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1667941163
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_61
timestamp 1667941163
transform 1 0 6716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_73
timestamp 1667941163
transform 1 0 7820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_85
timestamp 1667941163
transform 1 0 8924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_97
timestamp 1667941163
transform 1 0 10028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 1667941163
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_123
timestamp 1667941163
transform 1 0 12420 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_129
timestamp 1667941163
transform 1 0 12972 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_136
timestamp 1667941163
transform 1 0 13616 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_142
timestamp 1667941163
transform 1 0 14168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_146
timestamp 1667941163
transform 1 0 14536 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_153
timestamp 1667941163
transform 1 0 15180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1667941163
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_173
timestamp 1667941163
transform 1 0 17020 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_183
timestamp 1667941163
transform 1 0 17940 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_187
timestamp 1667941163
transform 1 0 18308 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_197
timestamp 1667941163
transform 1 0 19228 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_206
timestamp 1667941163
transform 1 0 20056 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_219
timestamp 1667941163
transform 1 0 21252 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1667941163
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_235
timestamp 1667941163
transform 1 0 22724 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_248
timestamp 1667941163
transform 1 0 23920 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_261
timestamp 1667941163
transform 1 0 25116 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_267
timestamp 1667941163
transform 1 0 25668 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_277
timestamp 1667941163
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_292
timestamp 1667941163
transform 1 0 27968 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_299
timestamp 1667941163
transform 1 0 28612 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_306
timestamp 1667941163
transform 1 0 29256 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_313
timestamp 1667941163
transform 1 0 29900 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_320
timestamp 1667941163
transform 1 0 30544 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_327
timestamp 1667941163
transform 1 0 31188 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 1667941163
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_341
timestamp 1667941163
transform 1 0 32476 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_347
timestamp 1667941163
transform 1 0 33028 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_353
timestamp 1667941163
transform 1 0 33580 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_365
timestamp 1667941163
transform 1 0 34684 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_377
timestamp 1667941163
transform 1 0 35788 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1667941163
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_397
timestamp 1667941163
transform 1 0 37628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1667941163
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1667941163
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_117
timestamp 1667941163
transform 1 0 11868 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_120
timestamp 1667941163
transform 1 0 12144 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_126
timestamp 1667941163
transform 1 0 12696 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_132
timestamp 1667941163
transform 1 0 13248 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1667941163
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_148
timestamp 1667941163
transform 1 0 14720 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_155
timestamp 1667941163
transform 1 0 15364 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_162
timestamp 1667941163
transform 1 0 16008 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_175
timestamp 1667941163
transform 1 0 17204 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_183
timestamp 1667941163
transform 1 0 17940 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1667941163
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_212
timestamp 1667941163
transform 1 0 20608 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_216
timestamp 1667941163
transform 1 0 20976 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_230
timestamp 1667941163
transform 1 0 22264 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_234
timestamp 1667941163
transform 1 0 22632 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1667941163
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_264
timestamp 1667941163
transform 1 0 25392 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_268
timestamp 1667941163
transform 1 0 25760 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_278
timestamp 1667941163
transform 1 0 26680 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_291
timestamp 1667941163
transform 1 0 27876 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1667941163
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_314
timestamp 1667941163
transform 1 0 29992 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_328
timestamp 1667941163
transform 1 0 31280 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_335
timestamp 1667941163
transform 1 0 31924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_342
timestamp 1667941163
transform 1 0 32568 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_348
timestamp 1667941163
transform 1 0 33120 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_360
timestamp 1667941163
transform 1 0 34224 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_393
timestamp 1667941163
transform 1 0 37260 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_396
timestamp 1667941163
transform 1 0 37536 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_402
timestamp 1667941163
transform 1 0 38088 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_406
timestamp 1667941163
transform 1 0 38456 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_9
timestamp 1667941163
transform 1 0 1932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_21
timestamp 1667941163
transform 1 0 3036 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_33
timestamp 1667941163
transform 1 0 4140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1667941163
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1667941163
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_125
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_128
timestamp 1667941163
transform 1 0 12880 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_134
timestamp 1667941163
transform 1 0 13432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_140
timestamp 1667941163
transform 1 0 13984 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_146
timestamp 1667941163
transform 1 0 14536 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp 1667941163
transform 1 0 15180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1667941163
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_173
timestamp 1667941163
transform 1 0 17020 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_177
timestamp 1667941163
transform 1 0 17388 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_190
timestamp 1667941163
transform 1 0 18584 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_207
timestamp 1667941163
transform 1 0 20148 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1667941163
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_240
timestamp 1667941163
transform 1 0 23184 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_253
timestamp 1667941163
transform 1 0 24380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_260
timestamp 1667941163
transform 1 0 25024 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1667941163
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1667941163
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_287
timestamp 1667941163
transform 1 0 27508 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_297
timestamp 1667941163
transform 1 0 28428 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_304
timestamp 1667941163
transform 1 0 29072 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_311
timestamp 1667941163
transform 1 0 29716 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_318
timestamp 1667941163
transform 1 0 30360 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_325
timestamp 1667941163
transform 1 0 31004 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_332
timestamp 1667941163
transform 1 0 31648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_342
timestamp 1667941163
transform 1 0 32568 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_348
timestamp 1667941163
transform 1 0 33120 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_360
timestamp 1667941163
transform 1 0 34224 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_372
timestamp 1667941163
transform 1 0 35328 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_384
timestamp 1667941163
transform 1 0 36432 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_399
timestamp 1667941163
transform 1 0 37812 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_402
timestamp 1667941163
transform 1 0 38088 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_406
timestamp 1667941163
transform 1 0 38456 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1667941163
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1667941163
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1667941163
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_121
timestamp 1667941163
transform 1 0 12236 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_126
timestamp 1667941163
transform 1 0 12696 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_132
timestamp 1667941163
transform 1 0 13248 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1667941163
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_149
timestamp 1667941163
transform 1 0 14812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_156
timestamp 1667941163
transform 1 0 15456 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1667941163
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_170
timestamp 1667941163
transform 1 0 16744 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_178
timestamp 1667941163
transform 1 0 17480 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_191
timestamp 1667941163
transform 1 0 18676 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1667941163
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_208
timestamp 1667941163
transform 1 0 20240 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_212
timestamp 1667941163
transform 1 0 20608 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_222
timestamp 1667941163
transform 1 0 21528 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_243
timestamp 1667941163
transform 1 0 23460 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1667941163
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_270
timestamp 1667941163
transform 1 0 25944 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_289
timestamp 1667941163
transform 1 0 27692 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1667941163
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_320
timestamp 1667941163
transform 1 0 30544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_327
timestamp 1667941163
transform 1 0 31188 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_334
timestamp 1667941163
transform 1 0 31832 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_341
timestamp 1667941163
transform 1 0 32476 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_348
timestamp 1667941163
transform 1 0 33120 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_360
timestamp 1667941163
transform 1 0 34224 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_7
timestamp 1667941163
transform 1 0 1748 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_19
timestamp 1667941163
transform 1 0 2852 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_31
timestamp 1667941163
transform 1 0 3956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_43
timestamp 1667941163
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1667941163
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1667941163
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1667941163
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_125
timestamp 1667941163
transform 1 0 12604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_135
timestamp 1667941163
transform 1 0 13524 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_141
timestamp 1667941163
transform 1 0 14076 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_147
timestamp 1667941163
transform 1 0 14628 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1667941163
transform 1 0 15180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_159
timestamp 1667941163
transform 1 0 15732 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1667941163
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_174
timestamp 1667941163
transform 1 0 17112 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_181
timestamp 1667941163
transform 1 0 17756 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_194
timestamp 1667941163
transform 1 0 18952 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_198
timestamp 1667941163
transform 1 0 19320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_202
timestamp 1667941163
transform 1 0 19688 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_209
timestamp 1667941163
transform 1 0 20332 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1667941163
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_230
timestamp 1667941163
transform 1 0 22264 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_237
timestamp 1667941163
transform 1 0 22908 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_250
timestamp 1667941163
transform 1 0 24104 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_263
timestamp 1667941163
transform 1 0 25300 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_275
timestamp 1667941163
transform 1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1667941163
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_291
timestamp 1667941163
transform 1 0 27876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_304
timestamp 1667941163
transform 1 0 29072 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_311
timestamp 1667941163
transform 1 0 29716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_318
timestamp 1667941163
transform 1 0 30360 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_324
timestamp 1667941163
transform 1 0 30912 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1667941163
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_342
timestamp 1667941163
transform 1 0 32568 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_348
timestamp 1667941163
transform 1 0 33120 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_360
timestamp 1667941163
transform 1 0 34224 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_372
timestamp 1667941163
transform 1 0 35328 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_384
timestamp 1667941163
transform 1 0 36432 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_397
timestamp 1667941163
transform 1 0 37628 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1667941163
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1667941163
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_90
timestamp 1667941163
transform 1 0 9384 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_102
timestamp 1667941163
transform 1 0 10488 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_114
timestamp 1667941163
transform 1 0 11592 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_126
timestamp 1667941163
transform 1 0 12696 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_134
timestamp 1667941163
transform 1 0 13432 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1667941163
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_147
timestamp 1667941163
transform 1 0 14628 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_153
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_166
timestamp 1667941163
transform 1 0 16376 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_170
timestamp 1667941163
transform 1 0 16744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_174
timestamp 1667941163
transform 1 0 17112 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_181
timestamp 1667941163
transform 1 0 17756 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1667941163
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_202
timestamp 1667941163
transform 1 0 19688 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_209
timestamp 1667941163
transform 1 0 20332 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_224
timestamp 1667941163
transform 1 0 21712 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_231
timestamp 1667941163
transform 1 0 22356 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_247
timestamp 1667941163
transform 1 0 23828 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1667941163
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_264
timestamp 1667941163
transform 1 0 25392 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_270
timestamp 1667941163
transform 1 0 25944 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_287
timestamp 1667941163
transform 1 0 27508 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_299
timestamp 1667941163
transform 1 0 28612 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1667941163
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_314
timestamp 1667941163
transform 1 0 29992 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_328
timestamp 1667941163
transform 1 0 31280 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_335
timestamp 1667941163
transform 1 0 31924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_341
timestamp 1667941163
transform 1 0 32476 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_347
timestamp 1667941163
transform 1 0 33028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_359
timestamp 1667941163
transform 1 0 34132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_401
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1667941163
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1667941163
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1667941163
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_137
timestamp 1667941163
transform 1 0 13708 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_145
timestamp 1667941163
transform 1 0 14444 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_149
timestamp 1667941163
transform 1 0 14812 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_159
timestamp 1667941163
transform 1 0 15732 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1667941163
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_182
timestamp 1667941163
transform 1 0 17848 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_193
timestamp 1667941163
transform 1 0 18860 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_210
timestamp 1667941163
transform 1 0 20424 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_216
timestamp 1667941163
transform 1 0 20976 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1667941163
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_232
timestamp 1667941163
transform 1 0 22448 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_245
timestamp 1667941163
transform 1 0 23644 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_258
timestamp 1667941163
transform 1 0 24840 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_270
timestamp 1667941163
transform 1 0 25944 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1667941163
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_294
timestamp 1667941163
transform 1 0 28152 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_306
timestamp 1667941163
transform 1 0 29256 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_318
timestamp 1667941163
transform 1 0 30360 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_325
timestamp 1667941163
transform 1 0 31004 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_332
timestamp 1667941163
transform 1 0 31648 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1667941163
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1667941163
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1667941163
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1667941163
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1667941163
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1667941163
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1667941163
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_153
timestamp 1667941163
transform 1 0 15180 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_158
timestamp 1667941163
transform 1 0 15640 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_166
timestamp 1667941163
transform 1 0 16376 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_170
timestamp 1667941163
transform 1 0 16744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_180
timestamp 1667941163
transform 1 0 17664 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1667941163
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_208
timestamp 1667941163
transform 1 0 20240 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1667941163
transform 1 0 20884 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_222
timestamp 1667941163
transform 1 0 21528 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_228
timestamp 1667941163
transform 1 0 22080 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_232
timestamp 1667941163
transform 1 0 22448 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_244
timestamp 1667941163
transform 1 0 23552 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1667941163
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_257
timestamp 1667941163
transform 1 0 24748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_270
timestamp 1667941163
transform 1 0 25944 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_282
timestamp 1667941163
transform 1 0 27048 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_295
timestamp 1667941163
transform 1 0 28244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_302
timestamp 1667941163
transform 1 0 28888 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_314
timestamp 1667941163
transform 1 0 29992 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_330
timestamp 1667941163
transform 1 0 31464 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_342
timestamp 1667941163
transform 1 0 32568 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_350
timestamp 1667941163
transform 1 0 33304 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_355
timestamp 1667941163
transform 1 0 33764 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1667941163
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_397
timestamp 1667941163
transform 1 0 37628 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_402
timestamp 1667941163
transform 1 0 38088 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_406
timestamp 1667941163
transform 1 0 38456 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1667941163
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1667941163
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1667941163
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1667941163
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1667941163
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1667941163
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1667941163
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1667941163
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1667941163
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_149
timestamp 1667941163
transform 1 0 14812 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_154
timestamp 1667941163
transform 1 0 15272 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_162
timestamp 1667941163
transform 1 0 16008 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1667941163
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_180
timestamp 1667941163
transform 1 0 17664 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_184
timestamp 1667941163
transform 1 0 18032 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_194
timestamp 1667941163
transform 1 0 18952 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_201
timestamp 1667941163
transform 1 0 19596 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_207
timestamp 1667941163
transform 1 0 20148 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_211
timestamp 1667941163
transform 1 0 20516 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_218
timestamp 1667941163
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_231
timestamp 1667941163
transform 1 0 22356 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_241
timestamp 1667941163
transform 1 0 23276 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_254
timestamp 1667941163
transform 1 0 24472 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_267
timestamp 1667941163
transform 1 0 25668 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_274
timestamp 1667941163
transform 1 0 26312 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_292
timestamp 1667941163
transform 1 0 27968 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_299
timestamp 1667941163
transform 1 0 28612 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_306
timestamp 1667941163
transform 1 0 29256 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_313
timestamp 1667941163
transform 1 0 29900 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_320
timestamp 1667941163
transform 1 0 30544 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_332
timestamp 1667941163
transform 1 0 31648 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1667941163
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1667941163
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1667941163
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1667941163
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1667941163
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_165
timestamp 1667941163
transform 1 0 16284 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_175
timestamp 1667941163
transform 1 0 17204 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_181
timestamp 1667941163
transform 1 0 17756 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_187
timestamp 1667941163
transform 1 0 18308 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1667941163
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_208
timestamp 1667941163
transform 1 0 20240 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_214
timestamp 1667941163
transform 1 0 20792 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_218
timestamp 1667941163
transform 1 0 21160 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_224
timestamp 1667941163
transform 1 0 21712 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_232
timestamp 1667941163
transform 1 0 22448 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_238
timestamp 1667941163
transform 1 0 23000 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1667941163
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_264
timestamp 1667941163
transform 1 0 25392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_281
timestamp 1667941163
transform 1 0 26956 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_293
timestamp 1667941163
transform 1 0 28060 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_300
timestamp 1667941163
transform 1 0 28704 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_306
timestamp 1667941163
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_313
timestamp 1667941163
transform 1 0 29900 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_319
timestamp 1667941163
transform 1 0 30452 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_331
timestamp 1667941163
transform 1 0 31556 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_343
timestamp 1667941163
transform 1 0 32660 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_355
timestamp 1667941163
transform 1 0 33764 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_401
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_405
timestamp 1667941163
transform 1 0 38364 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1667941163
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1667941163
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1667941163
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1667941163
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1667941163
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1667941163
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1667941163
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1667941163
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_161
timestamp 1667941163
transform 1 0 15916 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1667941163
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_174
timestamp 1667941163
transform 1 0 17112 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_180
timestamp 1667941163
transform 1 0 17664 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_183
timestamp 1667941163
transform 1 0 17940 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_189
timestamp 1667941163
transform 1 0 18492 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_195
timestamp 1667941163
transform 1 0 19044 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_201
timestamp 1667941163
transform 1 0 19596 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_208
timestamp 1667941163
transform 1 0 20240 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1667941163
transform 1 0 20884 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1667941163
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_236
timestamp 1667941163
transform 1 0 22816 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_243
timestamp 1667941163
transform 1 0 23460 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_251
timestamp 1667941163
transform 1 0 24196 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_261
timestamp 1667941163
transform 1 0 25116 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_267
timestamp 1667941163
transform 1 0 25668 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 1667941163
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_286
timestamp 1667941163
transform 1 0 27416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_300
timestamp 1667941163
transform 1 0 28704 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_306
timestamp 1667941163
transform 1 0 29256 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_312
timestamp 1667941163
transform 1 0 29808 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_324
timestamp 1667941163
transform 1 0 30912 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1667941163
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1667941163
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1667941163
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1667941163
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1667941163
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1667941163
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1667941163
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_165
timestamp 1667941163
transform 1 0 16284 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_176
timestamp 1667941163
transform 1 0 17296 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_182
timestamp 1667941163
transform 1 0 17848 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_188
timestamp 1667941163
transform 1 0 18400 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1667941163
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_202
timestamp 1667941163
transform 1 0 19688 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1667941163
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_222
timestamp 1667941163
transform 1 0 21528 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_230
timestamp 1667941163
transform 1 0 22264 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_234
timestamp 1667941163
transform 1 0 22632 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1667941163
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_257
timestamp 1667941163
transform 1 0 24748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_267
timestamp 1667941163
transform 1 0 25668 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_274
timestamp 1667941163
transform 1 0 26312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_281
timestamp 1667941163
transform 1 0 26956 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_288
timestamp 1667941163
transform 1 0 27600 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_295
timestamp 1667941163
transform 1 0 28244 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_302
timestamp 1667941163
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_313
timestamp 1667941163
transform 1 0 29900 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_325
timestamp 1667941163
transform 1 0 31004 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_337
timestamp 1667941163
transform 1 0 32108 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_349
timestamp 1667941163
transform 1 0 33212 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_361
timestamp 1667941163
transform 1 0 34316 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_9
timestamp 1667941163
transform 1 0 1932 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_21
timestamp 1667941163
transform 1 0 3036 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_33
timestamp 1667941163
transform 1 0 4140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_45
timestamp 1667941163
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1667941163
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1667941163
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1667941163
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1667941163
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1667941163
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1667941163
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1667941163
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_186
timestamp 1667941163
transform 1 0 18216 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_190
timestamp 1667941163
transform 1 0 18584 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_194
timestamp 1667941163
transform 1 0 18952 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_200
timestamp 1667941163
transform 1 0 19504 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_206
timestamp 1667941163
transform 1 0 20056 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_213
timestamp 1667941163
transform 1 0 20700 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1667941163
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_236
timestamp 1667941163
transform 1 0 22816 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_249
timestamp 1667941163
transform 1 0 24012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_257
timestamp 1667941163
transform 1 0 24748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_265
timestamp 1667941163
transform 1 0 25484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_269
timestamp 1667941163
transform 1 0 25852 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1667941163
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_286
timestamp 1667941163
transform 1 0 27416 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_292
timestamp 1667941163
transform 1 0 27968 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_298
timestamp 1667941163
transform 1 0 28520 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_304
timestamp 1667941163
transform 1 0 29072 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_310
timestamp 1667941163
transform 1 0 29624 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_322
timestamp 1667941163
transform 1 0 30728 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1667941163
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1667941163
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1667941163
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1667941163
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1667941163
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_101
timestamp 1667941163
transform 1 0 10396 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_107
timestamp 1667941163
transform 1 0 10948 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_119
timestamp 1667941163
transform 1 0 12052 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_131
timestamp 1667941163
transform 1 0 13156 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1667941163
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1667941163
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1667941163
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_177
timestamp 1667941163
transform 1 0 17388 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_182
timestamp 1667941163
transform 1 0 17848 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1667941163
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_201
timestamp 1667941163
transform 1 0 19596 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_204
timestamp 1667941163
transform 1 0 19872 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1667941163
transform 1 0 20424 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_217
timestamp 1667941163
transform 1 0 21068 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_229
timestamp 1667941163
transform 1 0 22172 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_242
timestamp 1667941163
transform 1 0 23368 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 1667941163
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_264
timestamp 1667941163
transform 1 0 25392 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_271
timestamp 1667941163
transform 1 0 26036 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_278
timestamp 1667941163
transform 1 0 26680 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_285
timestamp 1667941163
transform 1 0 27324 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_291
timestamp 1667941163
transform 1 0 27876 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_297
timestamp 1667941163
transform 1 0 28428 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_303
timestamp 1667941163
transform 1 0 28980 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1667941163
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1667941163
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_7
timestamp 1667941163
transform 1 0 1748 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_19
timestamp 1667941163
transform 1 0 2852 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_31
timestamp 1667941163
transform 1 0 3956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_43
timestamp 1667941163
transform 1 0 5060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1667941163
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_92
timestamp 1667941163
transform 1 0 9568 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_104
timestamp 1667941163
transform 1 0 10672 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1667941163
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1667941163
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1667941163
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1667941163
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1667941163
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1667941163
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1667941163
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_205
timestamp 1667941163
transform 1 0 19964 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1667941163
transform 1 0 20884 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1667941163
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_235
timestamp 1667941163
transform 1 0 22724 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_252
timestamp 1667941163
transform 1 0 24288 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_264
timestamp 1667941163
transform 1 0 25392 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_271
timestamp 1667941163
transform 1 0 26036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1667941163
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_285
timestamp 1667941163
transform 1 0 27324 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_291
timestamp 1667941163
transform 1 0 27876 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_303
timestamp 1667941163
transform 1 0 28980 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_315
timestamp 1667941163
transform 1 0 30084 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_327
timestamp 1667941163
transform 1 0 31188 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1667941163
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_9
timestamp 1667941163
transform 1 0 1932 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1667941163
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1667941163
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1667941163
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1667941163
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1667941163
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1667941163
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1667941163
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1667941163
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1667941163
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1667941163
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1667941163
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1667941163
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1667941163
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_221
timestamp 1667941163
transform 1 0 21436 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_224
timestamp 1667941163
transform 1 0 21712 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_231
timestamp 1667941163
transform 1 0 22356 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_247
timestamp 1667941163
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_266
timestamp 1667941163
transform 1 0 25576 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_273
timestamp 1667941163
transform 1 0 26220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_280
timestamp 1667941163
transform 1 0 26864 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_292
timestamp 1667941163
transform 1 0 27968 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_304
timestamp 1667941163
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1667941163
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1667941163
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1667941163
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1667941163
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1667941163
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1667941163
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1667941163
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1667941163
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1667941163
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1667941163
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1667941163
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1667941163
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1667941163
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1667941163
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1667941163
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1667941163
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_229
timestamp 1667941163
transform 1 0 22172 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_233
timestamp 1667941163
transform 1 0 22540 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_240
timestamp 1667941163
transform 1 0 23184 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_246
timestamp 1667941163
transform 1 0 23736 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_258
timestamp 1667941163
transform 1 0 24840 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_265
timestamp 1667941163
transform 1 0 25484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 1667941163
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1667941163
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_10
timestamp 1667941163
transform 1 0 2024 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_22
timestamp 1667941163
transform 1 0 3128 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1667941163
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1667941163
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1667941163
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1667941163
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1667941163
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1667941163
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1667941163
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1667941163
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1667941163
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1667941163
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1667941163
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1667941163
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_221
timestamp 1667941163
transform 1 0 21436 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_227
timestamp 1667941163
transform 1 0 21988 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_230
timestamp 1667941163
transform 1 0 22264 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_242
timestamp 1667941163
transform 1 0 23368 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1667941163
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_258
timestamp 1667941163
transform 1 0 24840 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_270
timestamp 1667941163
transform 1 0 25944 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_282
timestamp 1667941163
transform 1 0 27048 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_294
timestamp 1667941163
transform 1 0 28152 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_306
timestamp 1667941163
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_9
timestamp 1667941163
transform 1 0 1932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_21
timestamp 1667941163
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_33
timestamp 1667941163
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_45
timestamp 1667941163
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1667941163
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_66
timestamp 1667941163
transform 1 0 7176 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_72
timestamp 1667941163
transform 1 0 7728 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_84
timestamp 1667941163
transform 1 0 8832 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_96
timestamp 1667941163
transform 1 0 9936 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1667941163
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1667941163
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1667941163
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1667941163
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1667941163
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1667941163
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1667941163
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1667941163
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1667941163
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1667941163
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_249
timestamp 1667941163
transform 1 0 24012 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_257
timestamp 1667941163
transform 1 0 24748 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_261
timestamp 1667941163
transform 1 0 25116 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_269
timestamp 1667941163
transform 1 0 25852 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_277
timestamp 1667941163
transform 1 0 26588 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1667941163
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_341
timestamp 1667941163
transform 1 0 32476 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_345
timestamp 1667941163
transform 1 0 32844 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_351
timestamp 1667941163
transform 1 0 33396 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_363
timestamp 1667941163
transform 1 0 34500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_375
timestamp 1667941163
transform 1 0 35604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_387
timestamp 1667941163
transform 1 0 36708 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1667941163
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1667941163
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1667941163
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1667941163
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1667941163
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1667941163
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1667941163
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1667941163
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1667941163
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1667941163
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1667941163
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1667941163
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1667941163
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_233
timestamp 1667941163
transform 1 0 22540 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_239
timestamp 1667941163
transform 1 0 23092 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1667941163
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1667941163
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1667941163
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_401
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1667941163
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1667941163
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1667941163
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1667941163
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1667941163
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1667941163
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1667941163
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1667941163
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1667941163
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1667941163
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1667941163
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1667941163
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1667941163
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1667941163
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1667941163
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1667941163
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1667941163
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1667941163
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1667941163
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1667941163
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1667941163
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1667941163
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_7
timestamp 1667941163
transform 1 0 1748 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_19
timestamp 1667941163
transform 1 0 2852 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1667941163
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1667941163
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1667941163
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1667941163
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1667941163
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1667941163
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1667941163
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1667941163
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1667941163
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1667941163
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1667941163
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_233
timestamp 1667941163
transform 1 0 22540 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_239
timestamp 1667941163
transform 1 0 23092 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_243
timestamp 1667941163
transform 1 0 23460 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_249
timestamp 1667941163
transform 1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1667941163
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1667941163
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1667941163
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1667941163
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1667941163
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1667941163
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1667941163
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1667941163
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1667941163
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1667941163
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1667941163
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1667941163
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1667941163
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1667941163
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1667941163
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1667941163
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1667941163
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1667941163
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1667941163
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1667941163
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1667941163
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1667941163
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1667941163
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1667941163
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1667941163
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1667941163
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1667941163
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1667941163
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1667941163
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1667941163
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1667941163
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1667941163
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1667941163
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1667941163
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1667941163
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1667941163
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1667941163
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1667941163
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1667941163
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1667941163
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_401
timestamp 1667941163
transform 1 0 37996 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1667941163
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_7
timestamp 1667941163
transform 1 0 1748 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_19
timestamp 1667941163
transform 1 0 2852 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_31
timestamp 1667941163
transform 1 0 3956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_43
timestamp 1667941163
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1667941163
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1667941163
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1667941163
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1667941163
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1667941163
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1667941163
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1667941163
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1667941163
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1667941163
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1667941163
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1667941163
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1667941163
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1667941163
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1667941163
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1667941163
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1667941163
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1667941163
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1667941163
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_69
timestamp 1667941163
transform 1 0 7452 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_75
timestamp 1667941163
transform 1 0 8004 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_90
timestamp 1667941163
transform 1 0 9384 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_96
timestamp 1667941163
transform 1 0 9936 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_108
timestamp 1667941163
transform 1 0 11040 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_120
timestamp 1667941163
transform 1 0 12144 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_132
timestamp 1667941163
transform 1 0 13248 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1667941163
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1667941163
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1667941163
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1667941163
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1667941163
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1667941163
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1667941163
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1667941163
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1667941163
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1667941163
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1667941163
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1667941163
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1667941163
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1667941163
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1667941163
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_401
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1667941163
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1667941163
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1667941163
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1667941163
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1667941163
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1667941163
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1667941163
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1667941163
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1667941163
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1667941163
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1667941163
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1667941163
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1667941163
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1667941163
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1667941163
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1667941163
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1667941163
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1667941163
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1667941163
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1667941163
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1667941163
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1667941163
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1667941163
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1667941163
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1667941163
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1667941163
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1667941163
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1667941163
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1667941163
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1667941163
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1667941163
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_401
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_405
timestamp 1667941163
transform 1 0 38364 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_9
timestamp 1667941163
transform 1 0 1932 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_21
timestamp 1667941163
transform 1 0 3036 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_33
timestamp 1667941163
transform 1 0 4140 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_45
timestamp 1667941163
transform 1 0 5244 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1667941163
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1667941163
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1667941163
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1667941163
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1667941163
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1667941163
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1667941163
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1667941163
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1667941163
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1667941163
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1667941163
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1667941163
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1667941163
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1667941163
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1667941163
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1667941163
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1667941163
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_152
timestamp 1667941163
transform 1 0 15088 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_164
timestamp 1667941163
transform 1 0 16192 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_176
timestamp 1667941163
transform 1 0 17296 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_188
timestamp 1667941163
transform 1 0 18400 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1667941163
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1667941163
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1667941163
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1667941163
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_337
timestamp 1667941163
transform 1 0 32108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_341
timestamp 1667941163
transform 1 0 32476 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_353
timestamp 1667941163
transform 1 0 33580 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_361
timestamp 1667941163
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1667941163
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1667941163
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1667941163
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1667941163
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1667941163
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1667941163
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1667941163
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1667941163
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1667941163
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_181
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_47_190
timestamp 1667941163
transform 1 0 18584 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_199
timestamp 1667941163
transform 1 0 19412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_211
timestamp 1667941163
transform 1 0 20516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1667941163
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_230
timestamp 1667941163
transform 1 0 22264 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_242
timestamp 1667941163
transform 1 0 23368 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_254
timestamp 1667941163
transform 1 0 24472 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_268
timestamp 1667941163
transform 1 0 25760 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_275
timestamp 1667941163
transform 1 0 26404 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1667941163
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_299
timestamp 1667941163
transform 1 0 28612 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_311
timestamp 1667941163
transform 1 0 29716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_323
timestamp 1667941163
transform 1 0 30820 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_397
timestamp 1667941163
transform 1 0 37628 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_7
timestamp 1667941163
transform 1 0 1748 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_19
timestamp 1667941163
transform 1 0 2852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1667941163
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1667941163
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_160
timestamp 1667941163
transform 1 0 15824 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_172
timestamp 1667941163
transform 1 0 16928 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_184
timestamp 1667941163
transform 1 0 18032 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_203
timestamp 1667941163
transform 1 0 19780 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_207
timestamp 1667941163
transform 1 0 20148 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_213
timestamp 1667941163
transform 1 0 20700 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_225
timestamp 1667941163
transform 1 0 21804 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_237
timestamp 1667941163
transform 1 0 22908 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_249
timestamp 1667941163
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1667941163
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1667941163
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_9
timestamp 1667941163
transform 1 0 1932 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_21
timestamp 1667941163
transform 1 0 3036 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_33
timestamp 1667941163
transform 1 0 4140 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_45
timestamp 1667941163
transform 1 0 5244 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1667941163
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1667941163
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1667941163
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1667941163
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1667941163
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1667941163
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1667941163
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1667941163
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1667941163
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1667941163
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1667941163
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1667941163
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_233
timestamp 1667941163
transform 1 0 22540 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_241
timestamp 1667941163
transform 1 0 23276 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_247
timestamp 1667941163
transform 1 0 23828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1667941163
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1667941163
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1667941163
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_401
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_7
timestamp 1667941163
transform 1 0 1748 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_19
timestamp 1667941163
transform 1 0 2852 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_31
timestamp 1667941163
transform 1 0 3956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_43
timestamp 1667941163
transform 1 0 5060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1667941163
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1667941163
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1667941163
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1667941163
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1667941163
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1667941163
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1667941163
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1667941163
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1667941163
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1667941163
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1667941163
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1667941163
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_313
timestamp 1667941163
transform 1 0 29900 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_319
timestamp 1667941163
transform 1 0 30452 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_325
timestamp 1667941163
transform 1 0 31004 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_333
timestamp 1667941163
transform 1 0 31740 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_397
timestamp 1667941163
transform 1 0 37628 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_9
timestamp 1667941163
transform 1 0 1932 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_16
timestamp 1667941163
transform 1 0 2576 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_22
timestamp 1667941163
transform 1 0 3128 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1667941163
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1667941163
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1667941163
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1667941163
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1667941163
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1667941163
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1667941163
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1667941163
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_286
timestamp 1667941163
transform 1 0 27416 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_292
timestamp 1667941163
transform 1 0 27968 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1667941163
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1667941163
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1667941163
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1667941163
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1667941163
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1667941163
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1667941163
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1667941163
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1667941163
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1667941163
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1667941163
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1667941163
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1667941163
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_405
timestamp 1667941163
transform 1 0 38364 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_9
timestamp 1667941163
transform 1 0 1932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_21
timestamp 1667941163
transform 1 0 3036 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_33
timestamp 1667941163
transform 1 0 4140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1667941163
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1667941163
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_286
timestamp 1667941163
transform 1 0 27416 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_292
timestamp 1667941163
transform 1 0 27968 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_304
timestamp 1667941163
transform 1 0 29072 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_316
timestamp 1667941163
transform 1 0 30176 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_328
timestamp 1667941163
transform 1 0 31280 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1667941163
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1667941163
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1667941163
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1667941163
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1667941163
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_397
timestamp 1667941163
transform 1 0 37628 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_9
timestamp 1667941163
transform 1 0 1932 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_16
timestamp 1667941163
transform 1 0 2576 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_22
timestamp 1667941163
transform 1 0 3128 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_34
timestamp 1667941163
transform 1 0 4232 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_46
timestamp 1667941163
transform 1 0 5336 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_54
timestamp 1667941163
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_401
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_405
timestamp 1667941163
transform 1 0 38364 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1667941163
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1667941163
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1667941163
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1667941163
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_310
timestamp 1667941163
transform 1 0 29624 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_322
timestamp 1667941163
transform 1 0 30728 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_334
timestamp 1667941163
transform 1 0 31832 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_9
timestamp 1667941163
transform 1 0 1932 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_21
timestamp 1667941163
transform 1 0 3036 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1667941163
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_115
timestamp 1667941163
transform 1 0 11684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_127
timestamp 1667941163
transform 1 0 12788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_393
timestamp 1667941163
transform 1 0 37260 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_397
timestamp 1667941163
transform 1 0 37628 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_17
timestamp 1667941163
transform 1 0 2668 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_23
timestamp 1667941163
transform 1 0 3220 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_35
timestamp 1667941163
transform 1 0 4324 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_47
timestamp 1667941163
transform 1 0 5428 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1667941163
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_62
timestamp 1667941163
transform 1 0 6808 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_74
timestamp 1667941163
transform 1 0 7912 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_86
timestamp 1667941163
transform 1 0 9016 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_98
timestamp 1667941163
transform 1 0 10120 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1667941163
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1667941163
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1667941163
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1667941163
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1667941163
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1667941163
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1667941163
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1667941163
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_241
timestamp 1667941163
transform 1 0 23276 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_253
timestamp 1667941163
transform 1 0 24380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_265
timestamp 1667941163
transform 1 0 25484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_277
timestamp 1667941163
transform 1 0 26588 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_286
timestamp 1667941163
transform 1 0 27416 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_298
timestamp 1667941163
transform 1 0 28520 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_310
timestamp 1667941163
transform 1 0 29624 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_322
timestamp 1667941163
transform 1 0 30728 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_334
timestamp 1667941163
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_370
timestamp 1667941163
transform 1 0 35144 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_376
timestamp 1667941163
transform 1 0 35696 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_63_386
timestamp 1667941163
transform 1 0 36616 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_9
timestamp 1667941163
transform 1 0 1932 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_21
timestamp 1667941163
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1667941163
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_33
timestamp 1667941163
transform 1 0 4140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_37
timestamp 1667941163
transform 1 0 4508 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_42
timestamp 1667941163
transform 1 0 4968 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_48
timestamp 1667941163
transform 1 0 5520 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_54
timestamp 1667941163
transform 1 0 6072 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_63
timestamp 1667941163
transform 1 0 6900 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_71
timestamp 1667941163
transform 1 0 7636 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1667941163
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1667941163
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_90
timestamp 1667941163
transform 1 0 9384 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_98
timestamp 1667941163
transform 1 0 10120 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_110
timestamp 1667941163
transform 1 0 11224 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_125
timestamp 1667941163
transform 1 0 12604 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1667941163
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_145
timestamp 1667941163
transform 1 0 14444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_149
timestamp 1667941163
transform 1 0 14812 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_154
timestamp 1667941163
transform 1 0 15272 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_166
timestamp 1667941163
transform 1 0 16376 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_175
timestamp 1667941163
transform 1 0 17204 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_183
timestamp 1667941163
transform 1 0 17940 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1667941163
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1667941163
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_205
timestamp 1667941163
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_210
timestamp 1667941163
transform 1 0 20424 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_216
timestamp 1667941163
transform 1 0 20976 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1667941163
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_237
timestamp 1667941163
transform 1 0 22908 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1667941163
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1667941163
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_258
timestamp 1667941163
transform 1 0 24840 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_266
timestamp 1667941163
transform 1 0 25576 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_274
timestamp 1667941163
transform 1 0 26312 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_278
timestamp 1667941163
transform 1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_287
timestamp 1667941163
transform 1 0 27508 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_295
timestamp 1667941163
transform 1 0 28244 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1667941163
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1667941163
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_317
timestamp 1667941163
transform 1 0 30268 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_322
timestamp 1667941163
transform 1 0 30728 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_334
timestamp 1667941163
transform 1 0 31832 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_343
timestamp 1667941163
transform 1 0 32660 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_351
timestamp 1667941163
transform 1 0 33396 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1667941163
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1667941163
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_370
timestamp 1667941163
transform 1 0 35144 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_378
timestamp 1667941163
transform 1 0 35880 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_390
timestamp 1667941163
transform 1 0 36984 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_399
timestamp 1667941163
transform 1 0 37812 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _213_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 17480 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _214_
timestamp 1667941163
transform 1 0 23368 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _215_
timestamp 1667941163
transform 1 0 14904 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _216_
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1667941163
transform -1 0 17112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1667941163
transform -1 0 16836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1667941163
transform 1 0 30360 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1667941163
transform 1 0 14904 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _221_
timestamp 1667941163
transform -1 0 17664 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1667941163
transform -1 0 18308 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _223_
timestamp 1667941163
transform 1 0 20608 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _224_
timestamp 1667941163
transform 1 0 16836 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1667941163
transform 1 0 16100 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1667941163
transform -1 0 29900 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1667941163
transform 1 0 22356 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1667941163
transform 1 0 20608 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1667941163
transform 1 0 20240 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1667941163
transform -1 0 17388 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp 1667941163
transform 1 0 15824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _232_
timestamp 1667941163
transform 1 0 16560 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _233_
timestamp 1667941163
transform -1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _234_
timestamp 1667941163
transform 1 0 28336 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1667941163
transform 1 0 15088 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1667941163
transform 1 0 20884 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 1667941163
transform -1 0 29992 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1667941163
transform -1 0 31004 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1667941163
transform -1 0 28704 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1667941163
transform -1 0 29716 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1667941163
transform -1 0 31648 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1667941163
transform 1 0 19780 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1667941163
transform 1 0 18676 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1667941163
transform 1 0 17480 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1667941163
transform -1 0 20332 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1667941163
transform -1 0 31188 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1667941163
transform -1 0 25484 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1667941163
transform -1 0 26680 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1667941163
transform -1 0 29256 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1667941163
transform -1 0 28612 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1667941163
transform -1 0 26220 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1667941163
transform 1 0 22264 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1667941163
transform -1 0 26036 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1667941163
transform -1 0 25484 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1667941163
transform -1 0 24840 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1667941163
transform 1 0 21252 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1667941163
transform -1 0 22356 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1667941163
transform -1 0 24104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1667941163
transform 1 0 20424 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1667941163
transform -1 0 20332 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1667941163
transform 1 0 17480 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1667941163
transform 1 0 30360 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1667941163
transform -1 0 26680 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1667941163
transform -1 0 27324 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1667941163
transform -1 0 28704 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1667941163
transform -1 0 25024 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1667941163
transform 1 0 17112 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1667941163
transform 1 0 22172 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1667941163
transform 1 0 22080 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1667941163
transform -1 0 31832 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1667941163
transform 1 0 27140 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1667941163
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1667941163
transform 1 0 14260 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1667941163
transform -1 0 31924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1667941163
transform -1 0 26956 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1667941163
transform 1 0 19412 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1667941163
transform 1 0 16100 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _278_
timestamp 1667941163
transform -1 0 31832 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1667941163
transform 1 0 18676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1667941163
transform -1 0 30636 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _281_
timestamp 1667941163
transform -1 0 29716 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1667941163
transform -1 0 18584 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1667941163
transform 1 0 19688 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp 1667941163
transform -1 0 29072 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1667941163
transform 1 0 14904 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1667941163
transform -1 0 16100 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _287_
timestamp 1667941163
transform 1 0 13524 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _288_
timestamp 1667941163
transform -1 0 19688 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _289_
timestamp 1667941163
transform -1 0 30084 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _290_
timestamp 1667941163
transform -1 0 16744 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _291_
timestamp 1667941163
transform 1 0 13524 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1667941163
transform -1 0 17756 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1667941163
transform 1 0 16100 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1667941163
transform 1 0 32200 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1667941163
transform -1 0 28244 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1667941163
transform 1 0 30084 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1667941163
transform 1 0 19412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1667941163
transform 1 0 31004 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1667941163
transform 1 0 23184 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 1667941163
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1667941163
transform 1 0 22172 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _303_
timestamp 1667941163
transform -1 0 18952 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1667941163
transform -1 0 27968 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1667941163
transform -1 0 14536 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _306_
timestamp 1667941163
transform -1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1667941163
transform 1 0 14260 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1667941163
transform -1 0 24104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1667941163
transform -1 0 29256 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1667941163
transform -1 0 17388 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1667941163
transform -1 0 24840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 1667941163
transform 1 0 16100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1667941163
transform -1 0 31188 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1667941163
transform -1 0 15456 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1667941163
transform 1 0 15180 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1667941163
transform 1 0 16468 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 1667941163
transform -1 0 17112 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _318_
timestamp 1667941163
transform -1 0 32568 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 1667941163
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1667941163
transform -1 0 22908 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1667941163
transform -1 0 28612 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1667941163
transform 1 0 31648 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1667941163
transform -1 0 28060 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1667941163
transform 1 0 30360 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 1667941163
transform -1 0 30544 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1667941163
transform -1 0 32568 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1667941163
transform 1 0 31372 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1667941163
transform -1 0 29992 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 1667941163
transform -1 0 29900 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 1667941163
transform -1 0 15180 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp 1667941163
transform 1 0 18676 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1667941163
transform -1 0 16008 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1667941163
transform 1 0 16836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1667941163
transform 1 0 14260 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1667941163
transform 1 0 21252 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 1667941163
transform 1 0 14996 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1667941163
transform 1 0 17020 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1667941163
transform 1 0 24564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1667941163
transform -1 0 29992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1667941163
transform -1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1667941163
transform 1 0 16836 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1667941163
transform -1 0 31280 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp 1667941163
transform -1 0 23460 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1667941163
transform -1 0 2576 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1667941163
transform 1 0 9292 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1667941163
transform -1 0 22264 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1667941163
transform 1 0 13616 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1667941163
transform -1 0 19596 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1667941163
transform 1 0 10764 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1667941163
transform -1 0 29992 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1667941163
transform 1 0 33488 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1667941163
transform -1 0 32476 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1667941163
transform 1 0 26036 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1667941163
transform -1 0 29256 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1667941163
transform -1 0 32200 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1667941163
transform -1 0 26036 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1667941163
transform -1 0 28704 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1667941163
transform -1 0 2944 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1667941163
transform 1 0 19872 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1667941163
transform 1 0 14444 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _361_
timestamp 1667941163
transform 1 0 10120 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1667941163
transform 1 0 14812 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1667941163
transform 1 0 19964 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1667941163
transform -1 0 30544 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1667941163
transform 1 0 34868 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1667941163
transform -1 0 23092 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _367_
timestamp 1667941163
transform -1 0 33488 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1667941163
transform 1 0 13524 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1667941163
transform 1 0 13340 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1667941163
transform 1 0 21988 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1667941163
transform 1 0 21252 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1667941163
transform -1 0 9384 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1667941163
transform 1 0 12420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1667941163
transform -1 0 17020 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 1667941163
transform -1 0 27600 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp 1667941163
transform -1 0 32568 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp 1667941163
transform 1 0 31556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _378_
timestamp 1667941163
transform -1 0 18584 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _379_
timestamp 1667941163
transform -1 0 19412 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _380_
timestamp 1667941163
transform -1 0 28612 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _381_
timestamp 1667941163
transform 1 0 15548 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _382_
timestamp 1667941163
transform 1 0 20792 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _383_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 24748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _384_
timestamp 1667941163
transform -1 0 20148 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _385_
timestamp 1667941163
transform -1 0 17204 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _386_
timestamp 1667941163
transform -1 0 4876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _387_
timestamp 1667941163
transform 1 0 14260 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp 1667941163
transform -1 0 31464 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _389_
timestamp 1667941163
transform 1 0 12328 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _390_
timestamp 1667941163
transform 1 0 19044 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _391_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 16376 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _392_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13984 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _393_
timestamp 1667941163
transform -1 0 35144 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _394_
timestamp 1667941163
transform -1 0 35788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _395_
timestamp 1667941163
transform -1 0 33672 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _396_
timestamp 1667941163
transform -1 0 34132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _397_
timestamp 1667941163
transform -1 0 33488 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _398_
timestamp 1667941163
transform -1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _399_
timestamp 1667941163
transform 1 0 38088 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _400_
timestamp 1667941163
transform -1 0 37904 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _401_
timestamp 1667941163
transform -1 0 37260 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _402_
timestamp 1667941163
transform -1 0 36708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _403_
timestamp 1667941163
transform 1 0 14260 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _404_
timestamp 1667941163
transform -1 0 36800 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _405_
timestamp 1667941163
transform -1 0 36156 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _406_
timestamp 1667941163
transform -1 0 35788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _407_
timestamp 1667941163
transform -1 0 34408 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _408_
timestamp 1667941163
transform -1 0 36432 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _409_
timestamp 1667941163
transform -1 0 34776 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _410_
timestamp 1667941163
transform -1 0 33580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _411_
timestamp 1667941163
transform -1 0 35144 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _412_
timestamp 1667941163
transform -1 0 37720 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _413_
timestamp 1667941163
transform 1 0 38088 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _414_
timestamp 1667941163
transform 1 0 14260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _415_
timestamp 1667941163
transform -1 0 35788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _416_
timestamp 1667941163
transform -1 0 34224 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _417_
timestamp 1667941163
transform -1 0 33028 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _418_
timestamp 1667941163
transform -1 0 36708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _419_
timestamp 1667941163
transform -1 0 34776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _420_
timestamp 1667941163
transform -1 0 35420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _421_
timestamp 1667941163
transform -1 0 36064 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _422_
timestamp 1667941163
transform -1 0 34776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _423_
timestamp 1667941163
transform -1 0 34776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _424_
timestamp 1667941163
transform -1 0 37076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _425_
timestamp 1667941163
transform 1 0 13064 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _426_
timestamp 1667941163
transform -1 0 36432 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _427_
timestamp 1667941163
transform -1 0 36708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _428_
timestamp 1667941163
transform -1 0 37720 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _429_
timestamp 1667941163
transform -1 0 34316 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 1667941163
transform -1 0 32844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _431_
timestamp 1667941163
transform -1 0 35420 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 1667941163
transform -1 0 36432 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 1667941163
transform -1 0 36064 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _434_
timestamp 1667941163
transform -1 0 35144 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _435_
timestamp 1667941163
transform -1 0 35420 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _436_
timestamp 1667941163
transform 1 0 17388 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _437_
timestamp 1667941163
transform 1 0 15272 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _438_
timestamp 1667941163
transform 1 0 26404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _439_
timestamp 1667941163
transform 1 0 17572 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _440_
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _441_
timestamp 1667941163
transform 1 0 14904 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _442_
timestamp 1667941163
transform -1 0 13892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _443_
timestamp 1667941163
transform 1 0 14536 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _444_
timestamp 1667941163
transform 1 0 23828 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _445_
timestamp 1667941163
transform 1 0 17112 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _446_
timestamp 1667941163
transform 1 0 15824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _447_
timestamp 1667941163
transform 1 0 17572 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _448_
timestamp 1667941163
transform 1 0 14444 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _449_
timestamp 1667941163
transform 1 0 13524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _450_
timestamp 1667941163
transform 1 0 14260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _451_
timestamp 1667941163
transform 1 0 16100 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _452_
timestamp 1667941163
transform -1 0 35420 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _453_
timestamp 1667941163
transform 1 0 15180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _454_
timestamp 1667941163
transform 1 0 12880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _455_
timestamp 1667941163
transform 1 0 12972 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _456_
timestamp 1667941163
transform 1 0 13432 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _457_
timestamp 1667941163
transform 1 0 16468 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _458_
timestamp 1667941163
transform 1 0 11776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _459_
timestamp 1667941163
transform 1 0 12144 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _460_
timestamp 1667941163
transform -1 0 11868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _461_
timestamp 1667941163
transform -1 0 11960 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _462_
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _463_
timestamp 1667941163
transform 1 0 12328 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _464_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19688 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _465_
timestamp 1667941163
transform -1 0 23828 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _466_
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _467_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21988 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _468_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22080 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _469_
timestamp 1667941163
transform -1 0 29256 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _470_
timestamp 1667941163
transform 1 0 27416 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _471_
timestamp 1667941163
transform 1 0 32292 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _472_
timestamp 1667941163
transform 1 0 27508 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _473_
timestamp 1667941163
transform 1 0 29716 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _474_
timestamp 1667941163
transform 1 0 27140 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _475_
timestamp 1667941163
transform 1 0 27140 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _476_
timestamp 1667941163
transform 1 0 20608 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _477_
timestamp 1667941163
transform 1 0 19688 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _478_
timestamp 1667941163
transform -1 0 21528 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _479_
timestamp 1667941163
transform 1 0 24472 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _480_
timestamp 1667941163
transform 1 0 24564 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _481_
timestamp 1667941163
transform 1 0 21988 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _482_
timestamp 1667941163
transform -1 0 31556 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _483_
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _484_
timestamp 1667941163
transform 1 0 29716 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _485_
timestamp 1667941163
transform 1 0 25392 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _486_
timestamp 1667941163
transform 1 0 20884 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _487_
timestamp 1667941163
transform 1 0 24564 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _488_
timestamp 1667941163
transform 1 0 21988 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _489_
timestamp 1667941163
transform 1 0 19688 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _490_
timestamp 1667941163
transform 1 0 17480 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _491_
timestamp 1667941163
transform 1 0 24104 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _492_
timestamp 1667941163
transform 1 0 20516 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _493_
timestamp 1667941163
transform -1 0 29992 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _494_
timestamp 1667941163
transform -1 0 33764 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _495_
timestamp 1667941163
transform 1 0 32292 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _496_
timestamp 1667941163
transform -1 0 34132 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _497_
timestamp 1667941163
transform 1 0 25852 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _498_
timestamp 1667941163
transform 1 0 20516 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _499_
timestamp 1667941163
transform 1 0 25024 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _500_
timestamp 1667941163
transform -1 0 31556 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _501_
timestamp 1667941163
transform 1 0 31924 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _502_
timestamp 1667941163
transform 1 0 24656 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _503_
timestamp 1667941163
transform 1 0 27140 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _504_
timestamp 1667941163
transform -1 0 26588 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _505_
timestamp 1667941163
transform -1 0 30176 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _506_
timestamp 1667941163
transform -1 0 31556 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _507_
timestamp 1667941163
transform -1 0 31464 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _508_
timestamp 1667941163
transform 1 0 19688 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _509_
timestamp 1667941163
transform -1 0 21528 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _510_
timestamp 1667941163
transform -1 0 26312 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _511_
timestamp 1667941163
transform -1 0 29072 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _512_
timestamp 1667941163
transform -1 0 34132 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _513_
timestamp 1667941163
transform -1 0 28612 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _514_
timestamp 1667941163
transform 1 0 21988 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _515_
timestamp 1667941163
transform -1 0 22448 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _516_
timestamp 1667941163
transform -1 0 26312 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _517_
timestamp 1667941163
transform -1 0 30912 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _518_
timestamp 1667941163
transform 1 0 27508 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _519_
timestamp 1667941163
transform -1 0 21528 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _520_
timestamp 1667941163
transform -1 0 26404 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _521_
timestamp 1667941163
transform 1 0 21988 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _522_
timestamp 1667941163
transform -1 0 23092 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _523_
timestamp 1667941163
transform -1 0 31832 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _524_
timestamp 1667941163
transform -1 0 26404 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _525_
timestamp 1667941163
transform 1 0 24196 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _526_
timestamp 1667941163
transform -1 0 26404 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _527_
timestamp 1667941163
transform 1 0 22448 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _528_
timestamp 1667941163
transform -1 0 21528 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _529_
timestamp 1667941163
transform -1 0 29256 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _541_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9752 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _542_
timestamp 1667941163
transform 1 0 6900 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _543_
timestamp 1667941163
transform -1 0 2576 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _544_
timestamp 1667941163
transform -1 0 27416 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _545_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 16376 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _546_
timestamp 1667941163
transform 1 0 21252 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _547_
timestamp 1667941163
transform -1 0 32844 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _548_
timestamp 1667941163
transform 1 0 20884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _549_
timestamp 1667941163
transform -1 0 22448 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _550_
timestamp 1667941163
transform -1 0 6624 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _551_
timestamp 1667941163
transform -1 0 23184 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _552_
timestamp 1667941163
transform -1 0 27416 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _553_
timestamp 1667941163
transform 1 0 1748 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _554_
timestamp 1667941163
transform 1 0 34132 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _555_
timestamp 1667941163
transform 1 0 25484 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _556_
timestamp 1667941163
transform -1 0 28060 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _557_
timestamp 1667941163
transform 1 0 25116 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _558_
timestamp 1667941163
transform -1 0 27416 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _559_
timestamp 1667941163
transform -1 0 27324 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _560_
timestamp 1667941163
transform 1 0 7176 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _561_
timestamp 1667941163
transform 1 0 31556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _562_
timestamp 1667941163
transform -1 0 17480 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _563_
timestamp 1667941163
transform 1 0 10488 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _564_
timestamp 1667941163
transform -1 0 30452 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _565_
timestamp 1667941163
transform 1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _566_
timestamp 1667941163
transform 1 0 9108 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _567_
timestamp 1667941163
transform 1 0 5704 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _568_
timestamp 1667941163
transform 1 0 6532 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _569_
timestamp 1667941163
transform -1 0 38088 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _570_
timestamp 1667941163
transform -1 0 36708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _571_
timestamp 1667941163
transform 1 0 5060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _572_
timestamp 1667941163
transform -1 0 23276 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _573_
timestamp 1667941163
transform -1 0 37076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _574_
timestamp 1667941163
transform -1 0 26404 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _575_
timestamp 1667941163
transform 1 0 16836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _576_
timestamp 1667941163
transform -1 0 29624 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _577_
timestamp 1667941163
transform -1 0 37628 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _578_
timestamp 1667941163
transform -1 0 26680 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  _579_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 17664 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _580_
timestamp 1667941163
transform 1 0 15548 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _581_
timestamp 1667941163
transform -1 0 26588 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _582_
timestamp 1667941163
transform -1 0 25116 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _583__91 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17572 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _583_
timestamp 1667941163
transform 1 0 17388 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _584_
timestamp 1667941163
transform 1 0 16836 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _585_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19228 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _586_
timestamp 1667941163
transform 1 0 19872 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _587_
timestamp 1667941163
transform -1 0 20240 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _588_
timestamp 1667941163
transform 1 0 18308 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _589_
timestamp 1667941163
transform -1 0 22816 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _590_
timestamp 1667941163
transform 1 0 18952 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _591_
timestamp 1667941163
transform 1 0 29716 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _592__92
timestamp 1667941163
transform 1 0 30728 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _592_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 28612 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _593_
timestamp 1667941163
transform -1 0 27876 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _594_
timestamp 1667941163
transform 1 0 27600 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _595_
timestamp 1667941163
transform -1 0 24840 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _596_
timestamp 1667941163
transform 1 0 20700 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _597_
timestamp 1667941163
transform 1 0 28520 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _598_
timestamp 1667941163
transform 1 0 25668 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _599_
timestamp 1667941163
transform 1 0 28244 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _600_
timestamp 1667941163
transform 1 0 26312 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _601_
timestamp 1667941163
transform -1 0 30360 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _602_
timestamp 1667941163
transform 1 0 24564 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _603_
timestamp 1667941163
transform -1 0 16192 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _604_
timestamp 1667941163
transform -1 0 15180 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _605_
timestamp 1667941163
transform -1 0 27968 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _606__93
timestamp 1667941163
transform -1 0 17756 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _606_
timestamp 1667941163
transform 1 0 20700 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _607_
timestamp 1667941163
transform -1 0 17204 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _608_
timestamp 1667941163
transform -1 0 17940 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _609_
timestamp 1667941163
transform -1 0 25300 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _610_
timestamp 1667941163
transform -1 0 24104 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _611_
timestamp 1667941163
transform -1 0 15456 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _612_
timestamp 1667941163
transform -1 0 23644 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _613_
timestamp 1667941163
transform 1 0 15548 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _614_
timestamp 1667941163
transform 1 0 15548 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _615_
timestamp 1667941163
transform 1 0 28060 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _616_
timestamp 1667941163
transform 1 0 26312 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _617_
timestamp 1667941163
transform 1 0 23644 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _618__94
timestamp 1667941163
transform 1 0 26036 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _618_
timestamp 1667941163
transform -1 0 25668 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _619_
timestamp 1667941163
transform 1 0 14904 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _620_
timestamp 1667941163
transform -1 0 26220 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _621_
timestamp 1667941163
transform 1 0 20700 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _622_
timestamp 1667941163
transform 1 0 23552 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _623_
timestamp 1667941163
transform 1 0 26496 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _624_
timestamp 1667941163
transform 1 0 23184 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _625_
timestamp 1667941163
transform -1 0 16376 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _626_
timestamp 1667941163
transform 1 0 25116 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _627_
timestamp 1667941163
transform -1 0 16100 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _628_
timestamp 1667941163
transform -1 0 14904 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _629_
timestamp 1667941163
transform -1 0 27876 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _630_
timestamp 1667941163
transform -1 0 18952 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _630__95
timestamp 1667941163
transform -1 0 18676 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _631_
timestamp 1667941163
transform 1 0 16836 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _632_
timestamp 1667941163
transform 1 0 19412 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _633_
timestamp 1667941163
transform 1 0 16284 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _634_
timestamp 1667941163
transform -1 0 23920 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _635_
timestamp 1667941163
transform -1 0 18032 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _636_
timestamp 1667941163
transform 1 0 14076 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _637_
timestamp 1667941163
transform 1 0 15548 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _638_
timestamp 1667941163
transform -1 0 22264 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _639_
timestamp 1667941163
transform 1 0 31004 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _640_
timestamp 1667941163
transform 1 0 27324 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _641_
timestamp 1667941163
transform 1 0 17020 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _642__96
timestamp 1667941163
transform -1 0 20332 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _642_
timestamp 1667941163
transform 1 0 20700 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _643_
timestamp 1667941163
transform -1 0 25392 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _644_
timestamp 1667941163
transform -1 0 29256 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _645_
timestamp 1667941163
transform 1 0 17112 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _646_
timestamp 1667941163
transform -1 0 18860 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _647_
timestamp 1667941163
transform 1 0 27416 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _648_
timestamp 1667941163
transform 1 0 24840 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _649_
timestamp 1667941163
transform 1 0 19504 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _650_
timestamp 1667941163
transform 1 0 27140 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _651_
timestamp 1667941163
transform -1 0 23460 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _652_
timestamp 1667941163
transform -1 0 26956 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _653_
timestamp 1667941163
transform -1 0 28060 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _654__97
timestamp 1667941163
transform 1 0 27140 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _654_
timestamp 1667941163
transform -1 0 26680 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _655_
timestamp 1667941163
transform -1 0 23552 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _656_
timestamp 1667941163
transform -1 0 23828 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _657_
timestamp 1667941163
transform 1 0 18124 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _658_
timestamp 1667941163
transform 1 0 18124 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _659_
timestamp 1667941163
transform 1 0 21068 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _660_
timestamp 1667941163
transform -1 0 26496 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _661_
timestamp 1667941163
transform 1 0 21988 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _662_
timestamp 1667941163
transform 1 0 20700 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _663_
timestamp 1667941163
transform -1 0 24288 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _664_
timestamp 1667941163
transform -1 0 25576 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _665_
timestamp 1667941163
transform -1 0 24104 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _666_
timestamp 1667941163
transform -1 0 23828 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _666__98
timestamp 1667941163
transform 1 0 23736 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _667_
timestamp 1667941163
transform 1 0 21988 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _668_
timestamp 1667941163
transform 1 0 21436 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _669_
timestamp 1667941163
transform -1 0 25944 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _670_
timestamp 1667941163
transform 1 0 23368 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _671_
timestamp 1667941163
transform -1 0 25116 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _672_
timestamp 1667941163
transform -1 0 24840 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _673_
timestamp 1667941163
transform -1 0 25392 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _674_
timestamp 1667941163
transform -1 0 25392 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _675_
timestamp 1667941163
transform 1 0 21988 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _676_
timestamp 1667941163
transform -1 0 25944 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _677_
timestamp 1667941163
transform -1 0 26680 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _678__99
timestamp 1667941163
transform 1 0 30084 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _678_
timestamp 1667941163
transform -1 0 26220 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _679_
timestamp 1667941163
transform 1 0 18124 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _680_
timestamp 1667941163
transform 1 0 17756 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _681_
timestamp 1667941163
transform -1 0 25392 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _682_
timestamp 1667941163
transform 1 0 21988 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _683_
timestamp 1667941163
transform -1 0 23920 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _684_
timestamp 1667941163
transform 1 0 25760 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _685_
timestamp 1667941163
transform 1 0 19412 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _686_
timestamp 1667941163
transform 1 0 18400 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _687_
timestamp 1667941163
transform -1 0 16008 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _688_
timestamp 1667941163
transform -1 0 21252 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _689_
timestamp 1667941163
transform 1 0 22448 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _690__100
timestamp 1667941163
transform 1 0 21068 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _690_
timestamp 1667941163
transform 1 0 20884 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _691_
timestamp 1667941163
transform 1 0 14904 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _692_
timestamp 1667941163
transform -1 0 20608 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _693_
timestamp 1667941163
transform 1 0 19412 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _694_
timestamp 1667941163
transform 1 0 17848 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _695_
timestamp 1667941163
transform 1 0 18124 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _696_
timestamp 1667941163
transform 1 0 22540 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _697_
timestamp 1667941163
transform 1 0 18032 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _698_
timestamp 1667941163
transform -1 0 23644 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _699_
timestamp 1667941163
transform -1 0 17664 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _700__101
timestamp 1667941163
transform -1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _700_
timestamp 1667941163
transform 1 0 16376 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _701_
timestamp 1667941163
transform 1 0 18032 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _702_
timestamp 1667941163
transform -1 0 19320 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _703_
timestamp 1667941163
transform -1 0 23460 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _704_
timestamp 1667941163
transform 1 0 16836 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _705_
timestamp 1667941163
transform -1 0 16376 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _706_
timestamp 1667941163
transform -1 0 25392 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _707_
timestamp 1667941163
transform -1 0 25024 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 38088 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1667941163
transform -1 0 13800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1667941163
transform -1 0 38364 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1667941163
transform -1 0 38364 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1667941163
transform -1 0 38364 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1667941163
transform -1 0 38364 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1667941163
transform -1 0 38364 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1667941163
transform 1 0 1564 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1667941163
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1667941163
transform -1 0 38364 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1667941163
transform 1 0 1564 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1667941163
transform 1 0 1564 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1667941163
transform -1 0 38364 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1667941163
transform -1 0 37812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1667941163
transform 1 0 25208 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1667941163
transform 1 0 1564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1667941163
transform -1 0 38364 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1667941163
transform 1 0 1564 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1667941163
transform 1 0 1564 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1667941163
transform -1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1667941163
transform 1 0 35788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input23 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 38364 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1667941163
transform -1 0 38364 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1667941163
transform 1 0 27140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1667941163
transform 1 0 37444 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1667941163
transform 1 0 1564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1667941163
transform -1 0 38364 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 1667941163
transform 1 0 1564 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1667941163
transform -1 0 29256 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1667941163
transform -1 0 38364 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1667941163
transform 1 0 11684 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1667941163
transform 1 0 6532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1667941163
transform -1 0 19780 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1667941163
transform -1 0 2484 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1667941163
transform 1 0 23000 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1667941163
transform -1 0 13800 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1667941163
transform -1 0 23644 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1667941163
transform 1 0 9752 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1667941163
transform -1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1667941163
transform 1 0 37444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1667941163
transform -1 0 1932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1667941163
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1667941163
transform -1 0 15272 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1667941163
transform -1 0 17204 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1667941163
transform -1 0 18492 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1667941163
transform -1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1667941163
transform 1 0 35512 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1667941163
transform -1 0 2668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1667941163
transform -1 0 30728 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1667941163
transform -1 0 1932 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1667941163
transform 1 0 28428 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1667941163
transform -1 0 35236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1667941163
transform -1 0 20424 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1667941163
transform 1 0 37996 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1667941163
transform -1 0 24104 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1667941163
transform -1 0 1932 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1667941163
transform 1 0 36616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1667941163
transform 1 0 37996 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1667941163
transform -1 0 2668 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1667941163
transform -1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1667941163
transform -1 0 1932 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1667941163
transform -1 0 1932 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1667941163
transform 1 0 37996 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1667941163
transform -1 0 8188 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1667941163
transform -1 0 3496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1667941163
transform 1 0 33580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1667941163
transform -1 0 1932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1667941163
transform -1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1667941163
transform -1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1667941163
transform 1 0 30360 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1667941163
transform -1 0 16376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1667941163
transform 1 0 36616 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1667941163
transform -1 0 4968 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1667941163
transform 1 0 37996 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1667941163
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1667941163
transform -1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1667941163
transform -1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1667941163
transform 1 0 37996 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform -1 0 18952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform -1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 2668 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform -1 0 1932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform -1 0 1932 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform 1 0 37996 0 -1 19584
box -38 -48 406 592
<< labels >>
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
port 0 nsew signal tristate
flabel metal2 s 37370 39200 37426 39800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
port 1 nsew signal tristate
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
port 2 nsew signal tristate
flabel metal2 s 35438 200 35494 800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
port 3 nsew signal tristate
flabel metal2 s 14830 39200 14886 39800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_
port 4 nsew signal tristate
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_
port 5 nsew signal tristate
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_
port 6 nsew signal tristate
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_
port 7 nsew signal tristate
flabel metal3 s 39200 8168 39800 8288 0 FreeSans 480 0 0 0 ccff_head
port 8 nsew signal input
flabel metal2 s 35438 39200 35494 39800 0 FreeSans 224 90 0 0 ccff_tail
port 9 nsew signal tristate
flabel metal2 s 21914 39200 21970 39800 0 FreeSans 224 90 0 0 chanx_left_in[0]
port 10 nsew signal input
flabel metal2 s 13542 200 13598 800 0 FreeSans 224 90 0 0 chanx_left_in[10]
port 11 nsew signal input
flabel metal3 s 39200 11568 39800 11688 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 12 nsew signal input
flabel metal3 s 39200 17008 39800 17128 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 13 nsew signal input
flabel metal3 s 39200 35368 39800 35488 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 14 nsew signal input
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 15 nsew signal input
flabel metal3 s 39200 4768 39800 4888 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 16 nsew signal input
flabel metal3 s 200 28568 800 28688 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 17 nsew signal input
flabel metal2 s 8390 200 8446 800 0 FreeSans 224 90 0 0 chanx_left_in[17]
port 18 nsew signal input
flabel metal3 s 39200 26528 39800 26648 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 19 nsew signal input
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 20 nsew signal input
flabel metal3 s 200 14288 800 14408 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 21 nsew signal input
flabel metal3 s 39200 27888 39800 28008 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 22 nsew signal input
flabel metal2 s 37370 200 37426 800 0 FreeSans 224 90 0 0 chanx_left_in[4]
port 23 nsew signal input
flabel metal2 s 25134 39200 25190 39800 0 FreeSans 224 90 0 0 chanx_left_in[5]
port 24 nsew signal input
flabel metal2 s 1306 39200 1362 39800 0 FreeSans 224 90 0 0 chanx_left_in[6]
port 25 nsew signal input
flabel metal3 s 39200 29928 39800 30048 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 26 nsew signal input
flabel metal3 s 200 19728 800 19848 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 27 nsew signal input
flabel metal3 s 200 23128 800 23248 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 28 nsew signal input
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 29 nsew signal tristate
flabel metal2 s 30286 200 30342 800 0 FreeSans 224 90 0 0 chanx_left_out[10]
port 30 nsew signal tristate
flabel metal3 s 200 34008 800 34128 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 31 nsew signal tristate
flabel metal2 s 27066 39200 27122 39800 0 FreeSans 224 90 0 0 chanx_left_out[12]
port 32 nsew signal tristate
flabel metal2 s 28354 39200 28410 39800 0 FreeSans 224 90 0 0 chanx_left_out[13]
port 33 nsew signal tristate
flabel metal2 s 34150 200 34206 800 0 FreeSans 224 90 0 0 chanx_left_out[14]
port 34 nsew signal tristate
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chanx_left_out[15]
port 35 nsew signal tristate
flabel metal3 s 39200 33328 39800 33448 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 36 nsew signal tristate
flabel metal2 s 23846 200 23902 800 0 FreeSans 224 90 0 0 chanx_left_out[17]
port 37 nsew signal tristate
flabel metal3 s 200 21088 800 21208 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 38 nsew signal tristate
flabel metal3 s 39200 688 39800 808 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 39 nsew signal tristate
flabel metal3 s 39200 15648 39800 15768 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 40 nsew signal tristate
flabel metal3 s 200 39448 800 39568 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 41 nsew signal tristate
flabel metal3 s 200 10208 800 10328 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 42 nsew signal tristate
flabel metal3 s 200 31968 800 32088 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 43 nsew signal tristate
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 44 nsew signal tristate
flabel metal3 s 39200 37408 39800 37528 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 45 nsew signal tristate
flabel metal2 s 7746 39200 7802 39800 0 FreeSans 224 90 0 0 chanx_left_out[8]
port 46 nsew signal tristate
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chanx_left_out[9]
port 47 nsew signal tristate
flabel metal2 s 9678 200 9734 800 0 FreeSans 224 90 0 0 chanx_right_in[0]
port 48 nsew signal input
flabel metal2 s 32218 200 32274 800 0 FreeSans 224 90 0 0 chanx_right_in[10]
port 49 nsew signal input
flabel metal3 s 39200 13608 39800 13728 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 50 nsew signal input
flabel metal3 s 39200 6128 39800 6248 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 51 nsew signal input
flabel metal2 s 25134 200 25190 800 0 FreeSans 224 90 0 0 chanx_right_in[13]
port 52 nsew signal input
flabel metal3 s 200 37408 800 37528 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 53 nsew signal input
flabel metal2 s 39302 200 39358 800 0 FreeSans 224 90 0 0 chanx_right_in[15]
port 54 nsew signal input
flabel metal3 s 200 8848 800 8968 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 55 nsew signal input
flabel metal3 s 39200 10208 39800 10328 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 56 nsew signal input
flabel metal3 s 200 25168 800 25288 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 57 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 chanx_right_in[1]
port 58 nsew signal input
flabel metal3 s 39200 24488 39800 24608 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 59 nsew signal input
flabel metal2 s 11610 39200 11666 39800 0 FreeSans 224 90 0 0 chanx_right_in[3]
port 60 nsew signal input
flabel metal2 s 6458 39200 6514 39800 0 FreeSans 224 90 0 0 chanx_right_in[4]
port 61 nsew signal input
flabel metal2 s 18694 200 18750 800 0 FreeSans 224 90 0 0 chanx_right_in[5]
port 62 nsew signal input
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chanx_right_in[6]
port 63 nsew signal input
flabel metal2 s 21914 200 21970 800 0 FreeSans 224 90 0 0 chanx_right_in[7]
port 64 nsew signal input
flabel metal2 s 12898 39200 12954 39800 0 FreeSans 224 90 0 0 chanx_right_in[8]
port 65 nsew signal input
flabel metal2 s 23202 39200 23258 39800 0 FreeSans 224 90 0 0 chanx_right_in[9]
port 66 nsew signal input
flabel metal2 s 33506 39200 33562 39800 0 FreeSans 224 90 0 0 chanx_right_out[0]
port 67 nsew signal tristate
flabel metal3 s 200 26528 800 26648 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 68 nsew signal tristate
flabel metal2 s 4526 200 4582 800 0 FreeSans 224 90 0 0 chanx_right_out[11]
port 69 nsew signal tristate
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 chanx_right_out[12]
port 70 nsew signal tristate
flabel metal2 s 38658 39200 38714 39800 0 FreeSans 224 90 0 0 chanx_right_out[13]
port 71 nsew signal tristate
flabel metal2 s 30286 39200 30342 39800 0 FreeSans 224 90 0 0 chanx_right_out[14]
port 72 nsew signal tristate
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 chanx_right_out[15]
port 73 nsew signal tristate
flabel metal3 s 39200 38768 39800 38888 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 74 nsew signal tristate
flabel metal3 s 39200 2728 39800 2848 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 75 nsew signal tristate
flabel metal2 s 4526 39200 4582 39800 0 FreeSans 224 90 0 0 chanx_right_out[18]
port 76 nsew signal tristate
flabel metal3 s 39200 21088 39800 21208 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 77 nsew signal tristate
flabel metal2 s 6458 200 6514 800 0 FreeSans 224 90 0 0 chanx_right_out[2]
port 78 nsew signal tristate
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 chanx_right_out[3]
port 79 nsew signal tristate
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 80 nsew signal tristate
flabel metal3 s 39200 22448 39800 22568 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 81 nsew signal tristate
flabel metal2 s 19982 200 20038 800 0 FreeSans 224 90 0 0 chanx_right_out[6]
port 82 nsew signal tristate
flabel metal3 s 200 4768 800 4888 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 83 nsew signal tristate
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 chanx_right_out[8]
port 84 nsew signal tristate
flabel metal2 s 2594 39200 2650 39800 0 FreeSans 224 90 0 0 chanx_right_out[9]
port 85 nsew signal tristate
flabel metal2 s 9678 39200 9734 39800 0 FreeSans 224 90 0 0 pReset
port 86 nsew signal input
flabel metal2 s 27066 200 27122 800 0 FreeSans 224 90 0 0 prog_clk
port 87 nsew signal input
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_
port 88 nsew signal tristate
flabel metal3 s 200 36048 800 36168 0 FreeSans 480 0 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_
port 89 nsew signal tristate
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_
port 90 nsew signal tristate
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 91 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 91 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 92 nsew ground bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal2 21114 3723 21114 3723 0 _000_
rlabel metal1 35512 4454 35512 4454 0 _001_
rlabel metal1 32637 5610 32637 5610 0 _002_
rlabel metal1 32867 6358 32867 6358 0 _003_
rlabel metal1 24702 8568 24702 8568 0 _004_
rlabel metal1 34868 7446 34868 7446 0 _005_
rlabel metal1 37030 4488 37030 4488 0 _006_
rlabel metal1 37536 5542 37536 5542 0 _007_
rlabel metal1 34868 5746 34868 5746 0 _008_
rlabel metal1 31142 6807 31142 6807 0 _009_
rlabel metal1 28566 7337 28566 7337 0 _010_
rlabel metal1 35834 6358 35834 6358 0 _011_
rlabel metal2 21666 3230 21666 3230 0 _012_
rlabel metal2 34270 4930 34270 4930 0 _013_
rlabel via2 20654 2363 20654 2363 0 _014_
rlabel via2 34638 6443 34638 6443 0 _015_
rlabel metal1 33258 6766 33258 6766 0 _016_
rlabel metal2 35006 3213 35006 3213 0 _017_
rlabel metal1 33258 4726 33258 4726 0 _018_
rlabel metal1 31287 2346 31287 2346 0 _019_
rlabel metal2 32522 5032 32522 5032 0 _020_
rlabel metal2 34086 8432 34086 8432 0 _021_
rlabel metal2 31510 5967 31510 5967 0 _022_
rlabel metal2 34546 3723 34546 3723 0 _023_
rlabel metal1 34592 2822 34592 2822 0 _024_
rlabel metal1 21535 4182 21535 4182 0 _025_
rlabel metal1 17940 2618 17940 2618 0 _026_
rlabel metal1 28842 5032 28842 5032 0 _027_
rlabel metal2 34178 3621 34178 3621 0 _028_
rlabel metal1 33626 4488 33626 4488 0 _029_
rlabel metal1 33173 3434 33173 3434 0 _030_
rlabel metal2 36570 4624 36570 4624 0 _031_
rlabel metal2 33350 2553 33350 2553 0 _032_
rlabel metal1 27278 8983 27278 8983 0 _033_
rlabel via2 21942 10013 21942 10013 0 _034_
rlabel metal1 33626 2856 33626 2856 0 _035_
rlabel metal1 32062 3400 32062 3400 0 _036_
rlabel metal1 33403 4590 33403 4590 0 _037_
rlabel metal1 31418 5848 31418 5848 0 _038_
rlabel metal1 35052 6426 35052 6426 0 _039_
rlabel metal1 15870 4046 15870 4046 0 _040_
rlabel metal2 26542 4692 26542 4692 0 _041_
rlabel metal2 17710 4913 17710 4913 0 _042_
rlabel metal1 18768 3366 18768 3366 0 _043_
rlabel metal2 15042 5491 15042 5491 0 _044_
rlabel metal1 14812 5270 14812 5270 0 _045_
rlabel metal2 14674 4930 14674 4930 0 _046_
rlabel metal1 24334 4726 24334 4726 0 _047_
rlabel via2 17250 4539 17250 4539 0 _048_
rlabel metal2 15962 4352 15962 4352 0 _049_
rlabel metal1 14720 5882 14720 5882 0 _050_
rlabel metal1 13754 4794 13754 4794 0 _051_
rlabel metal2 14398 5185 14398 5185 0 _052_
rlabel metal1 16238 4148 16238 4148 0 _053_
rlabel metal1 35006 3910 35006 3910 0 _054_
rlabel metal1 15962 3162 15962 3162 0 _055_
rlabel metal1 16192 4726 16192 4726 0 _056_
rlabel metal1 19366 7412 19366 7412 0 _057_
rlabel metal1 13570 3944 13570 3944 0 _058_
rlabel metal1 17434 4454 17434 4454 0 _059_
rlabel metal2 11914 2346 11914 2346 0 _060_
rlabel metal2 12282 3927 12282 3927 0 _061_
rlabel metal2 22862 4658 22862 4658 0 _062_
rlabel metal1 20838 5304 20838 5304 0 _063_
rlabel metal2 20102 7140 20102 7140 0 _064_
rlabel via2 12466 5083 12466 5083 0 _065_
rlabel metal1 14168 2414 14168 2414 0 _066_
rlabel metal2 14214 3298 14214 3298 0 _067_
rlabel metal2 21574 3196 21574 3196 0 _068_
rlabel metal2 14582 2176 14582 2176 0 _069_
rlabel metal1 13524 3094 13524 3094 0 _070_
rlabel metal1 19734 3434 19734 3434 0 _071_
rlabel metal1 35420 4114 35420 4114 0 _072_
rlabel metal2 17434 16184 17434 16184 0 _073_
rlabel metal2 15778 14586 15778 14586 0 _074_
rlabel metal1 27830 11220 27830 11220 0 _075_
rlabel metal1 24794 10234 24794 10234 0 _076_
rlabel metal1 17388 17850 17388 17850 0 _077_
rlabel metal1 16100 16150 16100 16150 0 _078_
rlabel metal1 19320 15062 19320 15062 0 _079_
rlabel metal2 20102 11135 20102 11135 0 _080_
rlabel metal2 20010 17306 20010 17306 0 _081_
rlabel metal1 17756 9078 17756 9078 0 _082_
rlabel metal1 21988 18326 21988 18326 0 _083_
rlabel metal1 16882 12682 16882 12682 0 _084_
rlabel metal2 30314 13090 30314 13090 0 _085_
rlabel metal2 29394 15198 29394 15198 0 _086_
rlabel metal2 27646 14042 27646 14042 0 _087_
rlabel metal2 31786 12920 31786 12920 0 _088_
rlabel metal1 24610 15096 24610 15096 0 _089_
rlabel metal1 20930 12920 20930 12920 0 _090_
rlabel metal2 28750 15470 28750 15470 0 _091_
rlabel metal1 25990 13838 25990 13838 0 _092_
rlabel metal1 28474 14008 28474 14008 0 _093_
rlabel metal1 27232 15538 27232 15538 0 _094_
rlabel metal1 30130 14892 30130 14892 0 _095_
rlabel metal1 24840 16490 24840 16490 0 _096_
rlabel metal1 15640 4794 15640 4794 0 _097_
rlabel metal1 16376 6426 16376 6426 0 _098_
rlabel metal1 28359 11798 28359 11798 0 _099_
rlabel metal2 20102 10574 20102 10574 0 _100_
rlabel metal2 16974 12988 16974 12988 0 _101_
rlabel metal1 17158 13294 17158 13294 0 _102_
rlabel metal1 28658 13974 28658 13974 0 _103_
rlabel metal1 23920 11322 23920 11322 0 _104_
rlabel metal2 15870 5950 15870 5950 0 _105_
rlabel metal2 24702 9520 24702 9520 0 _106_
rlabel metal1 15824 12886 15824 12886 0 _107_
rlabel metal1 15088 9622 15088 9622 0 _108_
rlabel metal1 29118 13294 29118 13294 0 _109_
rlabel via2 28934 14467 28934 14467 0 _110_
rlabel metal1 23092 15674 23092 15674 0 _111_
rlabel metal1 27094 15674 27094 15674 0 _112_
rlabel metal1 14766 10506 14766 10506 0 _113_
rlabel metal2 27830 10370 27830 10370 0 _114_
rlabel metal1 20930 14008 20930 14008 0 _115_
rlabel metal1 24564 12886 24564 12886 0 _116_
rlabel metal1 30590 13192 30590 13192 0 _117_
rlabel metal1 23368 17306 23368 17306 0 _118_
rlabel metal2 18814 10914 18814 10914 0 _119_
rlabel metal1 25392 15402 25392 15402 0 _120_
rlabel metal2 16606 7684 16606 7684 0 _121_
rlabel metal1 15870 6834 15870 6834 0 _122_
rlabel metal1 29854 10710 29854 10710 0 _123_
rlabel metal1 19504 6834 19504 6834 0 _124_
rlabel metal1 16652 8058 16652 8058 0 _125_
rlabel metal1 19642 8840 19642 8840 0 _126_
rlabel metal1 15778 12614 15778 12614 0 _127_
rlabel metal1 27646 12614 27646 12614 0 _128_
rlabel metal3 18124 9860 18124 9860 0 _129_
rlabel metal1 13984 3706 13984 3706 0 _130_
rlabel viali 15774 8874 15774 8874 0 _131_
rlabel metal1 20746 8058 20746 8058 0 _132_
rlabel metal1 31464 11866 31464 11866 0 _133_
rlabel metal2 31786 14824 31786 14824 0 _134_
rlabel metal2 16238 14552 16238 14552 0 _135_
rlabel metal2 20930 13498 20930 13498 0 _136_
rlabel metal2 25162 11203 25162 11203 0 _137_
rlabel metal2 30498 11407 30498 11407 0 _138_
rlabel metal1 17204 10710 17204 10710 0 _139_
rlabel metal1 18676 15130 18676 15130 0 _140_
rlabel metal2 31694 14552 31694 14552 0 _141_
rlabel metal1 25070 17544 25070 17544 0 _142_
rlabel metal1 19090 8058 19090 8058 0 _143_
rlabel metal2 27370 16558 27370 16558 0 _144_
rlabel metal1 24058 12954 24058 12954 0 _145_
rlabel via2 28934 14603 28934 14603 0 _146_
rlabel metal1 28198 16626 28198 16626 0 _147_
rlabel metal1 26588 18258 26588 18258 0 _148_
rlabel metal1 22770 14586 22770 14586 0 _149_
rlabel metal2 23598 14620 23598 14620 0 _150_
rlabel metal1 17986 13974 17986 13974 0 _151_
rlabel metal1 19274 16150 19274 16150 0 _152_
rlabel metal1 21252 12138 21252 12138 0 _153_
rlabel metal2 26266 18258 26266 18258 0 _154_
rlabel metal1 18676 12614 18676 12614 0 _155_
rlabel metal2 20930 17816 20930 17816 0 _156_
rlabel metal1 24380 19686 24380 19686 0 _157_
rlabel metal1 25990 19754 25990 19754 0 _158_
rlabel metal1 24104 17646 24104 17646 0 _159_
rlabel metal1 23000 19890 23000 19890 0 _160_
rlabel metal2 22218 19516 22218 19516 0 _161_
rlabel metal1 21528 18802 21528 18802 0 _162_
rlabel metal2 25714 15470 25714 15470 0 _163_
rlabel metal2 23598 16983 23598 16983 0 _164_
rlabel metal1 30820 13498 30820 13498 0 _165_
rlabel metal2 26082 20196 26082 20196 0 _166_
rlabel metal2 25162 20026 25162 20026 0 _167_
rlabel metal1 25208 18802 25208 18802 0 _168_
rlabel metal1 20930 12682 20930 12682 0 _169_
rlabel metal2 27646 13311 27646 13311 0 _170_
rlabel metal1 27462 12410 27462 12410 0 _171_
rlabel metal2 27278 13532 27278 13532 0 _172_
rlabel metal1 18354 14280 18354 14280 0 _173_
rlabel metal1 17802 12886 17802 12886 0 _174_
rlabel metal1 25806 14314 25806 14314 0 _175_
rlabel metal2 22218 16864 22218 16864 0 _176_
rlabel metal1 28336 11594 28336 11594 0 _177_
rlabel metal1 26220 11050 26220 11050 0 _178_
rlabel metal2 18814 15878 18814 15878 0 _179_
rlabel metal1 18630 11832 18630 11832 0 _180_
rlabel metal1 16882 6698 16882 6698 0 _181_
rlabel metal1 29440 11526 29440 11526 0 _182_
rlabel metal1 21528 16150 21528 16150 0 _183_
rlabel metal2 21114 14824 21114 14824 0 _184_
rlabel metal2 14674 10472 14674 10472 0 _185_
rlabel metal1 17802 10166 17802 10166 0 _186_
rlabel metal1 19642 13192 19642 13192 0 _187_
rlabel metal2 18078 13770 18078 13770 0 _188_
rlabel metal1 18262 8058 18262 8058 0 _189_
rlabel metal1 22632 17850 22632 17850 0 _190_
rlabel metal1 17250 13430 17250 13430 0 _191_
rlabel metal2 20746 16014 20746 16014 0 _192_
rlabel metal1 17066 5882 17066 5882 0 _193_
rlabel metal2 16974 3298 16974 3298 0 _194_
rlabel metal1 17572 8058 17572 8058 0 _195_
rlabel metal1 16376 9350 16376 9350 0 _196_
rlabel metal1 21850 7718 21850 7718 0 _197_
rlabel metal1 16054 9146 16054 9146 0 _198_
rlabel metal1 17296 5814 17296 5814 0 _199_
rlabel metal1 25162 12104 25162 12104 0 _200_
rlabel metal1 23598 9146 23598 9146 0 _201_
rlabel metal3 1188 3468 1188 3468 0 bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 37536 37094 37536 37094 0 bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal3 1188 17748 1188 17748 0 bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal2 35466 1520 35466 1520 0 bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 14950 37094 14950 37094 0 bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_
rlabel metal1 16882 37094 16882 37094 0 bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_
rlabel metal1 18170 37094 18170 37094 0 bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_
rlabel metal2 14858 1520 14858 1520 0 bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_
rlabel metal2 38318 8347 38318 8347 0 ccff_head
rlabel metal1 35604 37094 35604 37094 0 ccff_tail
rlabel metal1 21988 37298 21988 37298 0 chanx_left_in[0]
rlabel metal1 12144 2346 12144 2346 0 chanx_left_in[10]
rlabel metal2 38226 11679 38226 11679 0 chanx_left_in[11]
rlabel via2 38318 17085 38318 17085 0 chanx_left_in[12]
rlabel metal2 38318 35343 38318 35343 0 chanx_left_in[13]
rlabel via2 38318 32011 38318 32011 0 chanx_left_in[14]
rlabel metal1 38180 5270 38180 5270 0 chanx_left_in[15]
rlabel via2 1610 28645 1610 28645 0 chanx_left_in[16]
rlabel metal1 8464 2278 8464 2278 0 chanx_left_in[17]
rlabel via2 38318 26571 38318 26571 0 chanx_left_in[18]
rlabel via2 1702 30651 1702 30651 0 chanx_left_in[1]
rlabel via2 1610 14365 1610 14365 0 chanx_left_in[2]
rlabel metal2 38226 27999 38226 27999 0 chanx_left_in[3]
rlabel metal1 37536 3026 37536 3026 0 chanx_left_in[4]
rlabel metal1 25254 37230 25254 37230 0 chanx_left_in[5]
rlabel metal1 1564 37230 1564 37230 0 chanx_left_in[6]
rlabel metal2 38226 30107 38226 30107 0 chanx_left_in[7]
rlabel via2 1702 19771 1702 19771 0 chanx_left_in[8]
rlabel via2 1610 23205 1610 23205 0 chanx_left_in[9]
rlabel metal3 1740 1428 1740 1428 0 chanx_left_out[0]
rlabel metal1 30406 2822 30406 2822 0 chanx_left_out[10]
rlabel metal3 1188 34068 1188 34068 0 chanx_left_out[11]
rlabel metal1 27232 37094 27232 37094 0 chanx_left_out[12]
rlabel metal1 28520 37094 28520 37094 0 chanx_left_out[13]
rlabel metal2 34178 1520 34178 1520 0 chanx_left_out[14]
rlabel metal1 20102 37094 20102 37094 0 chanx_left_out[15]
rlabel via2 38226 33371 38226 33371 0 chanx_left_out[16]
rlabel metal2 23874 2064 23874 2064 0 chanx_left_out[17]
rlabel metal3 1188 21148 1188 21148 0 chanx_left_out[18]
rlabel metal1 37030 2278 37030 2278 0 chanx_left_out[1]
rlabel metal2 38226 15793 38226 15793 0 chanx_left_out[2]
rlabel metal1 2668 36890 2668 36890 0 chanx_left_out[3]
rlabel metal3 1188 10268 1188 10268 0 chanx_left_out[4]
rlabel metal3 1188 32028 1188 32028 0 chanx_left_out[5]
rlabel metal3 1188 6868 1188 6868 0 chanx_left_out[6]
rlabel metal2 38226 37179 38226 37179 0 chanx_left_out[7]
rlabel metal1 7866 37094 7866 37094 0 chanx_left_out[8]
rlabel metal2 3266 1520 3266 1520 0 chanx_left_out[9]
rlabel metal1 9798 2414 9798 2414 0 chanx_right_in[0]
rlabel metal1 36064 3026 36064 3026 0 chanx_right_in[10]
rlabel metal2 38318 13787 38318 13787 0 chanx_right_in[11]
rlabel metal1 38272 6290 38272 6290 0 chanx_right_in[12]
rlabel metal2 25162 1761 25162 1761 0 chanx_right_in[13]
rlabel metal2 1702 37145 1702 37145 0 chanx_right_in[14]
rlabel metal1 37582 2482 37582 2482 0 chanx_right_in[15]
rlabel via2 1702 8891 1702 8891 0 chanx_right_in[16]
rlabel via2 38318 10251 38318 10251 0 chanx_right_in[17]
rlabel via2 1610 25245 1610 25245 0 chanx_right_in[18]
rlabel metal1 29440 3502 29440 3502 0 chanx_right_in[1]
rlabel metal2 38318 24463 38318 24463 0 chanx_right_in[2]
rlabel metal1 11684 36754 11684 36754 0 chanx_right_in[3]
rlabel metal1 6578 37230 6578 37230 0 chanx_right_in[4]
rlabel metal1 18906 3434 18906 3434 0 chanx_right_in[5]
rlabel metal1 1242 2414 1242 2414 0 chanx_right_in[6]
rlabel metal2 29026 4182 29026 4182 0 chanx_right_in[7]
rlabel metal1 13340 37298 13340 37298 0 chanx_right_in[8]
rlabel metal1 23368 37230 23368 37230 0 chanx_right_in[9]
rlabel metal1 33672 37094 33672 37094 0 chanx_right_out[0]
rlabel metal3 1188 26588 1188 26588 0 chanx_right_out[10]
rlabel metal2 4554 1520 4554 1520 0 chanx_right_out[11]
rlabel metal2 1334 1792 1334 1792 0 chanx_right_out[12]
rlabel metal1 38456 36346 38456 36346 0 chanx_right_out[13]
rlabel metal1 30452 37094 30452 37094 0 chanx_right_out[14]
rlabel metal2 16790 1520 16790 1520 0 chanx_right_out[15]
rlabel metal2 36846 38131 36846 38131 0 chanx_right_out[16]
rlabel metal2 38226 3077 38226 3077 0 chanx_right_out[17]
rlabel metal1 4692 37094 4692 37094 0 chanx_right_out[18]
rlabel metal2 38226 21233 38226 21233 0 chanx_right_out[1]
rlabel metal2 6486 1520 6486 1520 0 chanx_right_out[2]
rlabel metal2 11638 1520 11638 1520 0 chanx_right_out[3]
rlabel metal3 1188 15708 1188 15708 0 chanx_right_out[4]
rlabel via2 38226 22491 38226 22491 0 chanx_right_out[5]
rlabel metal2 20010 1656 20010 1656 0 chanx_right_out[6]
rlabel metal3 1188 4828 1188 4828 0 chanx_right_out[7]
rlabel metal1 32384 37094 32384 37094 0 chanx_right_out[8]
rlabel metal1 2852 37094 2852 37094 0 chanx_right_out[9]
rlabel metal1 21436 18258 21436 18258 0 mem_bottom_ipin_0.DFFR_0_.Q
rlabel metal2 14766 14195 14766 14195 0 mem_bottom_ipin_0.DFFR_1_.Q
rlabel metal1 17434 17646 17434 17646 0 mem_bottom_ipin_0.DFFR_2_.Q
rlabel metal1 15364 11730 15364 11730 0 mem_bottom_ipin_0.DFFR_3_.Q
rlabel metal1 21528 2618 21528 2618 0 mem_bottom_ipin_0.DFFR_4_.Q
rlabel metal2 21390 5542 21390 5542 0 mem_bottom_ipin_0.DFFR_5_.Q
rlabel metal2 31418 14943 31418 14943 0 mem_bottom_ipin_1.DFFR_0_.Q
rlabel metal2 29946 14705 29946 14705 0 mem_bottom_ipin_1.DFFR_1_.Q
rlabel metal1 30636 16082 30636 16082 0 mem_bottom_ipin_1.DFFR_2_.Q
rlabel metal1 32568 13906 32568 13906 0 mem_bottom_ipin_1.DFFR_3_.Q
rlabel metal1 33074 12818 33074 12818 0 mem_bottom_ipin_1.DFFR_4_.Q
rlabel metal1 29808 2618 29808 2618 0 mem_bottom_ipin_1.DFFR_5_.Q
rlabel metal1 27508 5746 27508 5746 0 mem_bottom_ipin_2.DFFR_0_.Q
rlabel metal1 19872 7174 19872 7174 0 mem_bottom_ipin_2.DFFR_1_.Q
rlabel metal1 15226 8942 15226 8942 0 mem_bottom_ipin_2.DFFR_2_.Q
rlabel metal2 20194 5066 20194 5066 0 mem_bottom_ipin_2.DFFR_3_.Q
rlabel metal2 19090 4811 19090 4811 0 mem_bottom_ipin_2.DFFR_4_.Q
rlabel metal2 21298 3060 21298 3060 0 mem_bottom_ipin_2.DFFR_5_.Q
rlabel metal2 13386 13124 13386 13124 0 mem_top_ipin_0.DFFR_0_.Q
rlabel metal1 17296 9486 17296 9486 0 mem_top_ipin_0.DFFR_1_.Q
rlabel metal1 21206 2312 21206 2312 0 mem_top_ipin_0.DFFR_2_.Q
rlabel metal1 19918 2618 19918 2618 0 mem_top_ipin_0.DFFR_3_.Q
rlabel metal1 15686 4624 15686 4624 0 mem_top_ipin_0.DFFR_4_.Q
rlabel metal2 22402 5389 22402 5389 0 mem_top_ipin_0.DFFR_5_.Q
rlabel metal2 21850 14761 21850 14761 0 mem_top_ipin_1.DFFR_0_.Q
rlabel metal2 20102 14756 20102 14756 0 mem_top_ipin_1.DFFR_1_.Q
rlabel metal1 29992 13906 29992 13906 0 mem_top_ipin_1.DFFR_2_.Q
rlabel metal1 32430 13226 32430 13226 0 mem_top_ipin_1.DFFR_3_.Q
rlabel metal1 31326 2618 31326 2618 0 mem_top_ipin_1.DFFR_4_.Q
rlabel metal2 29440 14076 29440 14076 0 mem_top_ipin_1.DFFR_5_.Q
rlabel metal1 11799 3434 11799 3434 0 mem_top_ipin_2.DFFR_0_.Q
rlabel metal1 18998 5134 18998 5134 0 mem_top_ipin_2.DFFR_1_.Q
rlabel metal1 19642 6800 19642 6800 0 mem_top_ipin_2.DFFR_2_.Q
rlabel metal1 19918 4046 19918 4046 0 mem_top_ipin_2.DFFR_3_.Q
rlabel metal2 20746 5338 20746 5338 0 mem_top_ipin_2.DFFR_4_.Q
rlabel metal2 21942 6273 21942 6273 0 mem_top_ipin_2.DFFR_5_.Q
rlabel metal1 21344 10098 21344 10098 0 mem_top_ipin_3.DFFR_0_.Q
rlabel metal2 13754 13702 13754 13702 0 mem_top_ipin_3.DFFR_1_.Q
rlabel metal1 16146 15878 16146 15878 0 mem_top_ipin_3.DFFR_2_.Q
rlabel metal1 32476 2550 32476 2550 0 mem_top_ipin_3.DFFR_3_.Q
rlabel metal1 33994 3910 33994 3910 0 mem_top_ipin_3.DFFR_4_.Q
rlabel metal1 31970 14382 31970 14382 0 mem_top_ipin_3.DFFR_5_.Q
rlabel metal1 17066 12818 17066 12818 0 mem_top_ipin_4.DFFR_0_.Q
rlabel metal2 17526 14246 17526 14246 0 mem_top_ipin_4.DFFR_1_.Q
rlabel metal1 17710 17578 17710 17578 0 mem_top_ipin_4.DFFR_2_.Q
rlabel metal1 26082 13498 26082 13498 0 mem_top_ipin_4.DFFR_3_.Q
rlabel metal2 32062 3655 32062 3655 0 mem_top_ipin_4.DFFR_4_.Q
rlabel metal1 30268 14382 30268 14382 0 mem_top_ipin_4.DFFR_5_.Q
rlabel metal1 25806 20434 25806 20434 0 mem_top_ipin_5.DFFR_0_.Q
rlabel metal2 29210 16252 29210 16252 0 mem_top_ipin_5.DFFR_1_.Q
rlabel metal2 22034 20604 22034 20604 0 mem_top_ipin_5.DFFR_2_.Q
rlabel metal1 31004 8534 31004 8534 0 mem_top_ipin_5.DFFR_3_.Q
rlabel metal1 28750 8432 28750 8432 0 mem_top_ipin_5.DFFR_4_.Q
rlabel metal1 29716 5814 29716 5814 0 mem_top_ipin_5.DFFR_5_.Q
rlabel metal1 17250 17034 17250 17034 0 mem_top_ipin_6.DFFR_0_.Q
rlabel via2 22034 14365 22034 14365 0 mem_top_ipin_6.DFFR_1_.Q
rlabel metal1 17526 14450 17526 14450 0 mem_top_ipin_6.DFFR_2_.Q
rlabel metal2 28290 7159 28290 7159 0 mem_top_ipin_6.DFFR_3_.Q
rlabel metal2 16330 12019 16330 12019 0 mem_top_ipin_6.DFFR_4_.Q
rlabel metal2 31878 12585 31878 12585 0 mem_top_ipin_6.DFFR_5_.Q
rlabel metal1 15824 13294 15824 13294 0 mem_top_ipin_7.DFFR_0_.Q
rlabel viali 16146 14993 16146 14993 0 mem_top_ipin_7.DFFR_1_.Q
rlabel metal1 16882 14348 16882 14348 0 mem_top_ipin_7.DFFR_2_.Q
rlabel metal1 18262 7820 18262 7820 0 mem_top_ipin_7.DFFR_3_.Q
rlabel metal2 19734 4862 19734 4862 0 mem_top_ipin_7.DFFR_4_.Q
rlabel metal1 22540 27846 22540 27846 0 mux_bottom_ipin_0.INVTX1_0_.out
rlabel metal1 14720 14314 14720 14314 0 mux_bottom_ipin_0.INVTX1_1_.out
rlabel metal1 18860 16014 18860 16014 0 mux_bottom_ipin_0.INVTX1_2_.out
rlabel metal2 18446 10404 18446 10404 0 mux_bottom_ipin_0.INVTX1_3_.out
rlabel metal1 25070 11798 25070 11798 0 mux_bottom_ipin_0.INVTX1_4_.out
rlabel metal2 27462 12002 27462 12002 0 mux_bottom_ipin_0.INVTX1_5_.out
rlabel metal1 23092 22950 23092 22950 0 mux_bottom_ipin_0.INVTX1_6_.out
rlabel metal2 16974 17680 16974 17680 0 mux_bottom_ipin_0.INVTX1_7_.out
rlabel metal1 19389 16626 19389 16626 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 20010 11016 20010 11016 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 17618 16184 17618 16184 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 2806 34578 2806 34578 0 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 24886 14926 24886 14926 0 mux_bottom_ipin_1.INVTX1_2_.out
rlabel metal1 25714 14926 25714 14926 0 mux_bottom_ipin_1.INVTX1_3_.out
rlabel metal2 25714 14212 25714 14212 0 mux_bottom_ipin_1.INVTX1_4_.out
rlabel metal1 28474 14994 28474 14994 0 mux_bottom_ipin_1.INVTX1_5_.out
rlabel metal1 29394 27302 29394 27302 0 mux_bottom_ipin_1.INVTX1_6_.out
rlabel metal2 28014 15232 28014 15232 0 mux_bottom_ipin_1.INVTX1_7_.out
rlabel metal2 24150 14178 24150 14178 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 29348 14790 29348 14790 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 27094 14042 27094 14042 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 33534 14586 33534 14586 0 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 15594 9486 15594 9486 0 mux_bottom_ipin_2.INVTX1_2_.out
rlabel metal1 25622 14450 25622 14450 0 mux_bottom_ipin_2.INVTX1_3_.out
rlabel metal1 16836 8398 16836 8398 0 mux_bottom_ipin_2.INVTX1_4_.out
rlabel metal1 19366 8874 19366 8874 0 mux_bottom_ipin_2.INVTX1_5_.out
rlabel metal2 17618 9588 17618 9588 0 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 18906 9452 18906 9452 0 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 5106 9554 5106 9554 0 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 23506 16014 23506 16014 0 mux_top_ipin_0.INVTX1_2_.out
rlabel metal1 15272 27302 15272 27302 0 mux_top_ipin_0.INVTX1_3_.out
rlabel via1 18262 14331 18262 14331 0 mux_top_ipin_0.INVTX1_4_.out
rlabel metal1 18078 12274 18078 12274 0 mux_top_ipin_0.INVTX1_5_.out
rlabel metal1 24380 10098 24380 10098 0 mux_top_ipin_0.INVTX1_6_.out
rlabel metal1 27692 11662 27692 11662 0 mux_top_ipin_0.INVTX1_7_.out
rlabel metal2 16330 9503 16330 9503 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 16192 12886 16192 12886 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 18170 9146 18170 9146 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 4899 5678 4899 5678 0 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 23598 12886 23598 12886 0 mux_top_ipin_1.INVTX1_2_.out
rlabel metal1 14858 11662 14858 11662 0 mux_top_ipin_1.INVTX1_3_.out
rlabel metal1 14352 11050 14352 11050 0 mux_top_ipin_1.INVTX1_4_.out
rlabel metal2 30130 10608 30130 10608 0 mux_top_ipin_1.INVTX1_5_.out
rlabel metal2 22678 20332 22678 20332 0 mux_top_ipin_1.INVTX1_6_.out
rlabel metal2 22586 16490 22586 16490 0 mux_top_ipin_1.INVTX1_7_.out
rlabel metal1 23690 12750 23690 12750 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 15594 11288 15594 11288 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 24058 17102 24058 17102 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 35236 36754 35236 36754 0 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 27048 16014 27048 16014 0 mux_top_ipin_2.INVTX1_2_.out
rlabel metal1 17066 7990 17066 7990 0 mux_top_ipin_2.INVTX1_3_.out
rlabel metal2 12558 3604 12558 3604 0 mux_top_ipin_2.INVTX1_6_.out
rlabel via2 29026 12291 29026 12291 0 mux_top_ipin_2.INVTX1_7_.out
rlabel metal2 21482 11356 21482 11356 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 17526 8670 17526 8670 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 18354 8874 18354 8874 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 11730 14382 11730 14382 0 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 17940 15402 17940 15402 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 20286 10540 20286 10540 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 21206 14110 21206 14110 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 31464 5202 31464 5202 0 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 19964 15946 19964 15946 0 mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 23138 15062 23138 15062 0 mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 25898 17306 25898 17306 0 mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 20102 27302 20102 27302 0 mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 22034 19244 22034 19244 0 mux_top_ipin_5.INVTX1_4_.out
rlabel metal1 16376 16762 16376 16762 0 mux_top_ipin_5.INVTX1_5_.out
rlabel metal1 26680 27914 26680 27914 0 mux_top_ipin_5.INVTX1_6_.out
rlabel metal1 24288 17714 24288 17714 0 mux_top_ipin_5.INVTX1_7_.out
rlabel metal2 24978 16082 24978 16082 0 mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 24426 19414 24426 19414 0 mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 23138 18768 23138 18768 0 mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 22080 27982 22080 27982 0 mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 23690 12274 23690 12274 0 mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 18906 13498 18906 13498 0 mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 25852 12750 25852 12750 0 mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 21896 28390 21896 28390 0 mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 18722 13226 18722 13226 0 mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 19320 12206 19320 12206 0 mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 21666 14280 21666 14280 0 mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 17802 6902 17802 6902 0 mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 35466 8602 35466 8602 0 net1
rlabel metal2 36846 7276 36846 7276 0 net10
rlabel metal2 21022 14620 21022 14620 0 net100
rlabel metal1 16238 3434 16238 3434 0 net101
rlabel metal1 23782 23290 23782 23290 0 net11
rlabel metal1 2070 30634 2070 30634 0 net12
rlabel metal2 5566 12750 5566 12750 0 net13
rlabel metal1 37996 27914 37996 27914 0 net14
rlabel metal1 37628 3094 37628 3094 0 net15
rlabel metal1 32936 21522 32936 21522 0 net16
rlabel metal2 1702 21692 1702 21692 0 net17
rlabel metal2 38134 22304 38134 22304 0 net18
rlabel metal1 27094 30702 27094 30702 0 net19
rlabel metal2 22310 36992 22310 36992 0 net2
rlabel metal2 1886 21182 1886 21182 0 net20
rlabel metal1 7682 3026 7682 3026 0 net21
rlabel metal1 33580 10642 33580 10642 0 net22
rlabel metal1 37766 14042 37766 14042 0 net23
rlabel metal2 37582 9214 37582 9214 0 net24
rlabel metal1 28290 32198 28290 32198 0 net25
rlabel metal1 2024 36618 2024 36618 0 net26
rlabel metal1 38088 2482 38088 2482 0 net27
rlabel metal2 1886 10676 1886 10676 0 net28
rlabel metal1 36248 10642 36248 10642 0 net29
rlabel metal1 13432 2550 13432 2550 0 net3
rlabel metal2 1978 20128 1978 20128 0 net30
rlabel metal2 32430 5916 32430 5916 0 net31
rlabel metal1 37950 24718 37950 24718 0 net32
rlabel metal1 6831 36754 6831 36754 0 net33
rlabel metal1 6716 37298 6716 37298 0 net34
rlabel metal1 9568 25262 9568 25262 0 net35
rlabel metal1 2346 2482 2346 2482 0 net36
rlabel metal1 30544 30226 30544 30226 0 net37
rlabel metal1 13478 37196 13478 37196 0 net38
rlabel metal1 20332 37366 20332 37366 0 net39
rlabel metal1 10258 5202 10258 5202 0 net4
rlabel metal1 10810 37298 10810 37298 0 net40
rlabel metal1 2346 3502 2346 3502 0 net41
rlabel metal2 36294 36992 36294 36992 0 net42
rlabel metal1 2990 18258 2990 18258 0 net43
rlabel metal1 35650 2380 35650 2380 0 net44
rlabel metal2 15226 32674 15226 32674 0 net45
rlabel metal1 18216 28186 18216 28186 0 net46
rlabel metal1 19228 28730 19228 28730 0 net47
rlabel metal1 15502 2448 15502 2448 0 net48
rlabel metal1 34914 37094 34914 37094 0 net49
rlabel metal1 26634 14994 26634 14994 0 net5
rlabel metal1 3864 3026 3864 3026 0 net50
rlabel metal1 31050 3026 31050 3026 0 net51
rlabel metal1 1978 34578 1978 34578 0 net52
rlabel metal1 26910 37230 26910 37230 0 net53
rlabel metal1 27922 37230 27922 37230 0 net54
rlabel metal1 35512 2482 35512 2482 0 net55
rlabel metal1 20838 37264 20838 37264 0 net56
rlabel metal1 37766 33490 37766 33490 0 net57
rlabel metal2 33810 4182 33810 4182 0 net58
rlabel metal2 1794 21318 1794 21318 0 net59
rlabel metal1 37720 35598 37720 35598 0 net6
rlabel metal2 36662 2618 36662 2618 0 net60
rlabel metal2 38042 15878 38042 15878 0 net61
rlabel metal1 4600 36754 4600 36754 0 net62
rlabel metal1 3818 10642 3818 10642 0 net63
rlabel metal1 5520 32402 5520 32402 0 net64
rlabel metal1 2116 7378 2116 7378 0 net65
rlabel metal1 37674 36754 37674 36754 0 net66
rlabel metal1 9338 36890 9338 36890 0 net67
rlabel via2 4094 2499 4094 2499 0 net68
rlabel metal1 30498 36890 30498 36890 0 net69
rlabel metal1 28980 35666 28980 35666 0 net7
rlabel metal1 4370 26962 4370 26962 0 net70
rlabel metal1 4922 2448 4922 2448 0 net71
rlabel metal1 2116 3026 2116 3026 0 net72
rlabel metal1 37812 36142 37812 36142 0 net73
rlabel metal1 29992 35802 29992 35802 0 net74
rlabel metal1 16606 2414 16606 2414 0 net75
rlabel metal1 36662 37196 36662 37196 0 net76
rlabel metal1 37536 3502 37536 3502 0 net77
rlabel metal1 5198 37230 5198 37230 0 net78
rlabel metal2 38042 20910 38042 20910 0 net79
rlabel metal1 20470 5678 20470 5678 0 net8
rlabel metal2 6578 4522 6578 4522 0 net80
rlabel metal1 10810 3706 10810 3706 0 net81
rlabel metal2 2438 15742 2438 15742 0 net82
rlabel metal2 36018 22134 36018 22134 0 net83
rlabel metal3 20171 2652 20171 2652 0 net84
rlabel metal1 2116 5202 2116 5202 0 net85
rlabel metal1 31510 37230 31510 37230 0 net86
rlabel metal1 2622 37230 2622 37230 0 net87
rlabel metal1 4416 9622 4416 9622 0 net88
rlabel metal1 2162 34714 2162 34714 0 net89
rlabel metal2 25622 28594 25622 28594 0 net9
rlabel metal1 35834 19346 35834 19346 0 net90
rlabel metal2 17526 18462 17526 18462 0 net91
rlabel metal2 28934 15079 28934 15079 0 net92
rlabel metal2 20838 10914 20838 10914 0 net93
rlabel metal1 25806 16014 25806 16014 0 net94
rlabel metal1 18722 7514 18722 7514 0 net95
rlabel metal2 20838 13668 20838 13668 0 net96
rlabel metal1 26910 18190 26910 18190 0 net97
rlabel metal2 23782 19312 23782 19312 0 net98
rlabel metal1 26081 12920 26081 12920 0 net99
rlabel metal1 9798 37230 9798 37230 0 pReset
rlabel metal1 12052 2618 12052 2618 0 prog_clk
rlabel metal3 1188 12308 1188 12308 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_
rlabel metal3 1188 36108 1188 36108 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_
rlabel via2 38226 19125 38226 19125 0 top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
