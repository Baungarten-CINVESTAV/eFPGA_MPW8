magic
tech sky130A
magscale 1 2
timestamp 1672417051
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 14 2128 39362 37664
<< metal2 >>
rect 662 39200 718 39800
rect 6458 39200 6514 39800
rect 11610 39200 11666 39800
rect 17406 39200 17462 39800
rect 23202 39200 23258 39800
rect 28354 39200 28410 39800
rect 34150 39200 34206 39800
rect 39302 39200 39358 39800
rect 18 200 74 800
rect 5170 200 5226 800
rect 10966 200 11022 800
rect 16118 200 16174 800
rect 21914 200 21970 800
rect 27710 200 27766 800
rect 32862 200 32918 800
rect 38658 200 38714 800
<< obsm2 >>
rect 20 39144 606 39250
rect 774 39144 6402 39250
rect 6570 39144 11554 39250
rect 11722 39144 17350 39250
rect 17518 39144 23146 39250
rect 23314 39144 28298 39250
rect 28466 39144 34094 39250
rect 34262 39144 39246 39250
rect 20 856 39356 39144
rect 130 734 5114 856
rect 5282 734 10910 856
rect 11078 734 16062 856
rect 16230 734 21858 856
rect 22026 734 27654 856
rect 27822 734 32806 856
rect 32974 734 38602 856
rect 38770 734 39356 856
<< metal3 >>
rect 200 34688 800 34808
rect 39200 34008 39800 34128
rect 200 29248 800 29368
rect 39200 27888 39800 28008
rect 200 23128 800 23248
rect 39200 22448 39800 22568
rect 200 17008 800 17128
rect 39200 16328 39800 16448
rect 200 11568 800 11688
rect 39200 10208 39800 10328
rect 200 5448 800 5568
rect 39200 4768 39800 4888
<< obsm3 >>
rect 800 34888 39200 37569
rect 880 34608 39200 34888
rect 800 34208 39200 34608
rect 800 33928 39120 34208
rect 800 29448 39200 33928
rect 880 29168 39200 29448
rect 800 28088 39200 29168
rect 800 27808 39120 28088
rect 800 23328 39200 27808
rect 880 23048 39200 23328
rect 800 22648 39200 23048
rect 800 22368 39120 22648
rect 800 17208 39200 22368
rect 880 16928 39200 17208
rect 800 16528 39200 16928
rect 800 16248 39120 16528
rect 800 11768 39200 16248
rect 880 11488 39200 11768
rect 800 10408 39200 11488
rect 800 10128 39120 10408
rect 800 5648 39200 10128
rect 880 5368 39200 5648
rect 800 4968 39200 5368
rect 800 4688 39120 4968
rect 800 2143 39200 4688
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< labels >>
rlabel metal3 s 200 5448 800 5568 6 ccff_head
port 1 nsew signal input
rlabel metal2 s 39302 39200 39358 39800 6 ccff_tail
port 2 nsew signal output
rlabel metal3 s 200 34688 800 34808 6 gfpga_pad_GPIO_PAD[0]
port 3 nsew signal bidirectional
rlabel metal3 s 200 11568 800 11688 6 gfpga_pad_GPIO_PAD[1]
port 4 nsew signal bidirectional
rlabel metal2 s 11610 39200 11666 39800 6 gfpga_pad_GPIO_PAD[2]
port 5 nsew signal bidirectional
rlabel metal2 s 17406 39200 17462 39800 6 gfpga_pad_GPIO_PAD[3]
port 6 nsew signal bidirectional
rlabel metal3 s 39200 10208 39800 10328 6 gfpga_pad_GPIO_PAD[4]
port 7 nsew signal bidirectional
rlabel metal2 s 34150 39200 34206 39800 6 gfpga_pad_GPIO_PAD[5]
port 8 nsew signal bidirectional
rlabel metal2 s 27710 200 27766 800 6 gfpga_pad_GPIO_PAD[6]
port 9 nsew signal bidirectional
rlabel metal3 s 39200 22448 39800 22568 6 gfpga_pad_GPIO_PAD[7]
port 10 nsew signal bidirectional
rlabel metal2 s 28354 39200 28410 39800 6 pReset
port 11 nsew signal input
rlabel metal2 s 38658 200 38714 800 6 prog_clk
port 12 nsew signal input
rlabel metal3 s 200 17008 800 17128 6 top_width_0_height_0_subtile_0__pin_inpad_0_
port 13 nsew signal output
rlabel metal2 s 6458 39200 6514 39800 6 top_width_0_height_0_subtile_0__pin_outpad_0_
port 14 nsew signal input
rlabel metal2 s 32862 200 32918 800 6 top_width_0_height_0_subtile_1__pin_inpad_0_
port 15 nsew signal output
rlabel metal2 s 18 200 74 800 6 top_width_0_height_0_subtile_1__pin_outpad_0_
port 16 nsew signal input
rlabel metal2 s 5170 200 5226 800 6 top_width_0_height_0_subtile_2__pin_inpad_0_
port 17 nsew signal output
rlabel metal2 s 10966 200 11022 800 6 top_width_0_height_0_subtile_2__pin_outpad_0_
port 18 nsew signal input
rlabel metal3 s 39200 4768 39800 4888 6 top_width_0_height_0_subtile_3__pin_inpad_0_
port 19 nsew signal output
rlabel metal2 s 16118 200 16174 800 6 top_width_0_height_0_subtile_3__pin_outpad_0_
port 20 nsew signal input
rlabel metal3 s 39200 27888 39800 28008 6 top_width_0_height_0_subtile_4__pin_inpad_0_
port 21 nsew signal output
rlabel metal3 s 39200 34008 39800 34128 6 top_width_0_height_0_subtile_4__pin_outpad_0_
port 22 nsew signal input
rlabel metal3 s 200 29248 800 29368 6 top_width_0_height_0_subtile_5__pin_inpad_0_
port 23 nsew signal output
rlabel metal2 s 23202 39200 23258 39800 6 top_width_0_height_0_subtile_5__pin_outpad_0_
port 24 nsew signal input
rlabel metal2 s 21914 200 21970 800 6 top_width_0_height_0_subtile_6__pin_inpad_0_
port 25 nsew signal output
rlabel metal3 s 200 23128 800 23248 6 top_width_0_height_0_subtile_6__pin_outpad_0_
port 26 nsew signal input
rlabel metal2 s 662 39200 718 39800 6 top_width_0_height_0_subtile_7__pin_inpad_0_
port 27 nsew signal output
rlabel metal3 s 39200 16328 39800 16448 6 top_width_0_height_0_subtile_7__pin_outpad_0_
port 28 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 29 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 29 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 30 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 600054
string GDS_FILE /home/baungarten/Proyectos_caravel/FPGA_3/openlane/grid_io_bottom/runs/22_12_30_10_17/results/signoff/grid_io_bottom.magic.gds
string GDS_START 94596
<< end >>

