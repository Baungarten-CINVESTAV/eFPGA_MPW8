magic
tech sky130A
magscale 1 2
timestamp 1672461796
<< obsli1 >>
rect 1090 1959 560818 587337
<< obsm1 >>
rect 0 1576 560878 587368
<< metal2 >>
rect 5156 589000 5212 589600
rect 21900 589000 21956 589600
rect 38644 589000 38700 589600
rect 55388 589000 55444 589600
rect 72132 589000 72188 589600
rect 88232 589000 88288 589600
rect 104976 589000 105032 589600
rect 121720 589000 121776 589600
rect 138464 589000 138520 589600
rect 155208 589000 155264 589600
rect 171308 589000 171364 589600
rect 188052 589000 188108 589600
rect 204796 589000 204852 589600
rect 221540 589000 221596 589600
rect 238284 589000 238340 589600
rect 254384 589000 254440 589600
rect 271128 589000 271184 589600
rect 287872 589000 287928 589600
rect 304616 589000 304672 589600
rect 321360 589000 321416 589600
rect 337460 589000 337516 589600
rect 354204 589000 354260 589600
rect 370948 589000 371004 589600
rect 387692 589000 387748 589600
rect 403792 589000 403848 589600
rect 420536 589000 420592 589600
rect 437280 589000 437336 589600
rect 454024 589000 454080 589600
rect 470768 589000 470824 589600
rect 486868 589000 486924 589600
rect 503612 589000 503668 589600
rect 520356 589000 520412 589600
rect 537100 589000 537156 589600
rect 553844 589000 553900 589600
rect 4 0 60 600
rect 16104 0 16160 600
rect 32848 0 32904 600
rect 49592 0 49648 600
rect 66336 0 66392 600
rect 82436 0 82492 600
rect 99180 0 99236 600
rect 115924 0 115980 600
rect 132668 0 132724 600
rect 149412 0 149468 600
rect 165512 0 165568 600
rect 182256 0 182312 600
rect 199000 0 199056 600
rect 215744 0 215800 600
rect 232488 0 232544 600
rect 248588 0 248644 600
rect 265332 0 265388 600
rect 282076 0 282132 600
rect 298820 0 298876 600
rect 315564 0 315620 600
rect 331664 0 331720 600
rect 348408 0 348464 600
rect 365152 0 365208 600
rect 381896 0 381952 600
rect 398640 0 398696 600
rect 414740 0 414796 600
rect 431484 0 431540 600
rect 448228 0 448284 600
rect 464972 0 465028 600
rect 481072 0 481128 600
rect 497816 0 497872 600
rect 514560 0 514616 600
rect 531304 0 531360 600
rect 548048 0 548104 600
<< obsm2 >>
rect 6 588944 5100 589034
rect 5268 588944 21844 589034
rect 22012 588944 38588 589034
rect 38756 588944 55332 589034
rect 55500 588944 72076 589034
rect 72244 588944 88176 589034
rect 88344 588944 104920 589034
rect 105088 588944 121664 589034
rect 121832 588944 138408 589034
rect 138576 588944 155152 589034
rect 155320 588944 171252 589034
rect 171420 588944 187996 589034
rect 188164 588944 204740 589034
rect 204908 588944 221484 589034
rect 221652 588944 238228 589034
rect 238396 588944 254328 589034
rect 254496 588944 271072 589034
rect 271240 588944 287816 589034
rect 287984 588944 304560 589034
rect 304728 588944 321304 589034
rect 321472 588944 337404 589034
rect 337572 588944 354148 589034
rect 354316 588944 370892 589034
rect 371060 588944 387636 589034
rect 387804 588944 403736 589034
rect 403904 588944 420480 589034
rect 420648 588944 437224 589034
rect 437392 588944 453968 589034
rect 454136 588944 470712 589034
rect 470880 588944 486812 589034
rect 486980 588944 503556 589034
rect 503724 588944 520300 589034
rect 520468 588944 537044 589034
rect 537212 588944 553788 589034
rect 553956 588944 560338 589034
rect 6 656 560338 588944
rect 116 534 16048 656
rect 16216 534 32792 656
rect 32960 534 49536 656
rect 49704 534 66280 656
rect 66448 534 82380 656
rect 82548 534 99124 656
rect 99292 534 115868 656
rect 116036 534 132612 656
rect 132780 534 149356 656
rect 149524 534 165456 656
rect 165624 534 182200 656
rect 182368 534 198944 656
rect 199112 534 215688 656
rect 215856 534 232432 656
rect 232600 534 248532 656
rect 248700 534 265276 656
rect 265444 534 282020 656
rect 282188 534 298764 656
rect 298932 534 315508 656
rect 315676 534 331608 656
rect 331776 534 348352 656
rect 348520 534 365096 656
rect 365264 534 381840 656
rect 382008 534 398584 656
rect 398752 534 414684 656
rect 414852 534 431428 656
rect 431596 534 448172 656
rect 448340 534 464916 656
rect 465084 534 481016 656
rect 481184 534 497760 656
rect 497928 534 514504 656
rect 514672 534 531248 656
rect 531416 534 547992 656
rect 548160 534 560338 656
<< metal3 >>
rect 561186 581208 561786 581328
rect 186 578488 786 578608
rect 561186 563528 561786 563648
rect 186 560808 786 560928
rect 561186 545848 561786 545968
rect 186 543128 786 543248
rect 561186 528168 561786 528288
rect 186 525448 786 525568
rect 561186 510488 561786 510608
rect 186 507768 786 507888
rect 561186 493488 561786 493608
rect 186 490768 786 490888
rect 561186 475808 561786 475928
rect 186 473088 786 473208
rect 561186 458128 561786 458248
rect 186 455408 786 455528
rect 561186 440448 561786 440568
rect 186 437728 786 437848
rect 561186 422768 561786 422888
rect 186 420728 786 420848
rect 561186 405768 561786 405888
rect 186 403048 786 403168
rect 561186 388088 561786 388208
rect 186 385368 786 385488
rect 561186 370408 561786 370528
rect 186 367688 786 367808
rect 561186 352728 561786 352848
rect 186 350008 786 350128
rect 561186 335728 561786 335848
rect 186 333008 786 333128
rect 561186 318048 561786 318168
rect 186 315328 786 315448
rect 561186 300368 561786 300488
rect 186 297648 786 297768
rect 561186 282688 561786 282808
rect 186 279968 786 280088
rect 561186 265008 561786 265128
rect 186 262288 786 262408
rect 561186 248008 561786 248128
rect 186 245288 786 245408
rect 561186 230328 561786 230448
rect 186 227608 786 227728
rect 561186 212648 561786 212768
rect 186 209928 786 210048
rect 561186 194968 561786 195088
rect 186 192248 786 192368
rect 561186 177288 561786 177408
rect 186 174568 786 174688
rect 561186 160288 561786 160408
rect 186 157568 786 157688
rect 561186 142608 561786 142728
rect 186 139888 786 140008
rect 561186 124928 561786 125048
rect 186 122208 786 122328
rect 561186 107248 561786 107368
rect 186 104528 786 104648
rect 561186 89568 561786 89688
rect 186 86848 786 86968
rect 561186 72568 561786 72688
rect 186 69848 786 69968
rect 561186 54888 561786 55008
rect 186 52168 786 52288
rect 561186 37208 561786 37328
rect 186 34488 786 34608
rect 561186 19528 561786 19648
rect 186 16808 786 16928
rect 561186 1848 561786 1968
<< obsm3 >>
rect 786 581408 561186 587353
rect 786 581128 561106 581408
rect 786 578688 561186 581128
rect 866 578408 561186 578688
rect 786 563728 561186 578408
rect 786 563448 561106 563728
rect 786 561008 561186 563448
rect 866 560728 561186 561008
rect 786 546048 561186 560728
rect 786 545768 561106 546048
rect 786 543328 561186 545768
rect 866 543048 561186 543328
rect 786 528368 561186 543048
rect 786 528088 561106 528368
rect 786 525648 561186 528088
rect 866 525368 561186 525648
rect 786 510688 561186 525368
rect 786 510408 561106 510688
rect 786 507968 561186 510408
rect 866 507688 561186 507968
rect 786 493688 561186 507688
rect 786 493408 561106 493688
rect 786 490968 561186 493408
rect 866 490688 561186 490968
rect 786 476008 561186 490688
rect 786 475728 561106 476008
rect 786 473288 561186 475728
rect 866 473008 561186 473288
rect 786 458328 561186 473008
rect 786 458048 561106 458328
rect 786 455608 561186 458048
rect 866 455328 561186 455608
rect 786 440648 561186 455328
rect 786 440368 561106 440648
rect 786 437928 561186 440368
rect 866 437648 561186 437928
rect 786 422968 561186 437648
rect 786 422688 561106 422968
rect 786 420928 561186 422688
rect 866 420648 561186 420928
rect 786 405968 561186 420648
rect 786 405688 561106 405968
rect 786 403248 561186 405688
rect 866 402968 561186 403248
rect 786 388288 561186 402968
rect 786 388008 561106 388288
rect 786 385568 561186 388008
rect 866 385288 561186 385568
rect 786 370608 561186 385288
rect 786 370328 561106 370608
rect 786 367888 561186 370328
rect 866 367608 561186 367888
rect 786 352928 561186 367608
rect 786 352648 561106 352928
rect 786 350208 561186 352648
rect 866 349928 561186 350208
rect 786 335928 561186 349928
rect 786 335648 561106 335928
rect 786 333208 561186 335648
rect 866 332928 561186 333208
rect 786 318248 561186 332928
rect 786 317968 561106 318248
rect 786 315528 561186 317968
rect 866 315248 561186 315528
rect 786 300568 561186 315248
rect 786 300288 561106 300568
rect 786 297848 561186 300288
rect 866 297568 561186 297848
rect 786 282888 561186 297568
rect 786 282608 561106 282888
rect 786 280168 561186 282608
rect 866 279888 561186 280168
rect 786 265208 561186 279888
rect 786 264928 561106 265208
rect 786 262488 561186 264928
rect 866 262208 561186 262488
rect 786 248208 561186 262208
rect 786 247928 561106 248208
rect 786 245488 561186 247928
rect 866 245208 561186 245488
rect 786 230528 561186 245208
rect 786 230248 561106 230528
rect 786 227808 561186 230248
rect 866 227528 561186 227808
rect 786 212848 561186 227528
rect 786 212568 561106 212848
rect 786 210128 561186 212568
rect 866 209848 561186 210128
rect 786 195168 561186 209848
rect 786 194888 561106 195168
rect 786 192448 561186 194888
rect 866 192168 561186 192448
rect 786 177488 561186 192168
rect 786 177208 561106 177488
rect 786 174768 561186 177208
rect 866 174488 561186 174768
rect 786 160488 561186 174488
rect 786 160208 561106 160488
rect 786 157768 561186 160208
rect 866 157488 561186 157768
rect 786 142808 561186 157488
rect 786 142528 561106 142808
rect 786 140088 561186 142528
rect 866 139808 561186 140088
rect 786 125128 561186 139808
rect 786 124848 561106 125128
rect 786 122408 561186 124848
rect 866 122128 561186 122408
rect 786 107448 561186 122128
rect 786 107168 561106 107448
rect 786 104728 561186 107168
rect 866 104448 561186 104728
rect 786 89768 561186 104448
rect 786 89488 561106 89768
rect 786 87048 561186 89488
rect 866 86768 561186 87048
rect 786 72768 561186 86768
rect 786 72488 561106 72768
rect 786 70048 561186 72488
rect 866 69768 561186 70048
rect 786 55088 561186 69768
rect 786 54808 561106 55088
rect 786 52368 561186 54808
rect 866 52088 561186 52368
rect 786 37408 561186 52088
rect 786 37128 561106 37408
rect 786 34688 561186 37128
rect 866 34408 561186 34688
rect 786 19728 561186 34408
rect 786 19448 561106 19728
rect 786 17008 561186 19448
rect 866 16728 561186 17008
rect 786 2048 561186 16728
rect 786 1768 561106 2048
rect 786 1739 561186 1768
<< metal4 >>
rect 2494 411016 2814 456808
rect 3230 411016 3550 456808
rect 2494 308744 2814 354536
rect 3230 308744 3550 354536
rect 2494 207016 2814 252808
rect 3230 207016 3550 252808
rect 2494 104744 2814 150536
rect 3230 104744 3550 150536
rect 8330 1928 8650 587368
rect 8990 1928 9310 587368
rect 22330 1928 22650 587368
rect 22990 1928 23310 587368
rect 36330 98409 36650 587368
rect 36990 98409 37310 587368
rect 50330 98409 50650 587368
rect 50990 98409 51310 587368
rect 64330 449649 64650 587368
rect 64990 449649 65310 587368
rect 78330 449649 78650 587368
rect 78990 449649 79310 587368
rect 64330 353225 64650 430231
rect 64990 353225 65310 430231
rect 78330 353225 78650 430231
rect 78990 353225 79310 430231
rect 64330 251225 64650 314903
rect 64990 251225 65310 314903
rect 78330 251225 78650 314903
rect 78990 251225 79310 314903
rect 64330 149225 64650 212903
rect 64990 149225 65310 212903
rect 78330 149225 78650 212903
rect 78990 149225 79310 212903
rect 36330 1928 36650 60495
rect 36990 1928 37310 60495
rect 50330 1928 50650 60495
rect 50990 1928 51310 60495
rect 64330 1928 64650 110903
rect 64990 1928 65310 110903
rect 78330 1928 78650 110903
rect 78990 1928 79310 110903
rect 92330 1928 92650 587368
rect 92990 455444 93310 587368
rect 106330 509252 106650 587368
rect 106990 503865 107310 587368
rect 120330 503865 120650 587368
rect 120990 503865 121310 587368
rect 134330 503865 134650 587368
rect 134990 503865 135310 587368
rect 92990 353444 93310 415868
rect 100934 413192 101254 458440
rect 101670 413192 101990 458440
rect 106330 407252 106650 465868
rect 106990 401865 107310 466767
rect 120330 454953 120650 466767
rect 120990 454953 121310 466767
rect 134330 454953 134650 466767
rect 120330 401865 120650 416087
rect 120990 401865 121310 416087
rect 134330 401865 134650 416087
rect 134990 401865 135310 466767
rect 92990 251444 93310 313868
rect 100934 310920 101254 356712
rect 101670 310920 101990 356712
rect 106330 305252 106650 363868
rect 106990 299865 107310 364767
rect 120330 299865 120650 364767
rect 120990 299865 121310 364767
rect 134330 299865 134650 364767
rect 134990 299865 135310 364767
rect 92990 149444 93310 211868
rect 102406 209192 102726 254440
rect 103142 209192 103462 254440
rect 106330 203252 106650 261868
rect 106990 197865 107310 262767
rect 120330 197865 120650 262767
rect 120990 197865 121310 262767
rect 134330 224977 134650 262767
rect 134330 197865 134650 212903
rect 134990 197865 135310 262767
rect 92990 1928 93310 109868
rect 100934 106920 101254 152712
rect 101670 106920 101990 152712
rect 106330 1928 106650 159868
rect 106990 1928 107310 160767
rect 120330 1928 120650 160767
rect 120990 1928 121310 160767
rect 134330 1928 134650 160767
rect 134990 1928 135310 160767
rect 148330 1928 148650 587368
rect 148990 1928 149310 587368
rect 162330 448929 162650 587368
rect 162990 448929 163310 587368
rect 176330 448929 176650 587368
rect 176990 448929 177310 587368
rect 162330 350465 162650 418359
rect 162990 350465 163310 418359
rect 176330 350465 176650 418359
rect 176990 350465 177310 418359
rect 190330 350465 190650 587368
rect 190990 505444 191310 587368
rect 190990 457444 191310 465868
rect 199558 462696 199878 508488
rect 200294 462696 200614 508488
rect 204330 503865 204650 587368
rect 204990 503865 205310 587368
rect 218330 503865 218650 587368
rect 218990 503865 219310 587368
rect 232330 503865 232650 587368
rect 232990 503865 233310 587368
rect 190990 403444 191310 417868
rect 201398 415368 201718 457896
rect 190990 355444 191310 363868
rect 199558 360968 199878 406760
rect 200294 360968 200614 406760
rect 204330 401865 204650 466767
rect 204990 401865 205310 466767
rect 218330 401865 218650 466767
rect 218990 401865 219310 466767
rect 232330 454953 232650 466767
rect 232990 454953 233310 466767
rect 232330 401865 232650 416087
rect 232990 401865 233310 416087
rect 162330 248465 162650 316087
rect 162990 248465 163310 316087
rect 176330 248465 176650 316087
rect 176990 248465 177310 316087
rect 190330 248465 190650 316087
rect 190990 301444 191310 315868
rect 201398 313096 201718 356712
rect 190990 253444 191310 261868
rect 199558 258696 199878 304488
rect 200294 258696 200614 304488
rect 204330 299865 204650 364767
rect 204990 299865 205310 364767
rect 218330 299865 218650 364767
rect 218990 299865 219310 364767
rect 232330 326977 232650 364767
rect 232990 326977 233310 364767
rect 232330 299865 232650 314903
rect 232990 299865 233310 314903
rect 162330 146465 162650 214087
rect 162990 146465 163310 214087
rect 176330 146465 176650 214087
rect 176990 146465 177310 214087
rect 190330 146465 190650 214087
rect 190990 199444 191310 213868
rect 201398 210824 201718 254440
rect 190990 151444 191310 159868
rect 199558 156968 199878 202760
rect 200294 156968 200614 202760
rect 204330 197865 204650 262767
rect 204990 197865 205310 262767
rect 218330 197865 218650 262767
rect 218990 197865 219310 262767
rect 232330 224977 232650 262767
rect 232990 224977 233310 262767
rect 232330 197865 232650 212903
rect 232990 197865 233310 212903
rect 162330 96505 162650 112087
rect 162990 96505 163310 112087
rect 176330 96505 176650 112087
rect 176990 96505 177310 112087
rect 162330 1928 162650 67159
rect 162990 1928 163310 67159
rect 176330 1928 176650 67159
rect 176990 1928 177310 67159
rect 190330 1928 190650 112087
rect 190990 99444 191310 111868
rect 201398 109640 201718 152168
rect 190990 1928 191310 59868
rect 201398 57416 201718 98856
rect 204330 1928 204650 160767
rect 204990 1928 205310 160767
rect 218330 1928 218650 160767
rect 218990 1928 219310 160767
rect 232330 122977 232650 160767
rect 232990 122977 233310 160767
rect 232330 75505 232650 110903
rect 232330 1928 232650 56223
rect 232990 1928 233310 110903
rect 246330 1928 246650 587368
rect 246990 1928 247310 587368
rect 252550 462696 252870 508488
rect 253286 462696 253606 508488
rect 251262 414824 251582 458440
rect 260330 448929 260650 587368
rect 260990 448929 261310 587368
rect 274330 448929 274650 587368
rect 274990 448929 275310 587368
rect 252550 360968 252870 406760
rect 253286 360968 253606 406760
rect 251262 313640 251582 356168
rect 260330 350465 260650 418359
rect 260990 350465 261310 418359
rect 274330 350465 274650 418359
rect 274990 350465 275310 418359
rect 288330 350465 288650 587368
rect 288990 350465 289310 587368
rect 252550 258696 252870 304488
rect 253286 258696 253606 304488
rect 251262 211368 251582 253896
rect 260330 248465 260650 316087
rect 260990 248465 261310 316087
rect 274330 248465 274650 316087
rect 274990 248465 275310 316087
rect 288330 248465 288650 316087
rect 288990 248465 289310 316087
rect 252550 156968 252870 202760
rect 253286 156968 253606 202760
rect 251262 109096 251582 152712
rect 260330 146465 260650 214087
rect 260990 146465 261310 214087
rect 274330 146465 274650 214087
rect 274990 146465 275310 214087
rect 288330 146465 288650 214087
rect 288990 146465 289310 214087
rect 251998 56872 252318 98856
rect 252734 56872 253054 98856
rect 260330 96505 260650 112087
rect 260990 96505 261310 112087
rect 274330 96505 274650 112087
rect 274990 96505 275310 112087
rect 260330 1928 260650 67159
rect 260990 1928 261310 67159
rect 274330 1928 274650 67159
rect 274990 1928 275310 67159
rect 288330 1928 288650 112087
rect 288990 1928 289310 112087
rect 302330 1928 302650 587368
rect 302990 1928 303310 587368
rect 316330 503865 316650 587368
rect 316990 561444 317310 587368
rect 316990 503865 317310 521868
rect 330330 503865 330650 587368
rect 330990 503865 331310 587368
rect 344330 503865 344650 587368
rect 344990 503865 345310 587368
rect 316330 401865 316650 466767
rect 316990 401865 317310 466767
rect 330330 454953 330650 466767
rect 330990 454953 331310 466767
rect 330330 401865 330650 416087
rect 330990 401865 331310 416087
rect 344330 401865 344650 466767
rect 344990 401865 345310 466767
rect 354486 462696 354806 508488
rect 355222 462696 355542 508488
rect 353014 414824 353334 458440
rect 353750 414824 354070 458440
rect 316330 299865 316650 364767
rect 316990 299865 317310 364767
rect 330330 299865 330650 364767
rect 330990 299865 331310 364767
rect 344330 299865 344650 364767
rect 344990 299865 345310 364767
rect 354486 360968 354806 406760
rect 355222 360968 355542 406760
rect 353014 313096 353334 356712
rect 353750 313096 354070 356712
rect 316330 197865 316650 262767
rect 316990 197865 317310 262767
rect 330330 197865 330650 262767
rect 330990 197865 331310 262767
rect 344330 197865 344650 262767
rect 344990 197865 345310 262767
rect 354486 258696 354806 304488
rect 355222 258696 355542 304488
rect 353014 210824 353334 254440
rect 353750 210824 354070 254440
rect 316330 1928 316650 160767
rect 316990 45444 317310 160767
rect 330330 75505 330650 160767
rect 330990 75505 331310 160767
rect 316990 1928 317310 5868
rect 330330 1928 330650 56223
rect 330990 1928 331310 56223
rect 344330 1928 344650 160767
rect 344990 1928 345310 160767
rect 354486 156968 354806 202760
rect 355222 156968 355542 202760
rect 353014 109096 353334 154888
rect 353750 109096 354070 154888
rect 353934 56872 354254 98856
rect 354670 56872 354990 98856
rect 358330 1928 358650 587368
rect 358990 448929 359310 587368
rect 372330 448929 372650 587368
rect 372990 448929 373310 587368
rect 386330 491489 386650 587368
rect 386990 491489 387310 587368
rect 358990 1928 359310 418359
rect 372330 350465 372650 418359
rect 372990 350465 373310 418359
rect 386330 389489 386650 471255
rect 386990 389489 387310 471255
rect 386330 350465 386650 369255
rect 386990 350465 387310 369255
rect 372330 248465 372650 316087
rect 372990 248465 373310 316087
rect 386330 287489 386650 316087
rect 386990 287489 387310 316087
rect 386330 248465 386650 267255
rect 386990 248465 387310 267255
rect 372330 146465 372650 214087
rect 372990 146465 373310 214087
rect 386330 185489 386650 214087
rect 386990 185489 387310 214087
rect 386330 146465 386650 165255
rect 386990 146465 387310 165255
rect 372330 96505 372650 112087
rect 372990 96505 373310 112087
rect 386330 96505 386650 112087
rect 386990 96505 387310 112087
rect 372330 1928 372650 67159
rect 372990 1928 373310 67159
rect 386330 1928 386650 67159
rect 386990 1928 387310 67159
rect 400330 1928 400650 587368
rect 400990 1928 401310 587368
rect 403430 466660 403750 508488
rect 403430 462696 403750 466600
rect 404166 466660 404486 508488
rect 414330 503865 414650 587368
rect 414990 503865 415310 587368
rect 428330 503865 428650 587368
rect 428990 503865 429310 587368
rect 442330 503865 442650 587368
rect 442990 509252 443310 587368
rect 404166 462696 404486 466600
rect 404902 414824 405222 458440
rect 405638 414824 405958 458440
rect 403430 364932 403750 406760
rect 403430 360968 403750 364872
rect 404166 364932 404486 406760
rect 414330 401865 414650 466767
rect 414990 455444 415310 466767
rect 428330 454953 428650 466767
rect 428990 454953 429310 466767
rect 414990 401865 415310 415868
rect 428330 401865 428650 416087
rect 428990 401865 429310 416087
rect 442330 401865 442650 466767
rect 442990 407252 443310 465868
rect 404166 360968 404486 364872
rect 404902 313096 405222 356712
rect 405638 313096 405958 356712
rect 403430 262660 403750 304488
rect 403430 258696 403750 262600
rect 404166 262660 404486 304488
rect 414330 299865 414650 364767
rect 414990 353444 415310 364767
rect 414990 299865 415310 313868
rect 428330 299865 428650 364767
rect 428990 299865 429310 364767
rect 442330 299865 442650 364767
rect 442990 305252 443310 363868
rect 404166 258696 404486 262600
rect 404902 210824 405222 255528
rect 405638 210824 405958 255528
rect 403430 160932 403750 202760
rect 403430 156968 403750 160872
rect 404166 160932 404486 202760
rect 414330 197865 414650 262767
rect 414990 252044 415310 262767
rect 414990 197865 415310 212468
rect 428330 197865 428650 262767
rect 428990 197865 429310 262767
rect 442330 197865 442650 262767
rect 442990 203252 443310 261868
rect 404166 156968 404486 160872
rect 404902 109096 405222 152712
rect 405638 109096 405958 152712
rect 404902 56872 405222 98856
rect 405638 56872 405958 98856
rect 414330 1928 414650 160767
rect 414990 149444 415310 160767
rect 414990 95444 415310 109868
rect 428330 75505 428650 160767
rect 428990 75505 429310 160767
rect 414990 1928 415310 55868
rect 428330 1928 428650 56223
rect 428990 1928 429310 56223
rect 442330 1928 442650 160767
rect 442990 1928 443310 159868
rect 456330 1928 456650 587368
rect 456990 1928 457310 587368
rect 470330 479729 470650 587368
rect 470990 479729 471310 587368
rect 470330 377729 470650 460855
rect 470990 377729 471310 460855
rect 484330 435257 484650 587368
rect 484990 437652 485310 587368
rect 470330 343865 470650 358855
rect 470990 343865 471310 358855
rect 484330 343865 484650 408767
rect 484990 343865 485310 407868
rect 470330 275729 470650 306359
rect 470990 275729 471310 306359
rect 470330 241865 470650 256855
rect 470990 241865 471310 256855
rect 484330 241865 484650 306359
rect 484990 241865 485310 306359
rect 470330 173729 470650 204359
rect 470990 173729 471310 204359
rect 470330 145865 470650 154855
rect 470990 145865 471310 154855
rect 484330 145865 484650 204359
rect 484990 145865 485310 204359
rect 470330 98545 470650 108359
rect 470990 98545 471310 108359
rect 484330 98545 484650 108359
rect 484990 98545 485310 108359
rect 470330 1928 470650 61719
rect 470990 1928 471310 61719
rect 484330 1928 484650 61719
rect 484990 1928 485310 61719
rect 498330 1928 498650 587368
rect 498990 437652 499310 587368
rect 506470 458888 506790 501416
rect 507206 458888 507526 501416
rect 498990 1928 499310 407868
rect 506470 357160 506790 399688
rect 507206 357160 507526 399688
rect 506470 254888 506790 297416
rect 507206 254888 507526 297416
rect 506470 153160 506790 195688
rect 507206 153160 507526 195688
rect 512330 1928 512650 587368
rect 512990 1928 513310 587368
rect 526330 1928 526650 587368
rect 526990 1928 527310 587368
rect 540330 1928 540650 587368
rect 540990 1928 541310 587368
rect 554330 1928 554650 587368
rect 554990 1928 555310 587368
rect 557990 458888 558310 504680
rect 558726 458888 559046 504680
rect 557990 357160 558310 402408
rect 558726 357160 559046 402408
rect 557990 254888 558310 300680
rect 558726 254888 559046 300680
rect 557990 153160 558310 198408
rect 558726 153160 559046 198408
<< obsm4 >>
rect 5381 1848 8250 587149
rect 8730 1848 8910 587149
rect 9390 1848 22250 587149
rect 22730 1848 22910 587149
rect 23390 98329 36250 587149
rect 36730 98329 36910 587149
rect 37390 98329 50250 587149
rect 50730 98329 50910 587149
rect 51390 449569 64250 587149
rect 64730 449569 64910 587149
rect 65390 449569 78250 587149
rect 78730 449569 78910 587149
rect 79390 449569 92250 587149
rect 51390 430311 92250 449569
rect 51390 353145 64250 430311
rect 64730 353145 64910 430311
rect 65390 353145 78250 430311
rect 78730 353145 78910 430311
rect 79390 353145 92250 430311
rect 51390 314983 92250 353145
rect 51390 251145 64250 314983
rect 64730 251145 64910 314983
rect 65390 251145 78250 314983
rect 78730 251145 78910 314983
rect 79390 251145 92250 314983
rect 51390 212983 92250 251145
rect 51390 149145 64250 212983
rect 64730 149145 64910 212983
rect 65390 149145 78250 212983
rect 78730 149145 78910 212983
rect 79390 149145 92250 212983
rect 51390 110983 92250 149145
rect 51390 98329 64250 110983
rect 23390 60575 64250 98329
rect 23390 1848 36250 60575
rect 36730 1848 36910 60575
rect 37390 1848 50250 60575
rect 50730 1848 50910 60575
rect 51390 1848 64250 60575
rect 64730 1848 64910 110983
rect 65390 1848 78250 110983
rect 78730 1848 78910 110983
rect 79390 1848 92250 110983
rect 92730 455364 92910 587149
rect 93390 509172 106250 587149
rect 106730 509172 106910 587149
rect 93390 503785 106910 509172
rect 107390 503785 120250 587149
rect 120730 503785 120910 587149
rect 121390 503785 134250 587149
rect 134730 503785 134910 587149
rect 135390 503785 148250 587149
rect 93390 466847 148250 503785
rect 93390 465948 106910 466847
rect 93390 458520 106250 465948
rect 93390 455364 100854 458520
rect 92730 415948 100854 455364
rect 92730 353364 92910 415948
rect 93390 413112 100854 415948
rect 101334 413112 101590 458520
rect 102070 413112 106250 458520
rect 93390 407172 106250 413112
rect 106730 407172 106910 465948
rect 93390 401785 106910 407172
rect 107390 454873 120250 466847
rect 120730 454873 120910 466847
rect 121390 454873 134250 466847
rect 134730 454873 134910 466847
rect 107390 416167 134910 454873
rect 107390 401785 120250 416167
rect 120730 401785 120910 416167
rect 121390 401785 134250 416167
rect 134730 401785 134910 416167
rect 135390 401785 148250 466847
rect 93390 364847 148250 401785
rect 93390 363948 106910 364847
rect 93390 356792 106250 363948
rect 93390 353364 100854 356792
rect 92730 313948 100854 353364
rect 92730 251364 92910 313948
rect 93390 310840 100854 313948
rect 101334 310840 101590 356792
rect 102070 310840 106250 356792
rect 93390 305172 106250 310840
rect 106730 305172 106910 363948
rect 93390 299785 106910 305172
rect 107390 299785 120250 364847
rect 120730 299785 120910 364847
rect 121390 299785 134250 364847
rect 134730 299785 134910 364847
rect 135390 299785 148250 364847
rect 93390 262847 148250 299785
rect 93390 261948 106910 262847
rect 93390 254520 106250 261948
rect 93390 251364 102326 254520
rect 92730 211948 102326 251364
rect 92730 149364 92910 211948
rect 93390 209112 102326 211948
rect 102806 209112 103062 254520
rect 103542 209112 106250 254520
rect 93390 203172 106250 209112
rect 106730 203172 106910 261948
rect 93390 197785 106910 203172
rect 107390 197785 120250 262847
rect 120730 197785 120910 262847
rect 121390 224897 134250 262847
rect 134730 224897 134910 262847
rect 121390 212983 134910 224897
rect 121390 197785 134250 212983
rect 134730 197785 134910 212983
rect 135390 197785 148250 262847
rect 93390 160847 148250 197785
rect 93390 159948 106910 160847
rect 93390 152792 106250 159948
rect 93390 149364 100854 152792
rect 92730 109948 100854 149364
rect 92730 1848 92910 109948
rect 93390 106840 100854 109948
rect 101334 106840 101590 152792
rect 102070 106840 106250 152792
rect 93390 1848 106250 106840
rect 106730 1848 106910 159948
rect 107390 1848 120250 160847
rect 120730 1848 120910 160847
rect 121390 1848 134250 160847
rect 134730 1848 134910 160847
rect 135390 1848 148250 160847
rect 148730 1848 148910 587149
rect 149390 448849 162250 587149
rect 162730 448849 162910 587149
rect 163390 448849 176250 587149
rect 176730 448849 176910 587149
rect 177390 448849 190250 587149
rect 149390 418439 190250 448849
rect 149390 350385 162250 418439
rect 162730 350385 162910 418439
rect 163390 350385 176250 418439
rect 176730 350385 176910 418439
rect 177390 350385 190250 418439
rect 190730 505364 190910 587149
rect 191390 508568 204250 587149
rect 191390 505364 199478 508568
rect 190730 465948 199478 505364
rect 190730 457364 190910 465948
rect 191390 462616 199478 465948
rect 199958 462616 200214 508568
rect 200694 503785 204250 508568
rect 204730 503785 204910 587149
rect 205390 503785 218250 587149
rect 218730 503785 218910 587149
rect 219390 503785 232250 587149
rect 232730 503785 232910 587149
rect 233390 503785 246250 587149
rect 200694 466847 246250 503785
rect 200694 462616 204250 466847
rect 191390 457976 204250 462616
rect 191390 457364 201318 457976
rect 190730 417948 201318 457364
rect 190730 403364 190910 417948
rect 191390 415288 201318 417948
rect 201798 415288 204250 457976
rect 191390 406840 204250 415288
rect 191390 403364 199478 406840
rect 190730 363948 199478 403364
rect 190730 355364 190910 363948
rect 191390 360888 199478 363948
rect 199958 360888 200214 406840
rect 200694 401785 204250 406840
rect 204730 401785 204910 466847
rect 205390 401785 218250 466847
rect 218730 401785 218910 466847
rect 219390 454873 232250 466847
rect 232730 454873 232910 466847
rect 233390 454873 246250 466847
rect 219390 416167 246250 454873
rect 219390 401785 232250 416167
rect 232730 401785 232910 416167
rect 233390 401785 246250 416167
rect 200694 364847 246250 401785
rect 200694 360888 204250 364847
rect 191390 356792 204250 360888
rect 191390 355364 201318 356792
rect 190730 350385 201318 355364
rect 149390 316167 201318 350385
rect 149390 248385 162250 316167
rect 162730 248385 162910 316167
rect 163390 248385 176250 316167
rect 176730 248385 176910 316167
rect 177390 248385 190250 316167
rect 190730 315948 201318 316167
rect 190730 301364 190910 315948
rect 191390 313016 201318 315948
rect 201798 313016 204250 356792
rect 191390 304568 204250 313016
rect 191390 301364 199478 304568
rect 190730 261948 199478 301364
rect 190730 253364 190910 261948
rect 191390 258616 199478 261948
rect 199958 258616 200214 304568
rect 200694 299785 204250 304568
rect 204730 299785 204910 364847
rect 205390 299785 218250 364847
rect 218730 299785 218910 364847
rect 219390 326897 232250 364847
rect 232730 326897 232910 364847
rect 233390 326897 246250 364847
rect 219390 314983 246250 326897
rect 219390 299785 232250 314983
rect 232730 299785 232910 314983
rect 233390 299785 246250 314983
rect 200694 262847 246250 299785
rect 200694 258616 204250 262847
rect 191390 254520 204250 258616
rect 191390 253364 201318 254520
rect 190730 248385 201318 253364
rect 149390 214167 201318 248385
rect 149390 146385 162250 214167
rect 162730 146385 162910 214167
rect 163390 146385 176250 214167
rect 176730 146385 176910 214167
rect 177390 146385 190250 214167
rect 190730 213948 201318 214167
rect 190730 199364 190910 213948
rect 191390 210744 201318 213948
rect 201798 210744 204250 254520
rect 191390 202840 204250 210744
rect 191390 199364 199478 202840
rect 190730 159948 199478 199364
rect 190730 151364 190910 159948
rect 191390 156888 199478 159948
rect 199958 156888 200214 202840
rect 200694 197785 204250 202840
rect 204730 197785 204910 262847
rect 205390 197785 218250 262847
rect 218730 197785 218910 262847
rect 219390 224897 232250 262847
rect 232730 224897 232910 262847
rect 233390 224897 246250 262847
rect 219390 212983 246250 224897
rect 219390 197785 232250 212983
rect 232730 197785 232910 212983
rect 233390 197785 246250 212983
rect 200694 160847 246250 197785
rect 200694 156888 204250 160847
rect 191390 152248 204250 156888
rect 191390 151364 201318 152248
rect 190730 146385 201318 151364
rect 149390 112167 201318 146385
rect 149390 96425 162250 112167
rect 162730 96425 162910 112167
rect 163390 96425 176250 112167
rect 176730 96425 176910 112167
rect 177390 96425 190250 112167
rect 149390 67239 190250 96425
rect 149390 1848 162250 67239
rect 162730 1848 162910 67239
rect 163390 1848 176250 67239
rect 176730 1848 176910 67239
rect 177390 1848 190250 67239
rect 190730 111948 201318 112167
rect 190730 99364 190910 111948
rect 191390 109560 201318 111948
rect 201798 109560 204250 152248
rect 191390 99364 204250 109560
rect 190730 98936 204250 99364
rect 190730 59948 201318 98936
rect 190730 1848 190910 59948
rect 191390 57336 201318 59948
rect 201798 57336 204250 98936
rect 191390 1848 204250 57336
rect 204730 1848 204910 160847
rect 205390 1848 218250 160847
rect 218730 1848 218910 160847
rect 219390 122897 232250 160847
rect 232730 122897 232910 160847
rect 233390 122897 246250 160847
rect 219390 110983 246250 122897
rect 219390 75425 232250 110983
rect 232730 75425 232910 110983
rect 219390 56303 232910 75425
rect 219390 1848 232250 56303
rect 232730 1848 232910 56303
rect 233390 1848 246250 110983
rect 246730 1848 246910 587149
rect 247390 508568 260250 587149
rect 247390 462616 252470 508568
rect 252950 462616 253206 508568
rect 253686 462616 260250 508568
rect 247390 458520 260250 462616
rect 247390 414744 251182 458520
rect 251662 448849 260250 458520
rect 260730 448849 260910 587149
rect 261390 448849 274250 587149
rect 274730 448849 274910 587149
rect 275390 448849 288250 587149
rect 251662 418439 288250 448849
rect 251662 414744 260250 418439
rect 247390 406840 260250 414744
rect 247390 360888 252470 406840
rect 252950 360888 253206 406840
rect 253686 360888 260250 406840
rect 247390 356248 260250 360888
rect 247390 313560 251182 356248
rect 251662 350385 260250 356248
rect 260730 350385 260910 418439
rect 261390 350385 274250 418439
rect 274730 350385 274910 418439
rect 275390 350385 288250 418439
rect 288730 350385 288910 587149
rect 289390 350385 302250 587149
rect 251662 316167 302250 350385
rect 251662 313560 260250 316167
rect 247390 304568 260250 313560
rect 247390 258616 252470 304568
rect 252950 258616 253206 304568
rect 253686 258616 260250 304568
rect 247390 253976 260250 258616
rect 247390 211288 251182 253976
rect 251662 248385 260250 253976
rect 260730 248385 260910 316167
rect 261390 248385 274250 316167
rect 274730 248385 274910 316167
rect 275390 248385 288250 316167
rect 288730 248385 288910 316167
rect 289390 248385 302250 316167
rect 251662 214167 302250 248385
rect 251662 211288 260250 214167
rect 247390 202840 260250 211288
rect 247390 156888 252470 202840
rect 252950 156888 253206 202840
rect 253686 156888 260250 202840
rect 247390 152792 260250 156888
rect 247390 109016 251182 152792
rect 251662 146385 260250 152792
rect 260730 146385 260910 214167
rect 261390 146385 274250 214167
rect 274730 146385 274910 214167
rect 275390 146385 288250 214167
rect 288730 146385 288910 214167
rect 289390 146385 302250 214167
rect 251662 112167 302250 146385
rect 251662 109016 260250 112167
rect 247390 98936 260250 109016
rect 247390 56792 251918 98936
rect 252398 56792 252654 98936
rect 253134 96425 260250 98936
rect 260730 96425 260910 112167
rect 261390 96425 274250 112167
rect 274730 96425 274910 112167
rect 275390 96425 288250 112167
rect 253134 67239 288250 96425
rect 253134 56792 260250 67239
rect 247390 1848 260250 56792
rect 260730 1848 260910 67239
rect 261390 1848 274250 67239
rect 274730 1848 274910 67239
rect 275390 1848 288250 67239
rect 288730 1848 288910 112167
rect 289390 1848 302250 112167
rect 302730 1848 302910 587149
rect 303390 503785 316250 587149
rect 316730 561364 316910 587149
rect 317390 561364 330250 587149
rect 316730 521948 330250 561364
rect 316730 503785 316910 521948
rect 317390 503785 330250 521948
rect 330730 503785 330910 587149
rect 331390 503785 344250 587149
rect 344730 503785 344910 587149
rect 345390 508568 358250 587149
rect 345390 503785 354406 508568
rect 303390 466847 354406 503785
rect 303390 401785 316250 466847
rect 316730 401785 316910 466847
rect 317390 454873 330250 466847
rect 330730 454873 330910 466847
rect 331390 454873 344250 466847
rect 317390 416167 344250 454873
rect 317390 401785 330250 416167
rect 330730 401785 330910 416167
rect 331390 401785 344250 416167
rect 344730 401785 344910 466847
rect 345390 462616 354406 466847
rect 354886 462616 355142 508568
rect 355622 462616 358250 508568
rect 345390 458520 358250 462616
rect 345390 414744 352934 458520
rect 353414 414744 353670 458520
rect 354150 414744 358250 458520
rect 345390 406840 358250 414744
rect 345390 401785 354406 406840
rect 303390 364847 354406 401785
rect 303390 299785 316250 364847
rect 316730 299785 316910 364847
rect 317390 299785 330250 364847
rect 330730 299785 330910 364847
rect 331390 299785 344250 364847
rect 344730 299785 344910 364847
rect 345390 360888 354406 364847
rect 354886 360888 355142 406840
rect 355622 360888 358250 406840
rect 345390 356792 358250 360888
rect 345390 313016 352934 356792
rect 353414 313016 353670 356792
rect 354150 313016 358250 356792
rect 345390 304568 358250 313016
rect 345390 299785 354406 304568
rect 303390 262847 354406 299785
rect 303390 197785 316250 262847
rect 316730 197785 316910 262847
rect 317390 197785 330250 262847
rect 330730 197785 330910 262847
rect 331390 197785 344250 262847
rect 344730 197785 344910 262847
rect 345390 258616 354406 262847
rect 354886 258616 355142 304568
rect 355622 258616 358250 304568
rect 345390 254520 358250 258616
rect 345390 210744 352934 254520
rect 353414 210744 353670 254520
rect 354150 210744 358250 254520
rect 345390 202840 358250 210744
rect 345390 197785 354406 202840
rect 303390 160847 354406 197785
rect 303390 1848 316250 160847
rect 316730 45364 316910 160847
rect 317390 75425 330250 160847
rect 330730 75425 330910 160847
rect 331390 75425 344250 160847
rect 317390 56303 344250 75425
rect 317390 45364 330250 56303
rect 316730 5948 330250 45364
rect 316730 1848 316910 5948
rect 317390 1848 330250 5948
rect 330730 1848 330910 56303
rect 331390 1848 344250 56303
rect 344730 1848 344910 160847
rect 345390 156888 354406 160847
rect 354886 156888 355142 202840
rect 355622 156888 358250 202840
rect 345390 154968 358250 156888
rect 345390 109016 352934 154968
rect 353414 109016 353670 154968
rect 354150 109016 358250 154968
rect 345390 98936 358250 109016
rect 345390 56792 353854 98936
rect 354334 56792 354590 98936
rect 355070 56792 358250 98936
rect 345390 1848 358250 56792
rect 358730 448849 358910 587149
rect 359390 448849 372250 587149
rect 372730 448849 372910 587149
rect 373390 491409 386250 587149
rect 386730 491409 386910 587149
rect 387390 491409 400250 587149
rect 373390 471335 400250 491409
rect 373390 448849 386250 471335
rect 358730 418439 386250 448849
rect 358730 1848 358910 418439
rect 359390 350385 372250 418439
rect 372730 350385 372910 418439
rect 373390 389409 386250 418439
rect 386730 389409 386910 471335
rect 387390 389409 400250 471335
rect 373390 369335 400250 389409
rect 373390 350385 386250 369335
rect 386730 350385 386910 369335
rect 387390 350385 400250 369335
rect 359390 316167 400250 350385
rect 359390 248385 372250 316167
rect 372730 248385 372910 316167
rect 373390 287409 386250 316167
rect 386730 287409 386910 316167
rect 387390 287409 400250 316167
rect 373390 267335 400250 287409
rect 373390 248385 386250 267335
rect 386730 248385 386910 267335
rect 387390 248385 400250 267335
rect 359390 214167 400250 248385
rect 359390 146385 372250 214167
rect 372730 146385 372910 214167
rect 373390 185409 386250 214167
rect 386730 185409 386910 214167
rect 387390 185409 400250 214167
rect 373390 165335 400250 185409
rect 373390 146385 386250 165335
rect 386730 146385 386910 165335
rect 387390 146385 400250 165335
rect 359390 112167 400250 146385
rect 359390 96425 372250 112167
rect 372730 96425 372910 112167
rect 373390 96425 386250 112167
rect 386730 96425 386910 112167
rect 387390 96425 400250 112167
rect 359390 67239 400250 96425
rect 359390 1848 372250 67239
rect 372730 1848 372910 67239
rect 373390 1848 386250 67239
rect 386730 1848 386910 67239
rect 387390 1848 400250 67239
rect 400730 1848 400910 587149
rect 401390 508568 414250 587149
rect 401390 462616 403350 508568
rect 403830 462616 404086 508568
rect 404566 503785 414250 508568
rect 414730 503785 414910 587149
rect 415390 503785 428250 587149
rect 428730 503785 428910 587149
rect 429390 503785 442250 587149
rect 442730 509172 442910 587149
rect 443390 509172 456250 587149
rect 442730 503785 456250 509172
rect 404566 466847 456250 503785
rect 404566 462616 414250 466847
rect 401390 458520 414250 462616
rect 401390 414744 404822 458520
rect 405302 414744 405558 458520
rect 406038 414744 414250 458520
rect 401390 406840 414250 414744
rect 401390 360888 403350 406840
rect 403830 360888 404086 406840
rect 404566 401785 414250 406840
rect 414730 455364 414910 466847
rect 415390 455364 428250 466847
rect 414730 454873 428250 455364
rect 428730 454873 428910 466847
rect 429390 454873 442250 466847
rect 414730 416167 442250 454873
rect 414730 415948 428250 416167
rect 414730 401785 414910 415948
rect 415390 401785 428250 415948
rect 428730 401785 428910 416167
rect 429390 401785 442250 416167
rect 442730 465948 456250 466847
rect 442730 407172 442910 465948
rect 443390 407172 456250 465948
rect 442730 401785 456250 407172
rect 404566 364847 456250 401785
rect 404566 360888 414250 364847
rect 401390 356792 414250 360888
rect 401390 313016 404822 356792
rect 405302 313016 405558 356792
rect 406038 313016 414250 356792
rect 401390 304568 414250 313016
rect 401390 258616 403350 304568
rect 403830 258616 404086 304568
rect 404566 299785 414250 304568
rect 414730 353364 414910 364847
rect 415390 353364 428250 364847
rect 414730 313948 428250 353364
rect 414730 299785 414910 313948
rect 415390 299785 428250 313948
rect 428730 299785 428910 364847
rect 429390 299785 442250 364847
rect 442730 363948 456250 364847
rect 442730 305172 442910 363948
rect 443390 305172 456250 363948
rect 442730 299785 456250 305172
rect 404566 262847 456250 299785
rect 404566 258616 414250 262847
rect 401390 255608 414250 258616
rect 401390 210744 404822 255608
rect 405302 210744 405558 255608
rect 406038 210744 414250 255608
rect 401390 202840 414250 210744
rect 401390 156888 403350 202840
rect 403830 156888 404086 202840
rect 404566 197785 414250 202840
rect 414730 251964 414910 262847
rect 415390 251964 428250 262847
rect 414730 212548 428250 251964
rect 414730 197785 414910 212548
rect 415390 197785 428250 212548
rect 428730 197785 428910 262847
rect 429390 197785 442250 262847
rect 442730 261948 456250 262847
rect 442730 203172 442910 261948
rect 443390 203172 456250 261948
rect 442730 197785 456250 203172
rect 404566 160847 456250 197785
rect 404566 156888 414250 160847
rect 401390 152792 414250 156888
rect 401390 109016 404822 152792
rect 405302 109016 405558 152792
rect 406038 109016 414250 152792
rect 401390 98936 414250 109016
rect 401390 56792 404822 98936
rect 405302 56792 405558 98936
rect 406038 56792 414250 98936
rect 401390 1848 414250 56792
rect 414730 149364 414910 160847
rect 415390 149364 428250 160847
rect 414730 109948 428250 149364
rect 414730 95364 414910 109948
rect 415390 95364 428250 109948
rect 414730 75425 428250 95364
rect 428730 75425 428910 160847
rect 429390 75425 442250 160847
rect 414730 56303 442250 75425
rect 414730 55948 428250 56303
rect 414730 1848 414910 55948
rect 415390 1848 428250 55948
rect 428730 1848 428910 56303
rect 429390 1848 442250 56303
rect 442730 159948 456250 160847
rect 442730 1848 442910 159948
rect 443390 1848 456250 159948
rect 456730 1848 456910 587149
rect 457390 479649 470250 587149
rect 470730 479649 470910 587149
rect 471390 479649 484250 587149
rect 457390 460935 484250 479649
rect 457390 377649 470250 460935
rect 470730 377649 470910 460935
rect 471390 435177 484250 460935
rect 484730 437572 484910 587149
rect 485390 437572 498250 587149
rect 484730 435177 498250 437572
rect 471390 408847 498250 435177
rect 471390 377649 484250 408847
rect 457390 358935 484250 377649
rect 457390 343785 470250 358935
rect 470730 343785 470910 358935
rect 471390 343785 484250 358935
rect 484730 407948 498250 408847
rect 484730 343785 484910 407948
rect 485390 343785 498250 407948
rect 457390 306439 498250 343785
rect 457390 275649 470250 306439
rect 470730 275649 470910 306439
rect 471390 275649 484250 306439
rect 457390 256935 484250 275649
rect 457390 241785 470250 256935
rect 470730 241785 470910 256935
rect 471390 241785 484250 256935
rect 484730 241785 484910 306439
rect 485390 241785 498250 306439
rect 457390 204439 498250 241785
rect 457390 173649 470250 204439
rect 470730 173649 470910 204439
rect 471390 173649 484250 204439
rect 457390 154935 484250 173649
rect 457390 145785 470250 154935
rect 470730 145785 470910 154935
rect 471390 145785 484250 154935
rect 484730 145785 484910 204439
rect 485390 145785 498250 204439
rect 457390 108439 498250 145785
rect 457390 98465 470250 108439
rect 470730 98465 470910 108439
rect 471390 98465 484250 108439
rect 484730 98465 484910 108439
rect 485390 98465 498250 108439
rect 457390 61799 498250 98465
rect 457390 1848 470250 61799
rect 470730 1848 470910 61799
rect 471390 1848 484250 61799
rect 484730 1848 484910 61799
rect 485390 1848 498250 61799
rect 498730 437572 498910 587149
rect 499390 501496 512250 587149
rect 499390 458808 506390 501496
rect 506870 458808 507126 501496
rect 507606 458808 512250 501496
rect 499390 437572 512250 458808
rect 498730 407948 512250 437572
rect 498730 1848 498910 407948
rect 499390 399768 512250 407948
rect 499390 357080 506390 399768
rect 506870 357080 507126 399768
rect 507606 357080 512250 399768
rect 499390 297496 512250 357080
rect 499390 254808 506390 297496
rect 506870 254808 507126 297496
rect 507606 254808 512250 297496
rect 499390 195768 512250 254808
rect 499390 153080 506390 195768
rect 506870 153080 507126 195768
rect 507606 153080 512250 195768
rect 499390 1848 512250 153080
rect 512730 1848 512910 587149
rect 513390 1848 526250 587149
rect 526730 1848 526910 587149
rect 527390 1848 540250 587149
rect 540730 1848 540910 587149
rect 541390 1848 553399 587149
rect 5381 1739 553399 1848
<< metal5 >>
rect 1042 579876 560866 580196
rect 1042 579216 560866 579536
rect 1042 564876 560866 565196
rect 1042 564216 560866 564536
rect 1042 549876 560866 550196
rect 1042 549216 560866 549536
rect 1042 534876 560866 535196
rect 1042 534216 560866 534536
rect 1042 519876 560866 520196
rect 1042 519216 560866 519536
rect 1042 504876 560866 505196
rect 1042 504216 560866 504536
rect 1042 489876 560866 490196
rect 1042 489216 560866 489536
rect 1042 474876 560866 475196
rect 1042 474216 560866 474536
rect 1042 459876 560866 460196
rect 1042 459216 560866 459536
rect 1042 444876 560866 445196
rect 1042 444216 560866 444536
rect 1042 429876 560866 430196
rect 1042 429216 560866 429536
rect 1042 414876 560866 415196
rect 1042 414216 560866 414536
rect 1042 399876 560866 400196
rect 1042 399216 560866 399536
rect 1042 384876 560866 385196
rect 1042 384216 560866 384536
rect 1042 369876 560866 370196
rect 1042 369216 560866 369536
rect 1042 354876 560866 355196
rect 1042 354216 560866 354536
rect 1042 339876 560866 340196
rect 1042 339216 560866 339536
rect 1042 324876 560866 325196
rect 1042 324216 560866 324536
rect 1042 309876 560866 310196
rect 1042 309216 560866 309536
rect 1042 294876 560866 295196
rect 1042 294216 560866 294536
rect 1042 279876 560866 280196
rect 1042 279216 560866 279536
rect 1042 264876 560866 265196
rect 1042 264216 560866 264536
rect 1042 249876 560866 250196
rect 1042 249216 560866 249536
rect 1042 234876 560866 235196
rect 1042 234216 560866 234536
rect 1042 219876 560866 220196
rect 1042 219216 560866 219536
rect 1042 204876 560866 205196
rect 1042 204216 560866 204536
rect 1042 189876 560866 190196
rect 1042 189216 560866 189536
rect 1042 174876 560866 175196
rect 1042 174216 560866 174536
rect 1042 159876 560866 160196
rect 1042 159216 560866 159536
rect 456330 150260 485310 150580
rect 456330 149580 485310 149900
rect 1042 144876 560866 145196
rect 1042 144216 560866 144536
rect 1042 129876 560866 130196
rect 1042 129216 560866 129536
rect 1042 114876 560866 115196
rect 1042 114216 560866 114536
rect 1042 99876 560866 100196
rect 1042 99216 560866 99536
rect 1042 84876 560866 85196
rect 1042 84216 560866 84536
rect 1042 69876 560866 70196
rect 1042 69216 560866 69536
rect 1042 54876 560866 55196
rect 1042 54216 560866 54536
rect 1042 39876 560866 40196
rect 1042 39216 560866 39536
rect 1042 24876 560866 25196
rect 1042 24216 560866 24536
rect 1042 9876 560866 10196
rect 1042 9216 560866 9536
<< labels >>
rlabel metal2 s 248588 0 248644 600 6 ccff_head
port 1 nsew signal input
rlabel metal2 s 204796 589000 204852 589600 6 ccff_tail
port 2 nsew signal output
rlabel metal2 s 448228 0 448284 600 6 clk
port 3 nsew signal input
rlabel metal2 s 497816 0 497872 600 6 gfpga_pad_GPIO_PAD_in[0]
port 4 nsew signal input
rlabel metal2 s 365152 0 365208 600 6 gfpga_pad_GPIO_PAD_in[10]
port 5 nsew signal input
rlabel metal2 s 254384 589000 254440 589600 6 gfpga_pad_GPIO_PAD_in[11]
port 6 nsew signal input
rlabel metal3 s 561186 19528 561786 19648 6 gfpga_pad_GPIO_PAD_in[12]
port 7 nsew signal input
rlabel metal3 s 561186 510488 561786 510608 6 gfpga_pad_GPIO_PAD_in[13]
port 8 nsew signal input
rlabel metal2 s 553844 589000 553900 589600 6 gfpga_pad_GPIO_PAD_in[14]
port 9 nsew signal input
rlabel metal2 s 337460 589000 337516 589600 6 gfpga_pad_GPIO_PAD_in[15]
port 10 nsew signal input
rlabel metal2 s 149412 0 149468 600 6 gfpga_pad_GPIO_PAD_in[16]
port 11 nsew signal input
rlabel metal3 s 186 122208 786 122328 6 gfpga_pad_GPIO_PAD_in[17]
port 12 nsew signal input
rlabel metal3 s 186 139888 786 140008 6 gfpga_pad_GPIO_PAD_in[18]
port 13 nsew signal input
rlabel metal3 s 186 104528 786 104648 6 gfpga_pad_GPIO_PAD_in[19]
port 14 nsew signal input
rlabel metal2 s 287872 589000 287928 589600 6 gfpga_pad_GPIO_PAD_in[1]
port 15 nsew signal input
rlabel metal2 s 55388 589000 55444 589600 6 gfpga_pad_GPIO_PAD_in[20]
port 16 nsew signal input
rlabel metal3 s 561186 458128 561786 458248 6 gfpga_pad_GPIO_PAD_in[21]
port 17 nsew signal input
rlabel metal3 s 186 420728 786 420848 6 gfpga_pad_GPIO_PAD_in[22]
port 18 nsew signal input
rlabel metal3 s 561186 475808 561786 475928 6 gfpga_pad_GPIO_PAD_in[23]
port 19 nsew signal input
rlabel metal2 s 165512 0 165568 600 6 gfpga_pad_GPIO_PAD_in[24]
port 20 nsew signal input
rlabel metal2 s 520356 589000 520412 589600 6 gfpga_pad_GPIO_PAD_in[25]
port 21 nsew signal input
rlabel metal2 s 370948 589000 371004 589600 6 gfpga_pad_GPIO_PAD_in[26]
port 22 nsew signal input
rlabel metal2 s 72132 589000 72188 589600 6 gfpga_pad_GPIO_PAD_in[27]
port 23 nsew signal input
rlabel metal2 s 271128 589000 271184 589600 6 gfpga_pad_GPIO_PAD_in[28]
port 24 nsew signal input
rlabel metal3 s 186 473088 786 473208 6 gfpga_pad_GPIO_PAD_in[29]
port 25 nsew signal input
rlabel metal3 s 561186 230328 561786 230448 6 gfpga_pad_GPIO_PAD_in[2]
port 26 nsew signal input
rlabel metal3 s 186 333008 786 333128 6 gfpga_pad_GPIO_PAD_in[30]
port 27 nsew signal input
rlabel metal3 s 561186 1848 561786 1968 6 gfpga_pad_GPIO_PAD_in[31]
port 28 nsew signal input
rlabel metal2 s 21900 589000 21956 589600 6 gfpga_pad_GPIO_PAD_in[32]
port 29 nsew signal input
rlabel metal2 s 182256 0 182312 600 6 gfpga_pad_GPIO_PAD_in[33]
port 30 nsew signal input
rlabel metal3 s 561186 248008 561786 248128 6 gfpga_pad_GPIO_PAD_in[34]
port 31 nsew signal input
rlabel metal2 s 232488 0 232544 600 6 gfpga_pad_GPIO_PAD_in[35]
port 32 nsew signal input
rlabel metal3 s 186 245288 786 245408 6 gfpga_pad_GPIO_PAD_in[36]
port 33 nsew signal input
rlabel metal2 s 88232 589000 88288 589600 6 gfpga_pad_GPIO_PAD_in[37]
port 34 nsew signal input
rlabel metal2 s 304616 589000 304672 589600 6 gfpga_pad_GPIO_PAD_in[38]
port 35 nsew signal input
rlabel metal2 s 470768 589000 470824 589600 6 gfpga_pad_GPIO_PAD_in[39]
port 36 nsew signal input
rlabel metal3 s 561186 352728 561786 352848 6 gfpga_pad_GPIO_PAD_in[3]
port 37 nsew signal input
rlabel metal3 s 561186 370408 561786 370528 6 gfpga_pad_GPIO_PAD_in[40]
port 38 nsew signal input
rlabel metal2 s 121720 589000 121776 589600 6 gfpga_pad_GPIO_PAD_in[41]
port 39 nsew signal input
rlabel metal2 s 454024 589000 454080 589600 6 gfpga_pad_GPIO_PAD_in[42]
port 40 nsew signal input
rlabel metal2 s 348408 0 348464 600 6 gfpga_pad_GPIO_PAD_in[43]
port 41 nsew signal input
rlabel metal2 s 282076 0 282132 600 6 gfpga_pad_GPIO_PAD_in[44]
port 42 nsew signal input
rlabel metal3 s 561186 405768 561786 405888 6 gfpga_pad_GPIO_PAD_in[45]
port 43 nsew signal input
rlabel metal2 s 548048 0 548104 600 6 gfpga_pad_GPIO_PAD_in[46]
port 44 nsew signal input
rlabel metal2 s 481072 0 481128 600 6 gfpga_pad_GPIO_PAD_in[47]
port 45 nsew signal input
rlabel metal3 s 561186 265008 561786 265128 6 gfpga_pad_GPIO_PAD_in[48]
port 46 nsew signal input
rlabel metal2 s 486868 589000 486924 589600 6 gfpga_pad_GPIO_PAD_in[49]
port 47 nsew signal input
rlabel metal2 s 298820 0 298876 600 6 gfpga_pad_GPIO_PAD_in[4]
port 48 nsew signal input
rlabel metal3 s 561186 177288 561786 177408 6 gfpga_pad_GPIO_PAD_in[50]
port 49 nsew signal input
rlabel metal2 s 132668 0 132724 600 6 gfpga_pad_GPIO_PAD_in[51]
port 50 nsew signal input
rlabel metal2 s 16104 0 16160 600 6 gfpga_pad_GPIO_PAD_in[52]
port 51 nsew signal input
rlabel metal3 s 561186 160288 561786 160408 6 gfpga_pad_GPIO_PAD_in[53]
port 52 nsew signal input
rlabel metal2 s 188052 589000 188108 589600 6 gfpga_pad_GPIO_PAD_in[54]
port 53 nsew signal input
rlabel metal3 s 186 297648 786 297768 6 gfpga_pad_GPIO_PAD_in[55]
port 54 nsew signal input
rlabel metal3 s 186 385368 786 385488 6 gfpga_pad_GPIO_PAD_in[56]
port 55 nsew signal input
rlabel metal3 s 561186 72568 561786 72688 6 gfpga_pad_GPIO_PAD_in[57]
port 56 nsew signal input
rlabel metal2 s 414740 0 414796 600 6 gfpga_pad_GPIO_PAD_in[58]
port 57 nsew signal input
rlabel metal3 s 561186 440448 561786 440568 6 gfpga_pad_GPIO_PAD_in[59]
port 58 nsew signal input
rlabel metal3 s 186 279968 786 280088 6 gfpga_pad_GPIO_PAD_in[5]
port 59 nsew signal input
rlabel metal2 s 215744 0 215800 600 6 gfpga_pad_GPIO_PAD_in[60]
port 60 nsew signal input
rlabel metal2 s 82436 0 82492 600 6 gfpga_pad_GPIO_PAD_in[61]
port 61 nsew signal input
rlabel metal2 s 537100 589000 537156 589600 6 gfpga_pad_GPIO_PAD_in[62]
port 62 nsew signal input
rlabel metal3 s 186 262288 786 262408 6 gfpga_pad_GPIO_PAD_in[63]
port 63 nsew signal input
rlabel metal3 s 186 69848 786 69968 6 gfpga_pad_GPIO_PAD_in[6]
port 64 nsew signal input
rlabel metal3 s 561186 318048 561786 318168 6 gfpga_pad_GPIO_PAD_in[7]
port 65 nsew signal input
rlabel metal2 s 138464 589000 138520 589600 6 gfpga_pad_GPIO_PAD_in[8]
port 66 nsew signal input
rlabel metal3 s 561186 581208 561786 581328 6 gfpga_pad_GPIO_PAD_in[9]
port 67 nsew signal input
rlabel metal3 s 186 403048 786 403168 6 gfpga_pad_GPIO_PAD_out[0]
port 68 nsew signal output
rlabel metal3 s 186 350008 786 350128 6 gfpga_pad_GPIO_PAD_out[10]
port 69 nsew signal output
rlabel metal2 s 38644 589000 38700 589600 6 gfpga_pad_GPIO_PAD_out[11]
port 70 nsew signal output
rlabel metal2 s 171308 589000 171364 589600 6 gfpga_pad_GPIO_PAD_out[12]
port 71 nsew signal output
rlabel metal2 s 221540 589000 221596 589600 6 gfpga_pad_GPIO_PAD_out[13]
port 72 nsew signal output
rlabel metal3 s 186 437728 786 437848 6 gfpga_pad_GPIO_PAD_out[14]
port 73 nsew signal output
rlabel metal3 s 186 86848 786 86968 6 gfpga_pad_GPIO_PAD_out[15]
port 74 nsew signal output
rlabel metal3 s 561186 194968 561786 195088 6 gfpga_pad_GPIO_PAD_out[16]
port 75 nsew signal output
rlabel metal3 s 561186 545848 561786 545968 6 gfpga_pad_GPIO_PAD_out[17]
port 76 nsew signal output
rlabel metal2 s 49592 0 49648 600 6 gfpga_pad_GPIO_PAD_out[18]
port 77 nsew signal output
rlabel metal3 s 561186 37208 561786 37328 6 gfpga_pad_GPIO_PAD_out[19]
port 78 nsew signal output
rlabel metal3 s 561186 212648 561786 212768 6 gfpga_pad_GPIO_PAD_out[1]
port 79 nsew signal output
rlabel metal2 s 387692 589000 387748 589600 6 gfpga_pad_GPIO_PAD_out[20]
port 80 nsew signal output
rlabel metal3 s 561186 124928 561786 125048 6 gfpga_pad_GPIO_PAD_out[21]
port 81 nsew signal output
rlabel metal3 s 186 578488 786 578608 6 gfpga_pad_GPIO_PAD_out[22]
port 82 nsew signal output
rlabel metal3 s 186 315328 786 315448 6 gfpga_pad_GPIO_PAD_out[23]
port 83 nsew signal output
rlabel metal3 s 561186 300368 561786 300488 6 gfpga_pad_GPIO_PAD_out[24]
port 84 nsew signal output
rlabel metal3 s 561186 563528 561786 563648 6 gfpga_pad_GPIO_PAD_out[25]
port 85 nsew signal output
rlabel metal3 s 186 227608 786 227728 6 gfpga_pad_GPIO_PAD_out[26]
port 86 nsew signal output
rlabel metal3 s 561186 89568 561786 89688 6 gfpga_pad_GPIO_PAD_out[27]
port 87 nsew signal output
rlabel metal2 s 331664 0 331720 600 6 gfpga_pad_GPIO_PAD_out[28]
port 88 nsew signal output
rlabel metal2 s 531304 0 531360 600 6 gfpga_pad_GPIO_PAD_out[29]
port 89 nsew signal output
rlabel metal2 s 238284 589000 238340 589600 6 gfpga_pad_GPIO_PAD_out[2]
port 90 nsew signal output
rlabel metal2 s 431484 0 431540 600 6 gfpga_pad_GPIO_PAD_out[30]
port 91 nsew signal output
rlabel metal2 s 66336 0 66392 600 6 gfpga_pad_GPIO_PAD_out[31]
port 92 nsew signal output
rlabel metal3 s 186 209928 786 210048 6 gfpga_pad_GPIO_PAD_out[32]
port 93 nsew signal output
rlabel metal3 s 561186 54888 561786 55008 6 gfpga_pad_GPIO_PAD_out[33]
port 94 nsew signal output
rlabel metal3 s 561186 422768 561786 422888 6 gfpga_pad_GPIO_PAD_out[34]
port 95 nsew signal output
rlabel metal3 s 186 16808 786 16928 6 gfpga_pad_GPIO_PAD_out[35]
port 96 nsew signal output
rlabel metal2 s 464972 0 465028 600 6 gfpga_pad_GPIO_PAD_out[36]
port 97 nsew signal output
rlabel metal3 s 186 367688 786 367808 6 gfpga_pad_GPIO_PAD_out[37]
port 98 nsew signal output
rlabel metal3 s 561186 142608 561786 142728 6 gfpga_pad_GPIO_PAD_out[38]
port 99 nsew signal output
rlabel metal3 s 186 490768 786 490888 6 gfpga_pad_GPIO_PAD_out[39]
port 100 nsew signal output
rlabel metal3 s 561186 335728 561786 335848 6 gfpga_pad_GPIO_PAD_out[3]
port 101 nsew signal output
rlabel metal3 s 561186 493488 561786 493608 6 gfpga_pad_GPIO_PAD_out[40]
port 102 nsew signal output
rlabel metal2 s 514560 0 514616 600 6 gfpga_pad_GPIO_PAD_out[41]
port 103 nsew signal output
rlabel metal3 s 561186 528168 561786 528288 6 gfpga_pad_GPIO_PAD_out[42]
port 104 nsew signal output
rlabel metal3 s 186 34488 786 34608 6 gfpga_pad_GPIO_PAD_out[43]
port 105 nsew signal output
rlabel metal3 s 186 525448 786 525568 6 gfpga_pad_GPIO_PAD_out[44]
port 106 nsew signal output
rlabel metal3 s 186 192248 786 192368 6 gfpga_pad_GPIO_PAD_out[45]
port 107 nsew signal output
rlabel metal2 s 4 0 60 600 6 gfpga_pad_GPIO_PAD_out[46]
port 108 nsew signal output
rlabel metal2 s 381896 0 381952 600 6 gfpga_pad_GPIO_PAD_out[47]
port 109 nsew signal output
rlabel metal3 s 186 560808 786 560928 6 gfpga_pad_GPIO_PAD_out[48]
port 110 nsew signal output
rlabel metal2 s 155208 589000 155264 589600 6 gfpga_pad_GPIO_PAD_out[49]
port 111 nsew signal output
rlabel metal2 s 354204 589000 354260 589600 6 gfpga_pad_GPIO_PAD_out[4]
port 112 nsew signal output
rlabel metal3 s 186 455408 786 455528 6 gfpga_pad_GPIO_PAD_out[50]
port 113 nsew signal output
rlabel metal2 s 99180 0 99236 600 6 gfpga_pad_GPIO_PAD_out[51]
port 114 nsew signal output
rlabel metal2 s 32848 0 32904 600 6 gfpga_pad_GPIO_PAD_out[52]
port 115 nsew signal output
rlabel metal2 s 437280 589000 437336 589600 6 gfpga_pad_GPIO_PAD_out[53]
port 116 nsew signal output
rlabel metal2 s 321360 589000 321416 589600 6 gfpga_pad_GPIO_PAD_out[54]
port 117 nsew signal output
rlabel metal2 s 265332 0 265388 600 6 gfpga_pad_GPIO_PAD_out[55]
port 118 nsew signal output
rlabel metal2 s 503612 589000 503668 589600 6 gfpga_pad_GPIO_PAD_out[56]
port 119 nsew signal output
rlabel metal3 s 561186 107248 561786 107368 6 gfpga_pad_GPIO_PAD_out[57]
port 120 nsew signal output
rlabel metal3 s 186 543128 786 543248 6 gfpga_pad_GPIO_PAD_out[58]
port 121 nsew signal output
rlabel metal3 s 186 174568 786 174688 6 gfpga_pad_GPIO_PAD_out[59]
port 122 nsew signal output
rlabel metal2 s 115924 0 115980 600 6 gfpga_pad_GPIO_PAD_out[5]
port 123 nsew signal output
rlabel metal2 s 199000 0 199056 600 6 gfpga_pad_GPIO_PAD_out[60]
port 124 nsew signal output
rlabel metal3 s 186 52168 786 52288 6 gfpga_pad_GPIO_PAD_out[61]
port 125 nsew signal output
rlabel metal3 s 561186 388088 561786 388208 6 gfpga_pad_GPIO_PAD_out[62]
port 126 nsew signal output
rlabel metal2 s 315564 0 315620 600 6 gfpga_pad_GPIO_PAD_out[63]
port 127 nsew signal output
rlabel metal2 s 420536 589000 420592 589600 6 gfpga_pad_GPIO_PAD_out[6]
port 128 nsew signal output
rlabel metal2 s 403792 589000 403848 589600 6 gfpga_pad_GPIO_PAD_out[7]
port 129 nsew signal output
rlabel metal2 s 5156 589000 5212 589600 6 gfpga_pad_GPIO_PAD_out[8]
port 130 nsew signal output
rlabel metal2 s 104976 589000 105032 589600 6 gfpga_pad_GPIO_PAD_out[9]
port 131 nsew signal output
rlabel metal2 s 398640 0 398696 600 6 pReset
port 132 nsew signal input
rlabel metal3 s 186 157568 786 157688 6 prog_clk
port 133 nsew signal input
rlabel metal3 s 186 507768 786 507888 6 reset
port 134 nsew signal input
rlabel metal3 s 561186 282688 561786 282808 6 set
port 135 nsew signal input
rlabel metal4 s 8330 1928 8650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 22330 1928 22650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 36330 1928 36650 60495 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 36330 98409 36650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 50330 1928 50650 60495 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 50330 98409 50650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 64330 1928 64650 110903 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 64330 149225 64650 212903 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 64330 251225 64650 314903 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 64330 353225 64650 430231 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 64330 449649 64650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 78330 1928 78650 110903 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 78330 149225 78650 212903 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 78330 251225 78650 314903 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 78330 353225 78650 430231 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 78330 449649 78650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 92330 1928 92650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 106330 1928 106650 159868 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 106330 203252 106650 261868 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 106330 305252 106650 363868 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 106330 407252 106650 465868 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 106330 509252 106650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 120330 1928 120650 160767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 120330 197865 120650 262767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 120330 299865 120650 364767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 120330 401865 120650 416087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 120330 454953 120650 466767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 120330 503865 120650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 134330 1928 134650 160767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 134330 197865 134650 212903 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 134330 224977 134650 262767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 134330 299865 134650 364767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 134330 401865 134650 416087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 134330 454953 134650 466767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 134330 503865 134650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 148330 1928 148650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 162330 1928 162650 67159 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 162330 96505 162650 112087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 162330 146465 162650 214087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 162330 248465 162650 316087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 162330 350465 162650 418359 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 162330 448929 162650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 176330 1928 176650 67159 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 176330 96505 176650 112087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 176330 146465 176650 214087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 176330 248465 176650 316087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 176330 350465 176650 418359 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 176330 448929 176650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 190330 1928 190650 112087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 190330 146465 190650 214087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 190330 248465 190650 316087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 190330 350465 190650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 204330 1928 204650 160767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 204330 197865 204650 262767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 204330 299865 204650 364767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 204330 401865 204650 466767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 204330 503865 204650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 218330 1928 218650 160767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 218330 197865 218650 262767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 218330 299865 218650 364767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 218330 401865 218650 466767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 218330 503865 218650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 232330 1928 232650 56223 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 232330 75505 232650 110903 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 232330 122977 232650 160767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 232330 197865 232650 212903 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 232330 224977 232650 262767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 232330 299865 232650 314903 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 232330 326977 232650 364767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 232330 401865 232650 416087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 232330 454953 232650 466767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 232330 503865 232650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 246330 1928 246650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 260330 1928 260650 67159 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 260330 96505 260650 112087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 260330 146465 260650 214087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 260330 248465 260650 316087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 260330 350465 260650 418359 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 260330 448929 260650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 274330 1928 274650 67159 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 274330 96505 274650 112087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 274330 146465 274650 214087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 274330 248465 274650 316087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 274330 350465 274650 418359 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 274330 448929 274650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 288330 1928 288650 112087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 288330 146465 288650 214087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 288330 248465 288650 316087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 288330 350465 288650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 302330 1928 302650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 316330 1928 316650 160767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 316330 197865 316650 262767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 316330 299865 316650 364767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 316330 401865 316650 466767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 316330 503865 316650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 330330 1928 330650 56223 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 330330 75505 330650 160767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 330330 197865 330650 262767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 330330 299865 330650 364767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 330330 401865 330650 416087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 330330 454953 330650 466767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 330330 503865 330650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 344330 1928 344650 160767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 344330 197865 344650 262767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 344330 299865 344650 364767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 344330 401865 344650 466767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 344330 503865 344650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 358330 1928 358650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 372330 1928 372650 67159 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 372330 96505 372650 112087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 372330 146465 372650 214087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 372330 248465 372650 316087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 372330 350465 372650 418359 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 372330 448929 372650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 386330 1928 386650 67159 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 386330 96505 386650 112087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 386330 146465 386650 165255 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 386330 185489 386650 214087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 386330 248465 386650 267255 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 386330 287489 386650 316087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 386330 350465 386650 369255 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 386330 389489 386650 471255 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 386330 491489 386650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 400330 1928 400650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 414330 1928 414650 160767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 414330 197865 414650 262767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 414330 299865 414650 364767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 414330 401865 414650 466767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 414330 503865 414650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 428330 1928 428650 56223 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 428330 75505 428650 160767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 428330 197865 428650 262767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 428330 299865 428650 364767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 428330 401865 428650 416087 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 428330 454953 428650 466767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 428330 503865 428650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 442330 1928 442650 160767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 442330 197865 442650 262767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 442330 299865 442650 364767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 442330 401865 442650 466767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 442330 503865 442650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 456330 1928 456650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 470330 1928 470650 61719 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 470330 98545 470650 108359 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 470330 145865 470650 154855 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 470330 173729 470650 204359 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 470330 241865 470650 256855 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 470330 275729 470650 306359 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 470330 343865 470650 358855 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 470330 377729 470650 460855 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 470330 479729 470650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 484330 1928 484650 61719 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 484330 98545 484650 108359 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 484330 145865 484650 204359 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 484330 241865 484650 306359 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 484330 343865 484650 408767 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 484330 435257 484650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 498330 1928 498650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 512330 1928 512650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 526330 1928 526650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 540330 1928 540650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 554330 1928 554650 587368 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 9216 560866 9536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 24216 560866 24536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 39216 560866 39536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 54216 560866 54536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 69216 560866 69536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 84216 560866 84536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 99216 560866 99536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 114216 560866 114536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 129216 560866 129536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 144216 560866 144536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 159216 560866 159536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 174216 560866 174536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 189216 560866 189536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 204216 560866 204536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 219216 560866 219536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 234216 560866 234536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 249216 560866 249536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 264216 560866 264536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 279216 560866 279536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 294216 560866 294536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 309216 560866 309536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 324216 560866 324536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 339216 560866 339536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 354216 560866 354536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 369216 560866 369536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 384216 560866 384536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 399216 560866 399536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 414216 560866 414536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 429216 560866 429536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 444216 560866 444536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 459216 560866 459536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 474216 560866 474536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 489216 560866 489536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 504216 560866 504536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 519216 560866 519536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 534216 560866 534536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 549216 560866 549536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 564216 560866 564536 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 1042 579216 560866 579536 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 2494 104744 2814 150536 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 102406 209192 102726 254440 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 251262 313640 251582 356168 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 353014 414824 353334 458440 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 403430 156968 403750 160872 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 506470 254888 506790 297416 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 557990 357160 558310 402408 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 2494 207016 2814 252808 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 100934 106920 101254 152712 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 199558 156968 199878 202760 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 251262 414824 251582 458440 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 353014 313096 353334 356712 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 404902 56872 405222 98856 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 506470 357160 506790 399688 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 557990 254888 558310 300680 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 2494 308744 2814 354536 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 100934 413192 101254 458440 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 251262 211368 251582 253896 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 353934 56872 354254 98856 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 403430 160932 403750 202760 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 506470 458888 506790 501416 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 2494 411016 2814 456808 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 100934 310920 101254 356712 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 251262 109096 251582 152712 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 354486 156968 354806 202760 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 403430 258696 403750 262600 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 557990 458888 558310 504680 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 199558 258696 199878 304488 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 251998 56872 252318 98856 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 353014 109096 353334 154888 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 404902 210824 405222 255528 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 252550 156968 252870 202760 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 353014 210824 353334 254440 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 404902 109096 405222 152712 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 199558 360968 199878 406760 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 252550 258696 252870 304488 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 354486 462696 354806 508488 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 404902 313096 405222 356712 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 506470 153160 506790 195688 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 252550 360968 252870 406760 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 354486 258696 354806 304488 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 403430 462696 403750 466600 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 557990 153160 558310 198408 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 199558 462696 199878 508488 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 354486 360968 354806 406760 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 403430 262660 403750 304488 6 vccd1
port 136 nsew power bidirectional
rlabel metal5 s 456330 149580 485310 149900 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 252550 462696 252870 508488 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 403430 360968 403750 364872 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 403430 364932 403750 406760 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 404902 414824 405222 458440 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 403430 466660 403750 508488 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 8990 1928 9310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 22990 1928 23310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 36990 1928 37310 60495 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 36990 98409 37310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 50990 1928 51310 60495 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 50990 98409 51310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 64990 1928 65310 110903 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 64990 149225 65310 212903 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 64990 251225 65310 314903 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 64990 353225 65310 430231 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 64990 449649 65310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 78990 1928 79310 110903 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 78990 149225 79310 212903 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 78990 251225 79310 314903 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 78990 353225 79310 430231 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 78990 449649 79310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 92990 1928 93310 109868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 92990 149444 93310 211868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 92990 251444 93310 313868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 92990 353444 93310 415868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 92990 455444 93310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 106990 1928 107310 160767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 106990 197865 107310 262767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 106990 299865 107310 364767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 106990 401865 107310 466767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 106990 503865 107310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 120990 1928 121310 160767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 120990 197865 121310 262767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 120990 299865 121310 364767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 120990 401865 121310 416087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 120990 454953 121310 466767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 120990 503865 121310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 134990 1928 135310 160767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 134990 197865 135310 262767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 134990 299865 135310 364767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 134990 401865 135310 466767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 134990 503865 135310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 148990 1928 149310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 162990 1928 163310 67159 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 162990 96505 163310 112087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 162990 146465 163310 214087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 162990 248465 163310 316087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 162990 350465 163310 418359 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 162990 448929 163310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 176990 1928 177310 67159 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 176990 96505 177310 112087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 176990 146465 177310 214087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 176990 248465 177310 316087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 176990 350465 177310 418359 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 176990 448929 177310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 190990 1928 191310 59868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 190990 99444 191310 111868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 190990 151444 191310 159868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 190990 199444 191310 213868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 190990 253444 191310 261868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 190990 301444 191310 315868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 190990 355444 191310 363868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 190990 403444 191310 417868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 190990 457444 191310 465868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 190990 505444 191310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 204990 1928 205310 160767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 204990 197865 205310 262767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 204990 299865 205310 364767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 204990 401865 205310 466767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 204990 503865 205310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 218990 1928 219310 160767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 218990 197865 219310 262767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 218990 299865 219310 364767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 218990 401865 219310 466767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 218990 503865 219310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 232990 1928 233310 110903 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 232990 122977 233310 160767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 232990 197865 233310 212903 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 232990 224977 233310 262767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 232990 299865 233310 314903 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 232990 326977 233310 364767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 232990 401865 233310 416087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 232990 454953 233310 466767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 232990 503865 233310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 246990 1928 247310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 260990 1928 261310 67159 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 260990 96505 261310 112087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 260990 146465 261310 214087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 260990 248465 261310 316087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 260990 350465 261310 418359 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 260990 448929 261310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 274990 1928 275310 67159 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 274990 96505 275310 112087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 274990 146465 275310 214087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 274990 248465 275310 316087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 274990 350465 275310 418359 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 274990 448929 275310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 288990 1928 289310 112087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 288990 146465 289310 214087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 288990 248465 289310 316087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 288990 350465 289310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 302990 1928 303310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 316990 1928 317310 5868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 316990 45444 317310 160767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 316990 197865 317310 262767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 316990 299865 317310 364767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 316990 401865 317310 466767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 316990 503865 317310 521868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 316990 561444 317310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 330990 1928 331310 56223 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 330990 75505 331310 160767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 330990 197865 331310 262767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 330990 299865 331310 364767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 330990 401865 331310 416087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 330990 454953 331310 466767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 330990 503865 331310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 344990 1928 345310 160767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 344990 197865 345310 262767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 344990 299865 345310 364767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 344990 401865 345310 466767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 344990 503865 345310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 358990 1928 359310 418359 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 358990 448929 359310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 372990 1928 373310 67159 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 372990 96505 373310 112087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 372990 146465 373310 214087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 372990 248465 373310 316087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 372990 350465 373310 418359 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 372990 448929 373310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 386990 1928 387310 67159 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 386990 96505 387310 112087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 386990 146465 387310 165255 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 386990 185489 387310 214087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 386990 248465 387310 267255 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 386990 287489 387310 316087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 386990 350465 387310 369255 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 386990 389489 387310 471255 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 386990 491489 387310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 400990 1928 401310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 414990 1928 415310 55868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 414990 95444 415310 109868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 414990 149444 415310 160767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 414990 197865 415310 212468 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 414990 252044 415310 262767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 414990 299865 415310 313868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 414990 353444 415310 364767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 414990 401865 415310 415868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 414990 455444 415310 466767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 414990 503865 415310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 428990 1928 429310 56223 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 428990 75505 429310 160767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 428990 197865 429310 262767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 428990 299865 429310 364767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 428990 401865 429310 416087 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 428990 454953 429310 466767 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 428990 503865 429310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 442990 1928 443310 159868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 442990 203252 443310 261868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 442990 305252 443310 363868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 442990 407252 443310 465868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 442990 509252 443310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 456990 1928 457310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 470990 1928 471310 61719 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 470990 98545 471310 108359 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 470990 145865 471310 154855 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 470990 173729 471310 204359 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 470990 241865 471310 256855 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 470990 275729 471310 306359 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 470990 343865 471310 358855 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 470990 377729 471310 460855 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 470990 479729 471310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 484990 1928 485310 61719 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 484990 98545 485310 108359 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 484990 145865 485310 204359 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 484990 241865 485310 306359 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 484990 343865 485310 407868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 484990 437652 485310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 498990 1928 499310 407868 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 498990 437652 499310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 512990 1928 513310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 526990 1928 527310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 540990 1928 541310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 554990 1928 555310 587368 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 9876 560866 10196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 24876 560866 25196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 39876 560866 40196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 54876 560866 55196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 69876 560866 70196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 84876 560866 85196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 99876 560866 100196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 114876 560866 115196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 129876 560866 130196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 144876 560866 145196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 159876 560866 160196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 174876 560866 175196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 189876 560866 190196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 204876 560866 205196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 219876 560866 220196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 234876 560866 235196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 249876 560866 250196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 264876 560866 265196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 279876 560866 280196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 294876 560866 295196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 309876 560866 310196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 324876 560866 325196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 339876 560866 340196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 354876 560866 355196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 369876 560866 370196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 384876 560866 385196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 399876 560866 400196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 414876 560866 415196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 429876 560866 430196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 444876 560866 445196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 459876 560866 460196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 474876 560866 475196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 489876 560866 490196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 504876 560866 505196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 519876 560866 520196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 534876 560866 535196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 549876 560866 550196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 564876 560866 565196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 1042 579876 560866 580196 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 3230 104744 3550 150536 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 103142 209192 103462 254440 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 201398 57416 201718 98856 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 353750 414824 354070 458440 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 404166 156968 404486 160872 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 507206 254888 507526 297416 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 558726 357160 559046 402408 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 3230 207016 3550 252808 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 101670 106920 101990 152712 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 200294 156968 200614 202760 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 353750 313096 354070 356712 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 405638 56872 405958 98856 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 507206 357160 507526 399688 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 558726 254888 559046 300680 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 3230 308744 3550 354536 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 101670 413192 101990 458440 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 201398 109640 201718 152168 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 354670 56872 354990 98856 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 404166 160932 404486 202760 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 507206 458888 507526 501416 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 3230 411016 3550 456808 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 101670 310920 101990 356712 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 201398 210824 201718 254440 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 355222 156968 355542 202760 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 404166 258696 404486 262600 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 558726 458888 559046 504680 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 200294 258696 200614 304488 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 252734 56872 253054 98856 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 353750 109096 354070 154888 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 405638 210824 405958 255528 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 201398 313096 201718 356712 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 253286 156968 253606 202760 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 353750 210824 354070 254440 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 405638 109096 405958 152712 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 200294 360968 200614 406760 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 253286 258696 253606 304488 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 355222 462696 355542 508488 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 405638 313096 405958 356712 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 507206 153160 507526 195688 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 201398 415368 201718 457896 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 253286 360968 253606 406760 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 355222 258696 355542 304488 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 404166 462696 404486 466600 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 558726 153160 559046 198408 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 200294 462696 200614 508488 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 355222 360968 355542 406760 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 404166 262660 404486 304488 6 vssd1
port 137 nsew ground bidirectional
rlabel metal5 s 456330 150260 485310 150580 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 253286 462696 253606 508488 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 404166 360968 404486 364872 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 404166 364932 404486 406760 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 405638 414824 405958 458440 6 vssd1
port 137 nsew ground bidirectional
rlabel metal4 s 404166 466660 404486 508488 6 vssd1
port 137 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 561786 589600
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 95819482
string GDS_FILE /home/baungarten/Proyectos_caravel/FPGA_3/openlane/fpga_top_2/runs/22_12_30_22_35/results/signoff/fpga_top.magic.gds
string GDS_START 37389160
<< end >>

