magic
tech sky130A
magscale 1 2
timestamp 1672416771
<< viali >>
rect 17693 37417 17727 37451
rect 12449 37281 12483 37315
rect 14473 37281 14507 37315
rect 14933 37281 14967 37315
rect 16313 37281 16347 37315
rect 17141 37281 17175 37315
rect 18153 37281 18187 37315
rect 21465 37281 21499 37315
rect 22017 37281 22051 37315
rect 35081 37281 35115 37315
rect 35541 37281 35575 37315
rect 36921 37281 36955 37315
rect 38301 37281 38335 37315
rect 1869 37213 1903 37247
rect 2973 37213 3007 37247
rect 4905 37213 4939 37247
rect 6837 37213 6871 37247
rect 7389 37213 7423 37247
rect 7941 37213 7975 37247
rect 10057 37213 10091 37247
rect 11989 37213 12023 37247
rect 13277 37213 13311 37247
rect 15209 37213 15243 37247
rect 16957 37213 16991 37247
rect 18337 37213 18371 37247
rect 20085 37213 20119 37247
rect 22293 37213 22327 37247
rect 23305 37213 23339 37247
rect 25237 37213 25271 37247
rect 27169 37213 27203 37247
rect 28457 37213 28491 37247
rect 30389 37213 30423 37247
rect 32321 37213 32355 37247
rect 33609 37213 33643 37247
rect 35817 37213 35851 37247
rect 38025 37213 38059 37247
rect 1685 37077 1719 37111
rect 2789 37077 2823 37111
rect 4721 37077 4755 37111
rect 5457 37077 5491 37111
rect 6653 37077 6687 37111
rect 8033 37077 8067 37111
rect 9873 37077 9907 37111
rect 11805 37077 11839 37111
rect 13093 37077 13127 37111
rect 20269 37077 20303 37111
rect 23489 37077 23523 37111
rect 25421 37077 25455 37111
rect 27353 37077 27387 37111
rect 28641 37077 28675 37111
rect 30573 37077 30607 37111
rect 32505 37077 32539 37111
rect 33793 37077 33827 37111
rect 22201 36873 22235 36907
rect 27997 36873 28031 36907
rect 37565 36873 37599 36907
rect 2421 36805 2455 36839
rect 1685 36737 1719 36771
rect 3065 36737 3099 36771
rect 10609 36737 10643 36771
rect 22017 36737 22051 36771
rect 27813 36737 27847 36771
rect 36737 36737 36771 36771
rect 37749 36737 37783 36771
rect 38209 36737 38243 36771
rect 1869 36601 1903 36635
rect 2513 36533 2547 36567
rect 10425 36533 10459 36567
rect 22753 36533 22787 36567
rect 36921 36533 36955 36567
rect 2421 36329 2455 36363
rect 37473 36329 37507 36363
rect 38209 36329 38243 36363
rect 1869 36125 1903 36159
rect 37289 36125 37323 36159
rect 38025 36125 38059 36159
rect 1685 35989 1719 36023
rect 36737 35989 36771 36023
rect 2145 35785 2179 35819
rect 2237 35649 2271 35683
rect 38025 35581 38059 35615
rect 38301 35581 38335 35615
rect 2789 35445 2823 35479
rect 20269 35241 20303 35275
rect 29929 35241 29963 35275
rect 38301 35241 38335 35275
rect 20085 35037 20119 35071
rect 20729 35037 20763 35071
rect 29745 35037 29779 35071
rect 30389 35037 30423 35071
rect 1869 34561 1903 34595
rect 2329 34493 2363 34527
rect 1685 34357 1719 34391
rect 7021 34153 7055 34187
rect 7113 33949 7147 33983
rect 7573 33949 7607 33983
rect 37473 33473 37507 33507
rect 38025 33473 38059 33507
rect 38209 33337 38243 33371
rect 1685 32385 1719 32419
rect 38025 32385 38059 32419
rect 38301 32317 38335 32351
rect 1777 32181 1811 32215
rect 1593 31977 1627 32011
rect 38301 31977 38335 32011
rect 27445 30889 27479 30923
rect 30849 30889 30883 30923
rect 27261 30685 27295 30719
rect 30757 30685 30791 30719
rect 31401 30685 31435 30719
rect 1685 30617 1719 30651
rect 1777 30549 1811 30583
rect 27997 30549 28031 30583
rect 1685 30345 1719 30379
rect 15393 30209 15427 30243
rect 38025 30209 38059 30243
rect 14749 30005 14783 30039
rect 15485 30005 15519 30039
rect 38209 30005 38243 30039
rect 38025 29801 38059 29835
rect 37841 29597 37875 29631
rect 38117 29257 38151 29291
rect 20545 29121 20579 29155
rect 1593 29053 1627 29087
rect 1869 29053 1903 29087
rect 20453 28985 20487 29019
rect 22293 28713 22327 28747
rect 1593 28645 1627 28679
rect 13277 28509 13311 28543
rect 21833 28509 21867 28543
rect 13369 28373 13403 28407
rect 21741 28373 21775 28407
rect 14473 28169 14507 28203
rect 14565 28033 14599 28067
rect 37473 28033 37507 28067
rect 38025 28033 38059 28067
rect 38209 27897 38243 27931
rect 15117 27829 15151 27863
rect 22109 27013 22143 27047
rect 1869 26945 1903 26979
rect 22293 26945 22327 26979
rect 30665 26945 30699 26979
rect 38025 26877 38059 26911
rect 38301 26877 38335 26911
rect 1685 26741 1719 26775
rect 22937 26741 22971 26775
rect 30573 26741 30607 26775
rect 38301 26537 38335 26571
rect 16497 26469 16531 26503
rect 15761 26333 15795 26367
rect 16313 26333 16347 26367
rect 18889 25993 18923 26027
rect 19073 25857 19107 25891
rect 19533 25857 19567 25891
rect 13001 25449 13035 25483
rect 28457 25449 28491 25483
rect 1593 25245 1627 25279
rect 1869 25245 1903 25279
rect 13737 25245 13771 25279
rect 16129 25245 16163 25279
rect 16773 25245 16807 25279
rect 27905 25245 27939 25279
rect 16221 25177 16255 25211
rect 13645 25109 13679 25143
rect 27813 25109 27847 25143
rect 1593 24905 1627 24939
rect 37565 24769 37599 24803
rect 38025 24769 38059 24803
rect 38209 24565 38243 24599
rect 31309 24361 31343 24395
rect 30757 24157 30791 24191
rect 30665 24021 30699 24055
rect 1869 23681 1903 23715
rect 1685 23477 1719 23511
rect 14841 22593 14875 22627
rect 15301 22593 15335 22627
rect 37565 22593 37599 22627
rect 38209 22593 38243 22627
rect 38025 22457 38059 22491
rect 14749 22389 14783 22423
rect 6561 21641 6595 21675
rect 19993 21641 20027 21675
rect 25881 21641 25915 21675
rect 1869 21505 1903 21539
rect 6745 21505 6779 21539
rect 19809 21505 19843 21539
rect 20453 21505 20487 21539
rect 25697 21505 25731 21539
rect 26341 21505 26375 21539
rect 38025 21505 38059 21539
rect 1685 21301 1719 21335
rect 7297 21301 7331 21335
rect 37473 21301 37507 21335
rect 38209 21301 38243 21335
rect 1777 21097 1811 21131
rect 1961 20893 1995 20927
rect 19441 20757 19475 20791
rect 19349 20485 19383 20519
rect 19441 20485 19475 20519
rect 19165 20349 19199 20383
rect 19993 20213 20027 20247
rect 2329 20009 2363 20043
rect 19533 20009 19567 20043
rect 23673 20009 23707 20043
rect 1869 19805 1903 19839
rect 2513 19805 2547 19839
rect 2973 19805 3007 19839
rect 18705 19805 18739 19839
rect 19625 19805 19659 19839
rect 20269 19805 20303 19839
rect 20729 19805 20763 19839
rect 23213 19805 23247 19839
rect 20177 19737 20211 19771
rect 1685 19669 1719 19703
rect 18153 19669 18187 19703
rect 18797 19669 18831 19703
rect 23121 19669 23155 19703
rect 1961 19465 1995 19499
rect 2145 19329 2179 19363
rect 9689 19329 9723 19363
rect 9781 19329 9815 19363
rect 12633 19329 12667 19363
rect 19625 19329 19659 19363
rect 20361 19329 20395 19363
rect 20453 19329 20487 19363
rect 38025 19329 38059 19363
rect 12817 19261 12851 19295
rect 20913 19261 20947 19295
rect 19165 19193 19199 19227
rect 22109 19193 22143 19227
rect 2697 19125 2731 19159
rect 11989 19125 12023 19159
rect 19717 19125 19751 19159
rect 23029 19125 23063 19159
rect 23673 19125 23707 19159
rect 38209 19125 38243 19159
rect 18245 18921 18279 18955
rect 20177 18785 20211 18819
rect 16865 18717 16899 18751
rect 22109 18717 22143 18751
rect 22753 18717 22787 18751
rect 23673 18717 23707 18751
rect 16221 18649 16255 18683
rect 20361 18649 20395 18683
rect 20453 18649 20487 18683
rect 21005 18649 21039 18683
rect 17417 18581 17451 18615
rect 18797 18581 18831 18615
rect 22293 18581 22327 18615
rect 23581 18581 23615 18615
rect 24593 18581 24627 18615
rect 25237 18581 25271 18615
rect 1777 18377 1811 18411
rect 4629 18377 4663 18411
rect 16221 18309 16255 18343
rect 17049 18309 17083 18343
rect 18889 18309 18923 18343
rect 20085 18309 20119 18343
rect 22569 18309 22603 18343
rect 22661 18309 22695 18343
rect 1685 18241 1719 18275
rect 4813 18241 4847 18275
rect 15669 18241 15703 18275
rect 16129 18241 16163 18275
rect 21281 18241 21315 18275
rect 23765 18241 23799 18275
rect 24593 18241 24627 18275
rect 25053 18241 25087 18275
rect 25697 18241 25731 18275
rect 16957 18173 16991 18207
rect 18797 18173 18831 18207
rect 19993 18173 20027 18207
rect 17509 18105 17543 18139
rect 19349 18105 19383 18139
rect 20545 18105 20579 18139
rect 22109 18105 22143 18139
rect 23857 18105 23891 18139
rect 5365 18037 5399 18071
rect 18245 18037 18279 18071
rect 21189 18037 21223 18071
rect 23305 18037 23339 18071
rect 24501 18037 24535 18071
rect 25145 18037 25179 18071
rect 22385 17833 22419 17867
rect 1593 17765 1627 17799
rect 24685 17765 24719 17799
rect 20269 17697 20303 17731
rect 20637 17697 20671 17731
rect 23029 17697 23063 17731
rect 14473 17629 14507 17663
rect 15025 17629 15059 17663
rect 15669 17629 15703 17663
rect 16681 17629 16715 17663
rect 17325 17629 17359 17663
rect 18337 17629 18371 17663
rect 19533 17629 19567 17663
rect 21557 17629 21591 17663
rect 22293 17629 22327 17663
rect 25973 17629 26007 17663
rect 26433 17629 26467 17663
rect 17877 17561 17911 17595
rect 19625 17561 19659 17595
rect 20361 17561 20395 17595
rect 23121 17561 23155 17595
rect 23673 17561 23707 17595
rect 25145 17561 25179 17595
rect 25237 17561 25271 17595
rect 15577 17493 15611 17527
rect 16589 17493 16623 17527
rect 17233 17493 17267 17527
rect 18429 17493 18463 17527
rect 21465 17493 21499 17527
rect 25881 17493 25915 17527
rect 27077 17493 27111 17527
rect 21005 17289 21039 17323
rect 16129 17221 16163 17255
rect 17049 17221 17083 17255
rect 19809 17221 19843 17255
rect 23489 17221 23523 17255
rect 24593 17221 24627 17255
rect 25421 17221 25455 17255
rect 14473 17153 14507 17187
rect 14933 17153 14967 17187
rect 18613 17153 18647 17187
rect 21097 17153 21131 17187
rect 22293 17153 22327 17187
rect 24685 17153 24719 17187
rect 26617 17153 26651 17187
rect 37565 17153 37599 17187
rect 38209 17153 38243 17187
rect 15945 17085 15979 17119
rect 16221 17085 16255 17119
rect 16957 17085 16991 17119
rect 18153 17085 18187 17119
rect 19901 17085 19935 17119
rect 22845 17085 22879 17119
rect 23397 17085 23431 17119
rect 24041 17085 24075 17119
rect 25329 17085 25363 17119
rect 27169 17085 27203 17119
rect 17509 17017 17543 17051
rect 19349 17017 19383 17051
rect 25881 17017 25915 17051
rect 38025 17017 38059 17051
rect 13185 16949 13219 16983
rect 13829 16949 13863 16983
rect 14381 16949 14415 16983
rect 15025 16949 15059 16983
rect 18705 16949 18739 16983
rect 22201 16949 22235 16983
rect 26525 16949 26559 16983
rect 19533 16745 19567 16779
rect 20821 16677 20855 16711
rect 22293 16677 22327 16711
rect 28273 16677 28307 16711
rect 14381 16609 14415 16643
rect 17877 16609 17911 16643
rect 25237 16609 25271 16643
rect 26065 16609 26099 16643
rect 26433 16609 26467 16643
rect 13093 16541 13127 16575
rect 13553 16541 13587 16575
rect 16037 16541 16071 16575
rect 16589 16541 16623 16575
rect 16681 16541 16715 16575
rect 17141 16541 17175 16575
rect 21557 16541 21591 16575
rect 27077 16541 27111 16575
rect 27169 16541 27203 16575
rect 27629 16541 27663 16575
rect 14473 16473 14507 16507
rect 15025 16473 15059 16507
rect 17969 16473 18003 16507
rect 18889 16473 18923 16507
rect 19625 16473 19659 16507
rect 20269 16473 20303 16507
rect 20361 16473 20395 16507
rect 22753 16473 22787 16507
rect 22845 16473 22879 16507
rect 24593 16473 24627 16507
rect 25145 16473 25179 16507
rect 26341 16473 26375 16507
rect 11437 16405 11471 16439
rect 12449 16405 12483 16439
rect 13001 16405 13035 16439
rect 13645 16405 13679 16439
rect 15945 16405 15979 16439
rect 17233 16405 17267 16439
rect 21465 16405 21499 16439
rect 23397 16405 23431 16439
rect 27721 16405 27755 16439
rect 28825 16405 28859 16439
rect 18337 16201 18371 16235
rect 26433 16201 26467 16235
rect 28641 16201 28675 16235
rect 13001 16133 13035 16167
rect 14197 16133 14231 16167
rect 14749 16133 14783 16167
rect 15761 16133 15795 16167
rect 17049 16133 17083 16167
rect 19625 16133 19659 16167
rect 20913 16133 20947 16167
rect 23765 16133 23799 16167
rect 24501 16133 24535 16167
rect 25697 16133 25731 16167
rect 27905 16133 27939 16167
rect 29101 16133 29135 16167
rect 1869 16065 1903 16099
rect 11161 16065 11195 16099
rect 12173 16065 12207 16099
rect 18429 16065 18463 16099
rect 19073 16065 19107 16099
rect 22017 16065 22051 16099
rect 22201 16065 22235 16099
rect 24685 16065 24719 16099
rect 26341 16065 26375 16099
rect 27169 16065 27203 16099
rect 27997 16065 28031 16099
rect 28457 16065 28491 16099
rect 37565 16065 37599 16099
rect 38209 16065 38243 16099
rect 12909 15997 12943 16031
rect 14105 15997 14139 16031
rect 15669 15997 15703 16031
rect 16957 15997 16991 16031
rect 19717 15997 19751 16031
rect 21005 15997 21039 16031
rect 23213 15997 23247 16031
rect 23857 15997 23891 16031
rect 25789 15997 25823 16031
rect 10149 15929 10183 15963
rect 13461 15929 13495 15963
rect 16221 15929 16255 15963
rect 17509 15929 17543 15963
rect 20453 15929 20487 15963
rect 25237 15929 25271 15963
rect 38025 15929 38059 15963
rect 1685 15861 1719 15895
rect 12265 15861 12299 15895
rect 27261 15861 27295 15895
rect 8125 15657 8159 15691
rect 9689 15657 9723 15691
rect 12541 15657 12575 15691
rect 18797 15657 18831 15691
rect 30941 15657 30975 15691
rect 15853 15589 15887 15623
rect 17049 15589 17083 15623
rect 24685 15589 24719 15623
rect 11897 15521 11931 15555
rect 13277 15521 13311 15555
rect 14381 15521 14415 15555
rect 19717 15521 19751 15555
rect 23121 15521 23155 15555
rect 23397 15521 23431 15555
rect 25237 15521 25271 15555
rect 8217 15453 8251 15487
rect 10241 15453 10275 15487
rect 11161 15453 11195 15487
rect 11805 15453 11839 15487
rect 12449 15453 12483 15487
rect 13093 15453 13127 15487
rect 18705 15453 18739 15487
rect 20361 15453 20395 15487
rect 22385 15453 22419 15487
rect 25789 15453 25823 15487
rect 27169 15453 27203 15487
rect 27629 15453 27663 15487
rect 28457 15453 28491 15487
rect 29745 15453 29779 15487
rect 30849 15453 30883 15487
rect 10333 15385 10367 15419
rect 14473 15385 14507 15419
rect 15025 15385 15059 15419
rect 16313 15385 16347 15419
rect 16405 15385 16439 15419
rect 17509 15385 17543 15419
rect 17601 15385 17635 15419
rect 20913 15385 20947 15419
rect 21005 15385 21039 15419
rect 21557 15385 21591 15419
rect 23213 15385 23247 15419
rect 25145 15385 25179 15419
rect 26341 15385 26375 15419
rect 26433 15385 26467 15419
rect 11253 15317 11287 15351
rect 13737 15317 13771 15351
rect 18153 15317 18187 15351
rect 20269 15317 20303 15351
rect 22477 15317 22511 15351
rect 27077 15317 27111 15351
rect 27721 15317 27755 15351
rect 28365 15317 28399 15351
rect 29009 15317 29043 15351
rect 11069 15113 11103 15147
rect 20361 15113 20395 15147
rect 21373 15113 21407 15147
rect 28549 15113 28583 15147
rect 9873 15045 9907 15079
rect 13001 15045 13035 15079
rect 13553 15045 13587 15079
rect 14197 15045 14231 15079
rect 15393 15045 15427 15079
rect 17049 15045 17083 15079
rect 18613 15045 18647 15079
rect 19165 15045 19199 15079
rect 22937 15045 22971 15079
rect 23581 15045 23615 15079
rect 24685 15045 24719 15079
rect 24777 15045 24811 15079
rect 25881 15045 25915 15079
rect 27905 15045 27939 15079
rect 9321 14977 9355 15011
rect 10333 14977 10367 15011
rect 10977 14977 11011 15011
rect 12173 14977 12207 15011
rect 19809 14977 19843 15011
rect 20453 14977 20487 15011
rect 21281 14977 21315 15011
rect 27353 14977 27387 15011
rect 27813 14977 27847 15011
rect 28641 14977 28675 15011
rect 29653 14977 29687 15011
rect 12909 14909 12943 14943
rect 14105 14909 14139 14943
rect 15301 14909 15335 14943
rect 15945 14909 15979 14943
rect 16957 14909 16991 14943
rect 17601 14909 17635 14943
rect 18521 14909 18555 14943
rect 22201 14909 22235 14943
rect 23029 14909 23063 14943
rect 25329 14909 25363 14943
rect 25973 14909 26007 14943
rect 8769 14841 8803 14875
rect 10425 14841 10459 14875
rect 14657 14841 14691 14875
rect 24225 14841 24259 14875
rect 12265 14773 12299 14807
rect 19717 14773 19751 14807
rect 26525 14773 26559 14807
rect 27261 14773 27295 14807
rect 29101 14773 29135 14807
rect 27997 14569 28031 14603
rect 9137 14501 9171 14535
rect 11161 14501 11195 14535
rect 12449 14501 12483 14535
rect 20913 14501 20947 14535
rect 23673 14501 23707 14535
rect 29745 14501 29779 14535
rect 8585 14433 8619 14467
rect 14565 14433 14599 14467
rect 16957 14433 16991 14467
rect 17601 14433 17635 14467
rect 18797 14433 18831 14467
rect 20361 14433 20395 14467
rect 22477 14433 22511 14467
rect 23121 14433 23155 14467
rect 24869 14433 24903 14467
rect 27353 14433 27387 14467
rect 1869 14365 1903 14399
rect 9321 14365 9355 14399
rect 9781 14365 9815 14399
rect 10425 14365 10459 14399
rect 10517 14365 10551 14399
rect 11253 14365 11287 14399
rect 12541 14365 12575 14399
rect 14473 14365 14507 14399
rect 16313 14365 16347 14399
rect 18153 14365 18187 14399
rect 19625 14365 19659 14399
rect 27445 14365 27479 14399
rect 28089 14365 28123 14399
rect 28549 14365 28583 14399
rect 9873 14297 9907 14331
rect 13093 14297 13127 14331
rect 13185 14297 13219 14331
rect 13737 14297 13771 14331
rect 15117 14297 15151 14331
rect 15669 14297 15703 14331
rect 15761 14297 15795 14331
rect 17509 14297 17543 14331
rect 18705 14297 18739 14331
rect 20453 14297 20487 14331
rect 21465 14297 21499 14331
rect 22385 14297 22419 14331
rect 23213 14297 23247 14331
rect 25421 14297 25455 14331
rect 25513 14297 25547 14331
rect 26065 14297 26099 14331
rect 26617 14297 26651 14331
rect 26709 14297 26743 14331
rect 28641 14297 28675 14331
rect 1685 14229 1719 14263
rect 11897 14229 11931 14263
rect 16405 14229 16439 14263
rect 19717 14229 19751 14263
rect 9229 14025 9263 14059
rect 18613 14025 18647 14059
rect 22017 14025 22051 14059
rect 29193 14025 29227 14059
rect 8033 13957 8067 13991
rect 10425 13957 10459 13991
rect 12817 13957 12851 13991
rect 12909 13957 12943 13991
rect 13645 13957 13679 13991
rect 15577 13957 15611 13991
rect 15669 13957 15703 13991
rect 17049 13957 17083 13991
rect 19165 13957 19199 13991
rect 19717 13957 19751 13991
rect 20637 13957 20671 13991
rect 23305 13957 23339 13991
rect 23397 13957 23431 13991
rect 23949 13957 23983 13991
rect 25513 13957 25547 13991
rect 26065 13957 26099 13991
rect 28549 13957 28583 13991
rect 8585 13889 8619 13923
rect 9873 13889 9907 13923
rect 10517 13889 10551 13923
rect 10977 13889 11011 13923
rect 11713 13889 11747 13923
rect 16221 13889 16255 13923
rect 18705 13889 18739 13923
rect 20545 13889 20579 13923
rect 21373 13889 21407 13923
rect 22477 13889 22511 13923
rect 24409 13889 24443 13923
rect 27353 13889 27387 13923
rect 27997 13889 28031 13923
rect 28641 13889 28675 13923
rect 29285 13889 29319 13923
rect 30297 13889 30331 13923
rect 37565 13889 37599 13923
rect 38209 13889 38243 13923
rect 11069 13821 11103 13855
rect 13553 13821 13587 13855
rect 14473 13821 14507 13855
rect 16957 13821 16991 13855
rect 17601 13821 17635 13855
rect 19809 13821 19843 13855
rect 21281 13821 21315 13855
rect 22661 13821 22695 13855
rect 24501 13821 24535 13855
rect 26157 13821 26191 13855
rect 27905 13821 27939 13855
rect 29745 13821 29779 13855
rect 38025 13821 38059 13855
rect 9689 13753 9723 13787
rect 12357 13753 12391 13787
rect 27261 13685 27295 13719
rect 9413 13481 9447 13515
rect 27077 13481 27111 13515
rect 28917 13481 28951 13515
rect 12541 13413 12575 13447
rect 13645 13413 13679 13447
rect 16037 13413 16071 13447
rect 8585 13345 8619 13379
rect 15485 13345 15519 13379
rect 18521 13345 18555 13379
rect 18797 13345 18831 13379
rect 19533 13345 19567 13379
rect 21741 13345 21775 13379
rect 23029 13345 23063 13379
rect 24041 13345 24075 13379
rect 24961 13345 24995 13379
rect 25237 13345 25271 13379
rect 25881 13345 25915 13379
rect 29745 13345 29779 13379
rect 6929 13277 6963 13311
rect 9321 13277 9355 13311
rect 9965 13277 9999 13311
rect 10793 13277 10827 13311
rect 11253 13277 11287 13311
rect 11897 13277 11931 13311
rect 12081 13277 12115 13311
rect 14473 13277 14507 13311
rect 26525 13277 26559 13311
rect 26985 13277 27019 13311
rect 7481 13209 7515 13243
rect 10057 13209 10091 13243
rect 13093 13209 13127 13243
rect 13185 13209 13219 13243
rect 15577 13209 15611 13243
rect 16681 13209 16715 13243
rect 16773 13209 16807 13243
rect 17325 13209 17359 13243
rect 18705 13209 18739 13243
rect 19625 13209 19659 13243
rect 20177 13209 20211 13243
rect 21925 13209 21959 13243
rect 22017 13209 22051 13243
rect 23121 13209 23155 13243
rect 25145 13209 25179 13243
rect 25973 13209 26007 13243
rect 27629 13209 27663 13243
rect 28181 13209 28215 13243
rect 28273 13209 28307 13243
rect 8033 13141 8067 13175
rect 11345 13141 11379 13175
rect 14381 13141 14415 13175
rect 7849 12937 7883 12971
rect 9137 12937 9171 12971
rect 19625 12937 19659 12971
rect 25973 12937 26007 12971
rect 28549 12937 28583 12971
rect 6745 12869 6779 12903
rect 11805 12869 11839 12903
rect 11897 12869 11931 12903
rect 13369 12869 13403 12903
rect 14933 12869 14967 12903
rect 15761 12869 15795 12903
rect 18061 12869 18095 12903
rect 20453 12869 20487 12903
rect 20545 12869 20579 12903
rect 21465 12869 21499 12903
rect 22845 12869 22879 12903
rect 23489 12869 23523 12903
rect 24041 12869 24075 12903
rect 24685 12869 24719 12903
rect 25260 12869 25294 12903
rect 27261 12869 27295 12903
rect 29653 12869 29687 12903
rect 1869 12801 1903 12835
rect 7757 12801 7791 12835
rect 8401 12801 8435 12835
rect 9045 12801 9079 12835
rect 9873 12801 9907 12835
rect 10517 12801 10551 12835
rect 10977 12801 11011 12835
rect 16313 12801 16347 12835
rect 17417 12801 17451 12835
rect 26065 12801 26099 12835
rect 27353 12801 27387 12835
rect 27997 12801 28031 12835
rect 28641 12801 28675 12835
rect 30757 12801 30791 12835
rect 7297 12733 7331 12767
rect 9781 12733 9815 12767
rect 13277 12733 13311 12767
rect 14749 12733 14783 12767
rect 15025 12733 15059 12767
rect 15669 12733 15703 12767
rect 17969 12733 18003 12767
rect 18521 12733 18555 12767
rect 22293 12733 22327 12767
rect 22937 12733 22971 12767
rect 24133 12733 24167 12767
rect 25329 12733 25363 12767
rect 30205 12733 30239 12767
rect 8493 12665 8527 12699
rect 12357 12665 12391 12699
rect 13829 12665 13863 12699
rect 17325 12665 17359 12699
rect 26525 12665 26559 12699
rect 27905 12665 27939 12699
rect 1685 12597 1719 12631
rect 10425 12597 10459 12631
rect 11069 12597 11103 12631
rect 29101 12597 29135 12631
rect 7849 12393 7883 12427
rect 9321 12393 9355 12427
rect 10609 12393 10643 12427
rect 11253 12393 11287 12427
rect 21649 12393 21683 12427
rect 27721 12393 27755 12427
rect 29837 12393 29871 12427
rect 7297 12325 7331 12359
rect 12449 12325 12483 12359
rect 18797 12325 18831 12359
rect 22845 12325 22879 12359
rect 24685 12325 24719 12359
rect 27077 12325 27111 12359
rect 13093 12257 13127 12291
rect 13737 12257 13771 12291
rect 15761 12257 15795 12291
rect 18245 12257 18279 12291
rect 20177 12257 20211 12291
rect 23397 12257 23431 12291
rect 7941 12189 7975 12223
rect 8585 12189 8619 12223
rect 9229 12189 9263 12223
rect 9873 12189 9907 12223
rect 10701 12189 10735 12223
rect 11345 12189 11379 12223
rect 17509 12189 17543 12223
rect 19441 12189 19475 12223
rect 22109 12189 22143 12223
rect 22293 12189 22327 12223
rect 26525 12189 26559 12223
rect 27169 12189 27203 12223
rect 27629 12189 27663 12223
rect 28457 12189 28491 12223
rect 29101 12189 29135 12223
rect 30297 12189 30331 12223
rect 9965 12121 9999 12155
rect 11897 12121 11931 12155
rect 11989 12121 12023 12155
rect 13185 12121 13219 12155
rect 14565 12121 14599 12155
rect 15117 12121 15151 12155
rect 15209 12121 15243 12155
rect 16681 12121 16715 12155
rect 16773 12121 16807 12155
rect 18337 12121 18371 12155
rect 20269 12121 20303 12155
rect 21189 12121 21223 12155
rect 23489 12121 23523 12155
rect 24041 12121 24075 12155
rect 25145 12121 25179 12155
rect 25237 12121 25271 12155
rect 25881 12121 25915 12155
rect 25973 12121 26007 12155
rect 29009 12121 29043 12155
rect 6653 12053 6687 12087
rect 8493 12053 8527 12087
rect 17601 12053 17635 12087
rect 19533 12053 19567 12087
rect 28365 12053 28399 12087
rect 7941 11849 7975 11883
rect 10425 11849 10459 11883
rect 11069 11849 11103 11883
rect 12173 11849 12207 11883
rect 28549 11849 28583 11883
rect 9873 11781 9907 11815
rect 12817 11781 12851 11815
rect 13369 11781 13403 11815
rect 14013 11781 14047 11815
rect 14933 11781 14967 11815
rect 15669 11781 15703 11815
rect 15761 11781 15795 11815
rect 18245 11781 18279 11815
rect 19073 11781 19107 11815
rect 20269 11781 20303 11815
rect 22201 11781 22235 11815
rect 23305 11781 23339 11815
rect 23857 11781 23891 11815
rect 24869 11781 24903 11815
rect 25421 11781 25455 11815
rect 26157 11781 26191 11815
rect 8401 11713 8435 11747
rect 9045 11713 9079 11747
rect 10517 11713 10551 11747
rect 11161 11713 11195 11747
rect 16313 11713 16347 11747
rect 17049 11713 17083 11747
rect 21373 11713 21407 11747
rect 21465 11713 21499 11747
rect 22753 11713 22787 11747
rect 26249 11713 26283 11747
rect 27353 11713 27387 11747
rect 27813 11713 27847 11747
rect 28457 11713 28491 11747
rect 37565 11713 37599 11747
rect 38209 11713 38243 11747
rect 12725 11645 12759 11679
rect 13921 11645 13955 11679
rect 17877 11645 17911 11679
rect 18337 11645 18371 11679
rect 18981 11645 19015 11679
rect 20177 11645 20211 11679
rect 20453 11645 20487 11679
rect 22109 11645 22143 11679
rect 23949 11645 23983 11679
rect 25513 11645 25547 11679
rect 29101 11645 29135 11679
rect 8493 11577 8527 11611
rect 19533 11577 19567 11611
rect 27905 11577 27939 11611
rect 38025 11577 38059 11611
rect 7297 11509 7331 11543
rect 9137 11509 9171 11543
rect 17141 11509 17175 11543
rect 27261 11509 27295 11543
rect 29653 11509 29687 11543
rect 11253 11305 11287 11339
rect 14289 11305 14323 11339
rect 16681 11237 16715 11271
rect 21189 11237 21223 11271
rect 24685 11237 24719 11271
rect 10425 11169 10459 11203
rect 12173 11169 12207 11203
rect 13093 11169 13127 11203
rect 14749 11169 14783 11203
rect 15485 11169 15519 11203
rect 16129 11169 16163 11203
rect 19901 11169 19935 11203
rect 20085 11169 20119 11203
rect 21833 11169 21867 11203
rect 23581 11169 23615 11203
rect 25237 11169 25271 11203
rect 25789 11169 25823 11203
rect 26433 11169 26467 11203
rect 27353 11169 27387 11203
rect 8033 11101 8067 11135
rect 9137 11101 9171 11135
rect 11345 11101 11379 11135
rect 13737 11101 13771 11135
rect 14933 11101 14967 11135
rect 18429 11101 18463 11135
rect 19441 11101 19475 11135
rect 28365 11101 28399 11135
rect 28825 11101 28859 11135
rect 29745 11101 29779 11135
rect 8585 11033 8619 11067
rect 9781 11033 9815 11067
rect 10333 11033 10367 11067
rect 11897 11033 11931 11067
rect 11989 11033 12023 11067
rect 13185 11033 13219 11067
rect 15577 11033 15611 11067
rect 18153 11033 18187 11067
rect 20637 11033 20671 11067
rect 20729 11033 20763 11067
rect 21925 11033 21959 11067
rect 22477 11033 22511 11067
rect 22937 11033 22971 11067
rect 23489 11033 23523 11067
rect 25145 11033 25179 11067
rect 26341 11033 26375 11067
rect 27077 11033 27111 11067
rect 27169 11033 27203 11067
rect 9229 10965 9263 10999
rect 28273 10965 28307 10999
rect 8769 10761 8803 10795
rect 21373 10761 21407 10795
rect 10425 10693 10459 10727
rect 12541 10693 12575 10727
rect 13369 10693 13403 10727
rect 13921 10693 13955 10727
rect 14565 10693 14599 10727
rect 15761 10693 15795 10727
rect 16313 10693 16347 10727
rect 24317 10693 24351 10727
rect 24869 10693 24903 10727
rect 25697 10693 25731 10727
rect 27353 10693 27387 10727
rect 1685 10625 1719 10659
rect 9689 10625 9723 10659
rect 10517 10625 10551 10659
rect 11161 10625 11195 10659
rect 11989 10625 12023 10659
rect 17233 10625 17267 10659
rect 19625 10625 19659 10659
rect 28917 10625 28951 10659
rect 37565 10625 37599 10659
rect 38209 10625 38243 10659
rect 12633 10557 12667 10591
rect 13277 10557 13311 10591
rect 14473 10557 14507 10591
rect 15669 10557 15703 10591
rect 17509 10557 17543 10591
rect 18981 10557 19015 10591
rect 19901 10557 19935 10591
rect 22017 10557 22051 10591
rect 22293 10557 22327 10591
rect 24961 10557 24995 10591
rect 25605 10557 25639 10591
rect 25881 10557 25915 10591
rect 27261 10557 27295 10591
rect 27905 10557 27939 10591
rect 28733 10557 28767 10591
rect 1869 10489 1903 10523
rect 9781 10489 9815 10523
rect 15025 10489 15059 10523
rect 29929 10489 29963 10523
rect 38025 10489 38059 10523
rect 8125 10421 8159 10455
rect 11069 10421 11103 10455
rect 23765 10421 23799 10455
rect 29377 10421 29411 10455
rect 1593 10217 1627 10251
rect 8585 10217 8619 10251
rect 23949 10217 23983 10251
rect 11161 10149 11195 10183
rect 13553 10149 13587 10183
rect 16313 10149 16347 10183
rect 26525 10149 26559 10183
rect 9873 10081 9907 10115
rect 12357 10081 12391 10115
rect 17049 10081 17083 10115
rect 17325 10081 17359 10115
rect 20729 10081 20763 10115
rect 21005 10081 21039 10115
rect 21649 10081 21683 10115
rect 9781 10013 9815 10047
rect 10617 10023 10651 10057
rect 11069 10013 11103 10047
rect 11713 10013 11747 10047
rect 14565 10013 14599 10047
rect 19441 10013 19475 10047
rect 27813 10013 27847 10047
rect 29009 10013 29043 10047
rect 30205 10013 30239 10047
rect 10517 9945 10551 9979
rect 12265 9945 12299 9979
rect 13001 9945 13035 9979
rect 13093 9945 13127 9979
rect 14841 9945 14875 9979
rect 20913 9945 20947 9979
rect 21925 9945 21959 9979
rect 24961 9945 24995 9979
rect 25053 9945 25087 9979
rect 25973 9945 26007 9979
rect 26985 9945 27019 9979
rect 27077 9945 27111 9979
rect 28733 9945 28767 9979
rect 29929 9945 29963 9979
rect 9321 9877 9355 9911
rect 18797 9877 18831 9911
rect 19533 9877 19567 9911
rect 23397 9877 23431 9911
rect 27721 9877 27755 9911
rect 14013 9673 14047 9707
rect 9781 9605 9815 9639
rect 10425 9605 10459 9639
rect 13001 9605 13035 9639
rect 17509 9605 17543 9639
rect 17601 9605 17635 9639
rect 21373 9605 21407 9639
rect 24409 9605 24443 9639
rect 24961 9605 24995 9639
rect 25513 9605 25547 9639
rect 27261 9605 27295 9639
rect 27905 9605 27939 9639
rect 28917 9605 28951 9639
rect 30849 9605 30883 9639
rect 10517 9537 10551 9571
rect 11161 9537 11195 9571
rect 11989 9537 12023 9571
rect 16957 9537 16991 9571
rect 20177 9537 20211 9571
rect 20637 9537 20671 9571
rect 21281 9537 21315 9571
rect 22017 9537 22051 9571
rect 24317 9537 24351 9571
rect 26341 9537 26375 9571
rect 27353 9537 27387 9571
rect 27997 9537 28031 9571
rect 34253 9537 34287 9571
rect 9321 9469 9355 9503
rect 13093 9469 13127 9503
rect 14473 9469 14507 9503
rect 16221 9469 16255 9503
rect 18153 9469 18187 9503
rect 19901 9469 19935 9503
rect 22293 9469 22327 9503
rect 25605 9469 25639 9503
rect 26249 9469 26283 9503
rect 28825 9469 28859 9503
rect 29101 9469 29135 9503
rect 31401 9469 31435 9503
rect 10977 9401 11011 9435
rect 12541 9401 12575 9435
rect 8769 9333 8803 9367
rect 11897 9333 11931 9367
rect 14736 9333 14770 9367
rect 20729 9333 20763 9367
rect 23765 9333 23799 9367
rect 30297 9333 30331 9367
rect 34345 9333 34379 9367
rect 11529 9129 11563 9163
rect 24685 9129 24719 9163
rect 30757 9129 30791 9163
rect 33517 9129 33551 9163
rect 19533 9061 19567 9095
rect 28825 9061 28859 9095
rect 1869 8993 1903 9027
rect 9781 8993 9815 9027
rect 12633 8993 12667 9027
rect 13645 8993 13679 9027
rect 16405 8993 16439 9027
rect 16865 8993 16899 9027
rect 18889 8993 18923 9027
rect 20269 8993 20303 9027
rect 23581 8993 23615 9027
rect 25789 8993 25823 9027
rect 26065 8993 26099 9027
rect 26985 8993 27019 9027
rect 27261 8993 27295 9027
rect 1593 8925 1627 8959
rect 10977 8925 11011 8959
rect 11437 8925 11471 8959
rect 13737 8925 13771 8959
rect 14381 8925 14415 8959
rect 19625 8925 19659 8959
rect 20177 8925 20211 8959
rect 20821 8925 20855 8959
rect 21557 8925 21591 8959
rect 24777 8925 24811 8959
rect 28089 8925 28123 8959
rect 28181 8925 28215 8959
rect 28917 8925 28951 8959
rect 30205 8925 30239 8959
rect 32505 8925 32539 8959
rect 32873 8925 32907 8959
rect 10333 8857 10367 8891
rect 12173 8857 12207 8891
rect 12265 8857 12299 8891
rect 14657 8857 14691 8891
rect 17141 8857 17175 8891
rect 20913 8857 20947 8891
rect 23305 8857 23339 8891
rect 25881 8857 25915 8891
rect 27077 8857 27111 8891
rect 29929 8857 29963 8891
rect 10885 8789 10919 8823
rect 1593 8585 1627 8619
rect 14013 8585 14047 8619
rect 24317 8585 24351 8619
rect 27905 8585 27939 8619
rect 29193 8585 29227 8619
rect 11161 8517 11195 8551
rect 14749 8517 14783 8551
rect 25053 8517 25087 8551
rect 25605 8517 25639 8551
rect 38025 8517 38059 8551
rect 2881 8449 2915 8483
rect 12265 8449 12299 8483
rect 17325 8449 17359 8483
rect 19993 8449 20027 8483
rect 20637 8449 20671 8483
rect 21189 8449 21223 8483
rect 21281 8449 21315 8483
rect 22017 8449 22051 8483
rect 26065 8449 26099 8483
rect 27353 8449 27387 8483
rect 27997 8449 28031 8483
rect 28641 8449 28675 8483
rect 29101 8449 29135 8483
rect 29929 8449 29963 8483
rect 30573 8449 30607 8483
rect 37565 8449 37599 8483
rect 38209 8449 38243 8483
rect 10609 8381 10643 8415
rect 11713 8381 11747 8415
rect 12541 8381 12575 8415
rect 14473 8381 14507 8415
rect 17969 8381 18003 8415
rect 18245 8381 18279 8415
rect 20545 8381 20579 8415
rect 22293 8381 22327 8415
rect 23765 8381 23799 8415
rect 24961 8381 24995 8415
rect 28549 8381 28583 8415
rect 29837 8381 29871 8415
rect 2789 8313 2823 8347
rect 16221 8313 16255 8347
rect 17509 8313 17543 8347
rect 27261 8313 27295 8347
rect 30481 8313 30515 8347
rect 26157 8245 26191 8279
rect 10885 8041 10919 8075
rect 12633 8041 12667 8075
rect 13277 8041 13311 8075
rect 16313 8041 16347 8075
rect 18797 8041 18831 8075
rect 24869 8041 24903 8075
rect 25513 8041 25547 8075
rect 26157 8041 26191 8075
rect 26801 8041 26835 8075
rect 28089 8041 28123 8075
rect 30481 8041 30515 8075
rect 29837 7973 29871 8007
rect 17049 7905 17083 7939
rect 19441 7905 19475 7939
rect 21741 7905 21775 7939
rect 28733 7905 28767 7939
rect 12725 7837 12759 7871
rect 13369 7837 13403 7871
rect 14565 7837 14599 7871
rect 24777 7837 24811 7871
rect 25605 7837 25639 7871
rect 26249 7837 26283 7871
rect 26893 7837 26927 7871
rect 27537 7837 27571 7871
rect 28181 7837 28215 7871
rect 28825 7837 28859 7871
rect 29929 7837 29963 7871
rect 30573 7837 30607 7871
rect 14841 7769 14875 7803
rect 17325 7769 17359 7803
rect 19717 7769 19751 7803
rect 22017 7769 22051 7803
rect 11437 7701 11471 7735
rect 11989 7701 12023 7735
rect 21189 7701 21223 7735
rect 23489 7701 23523 7735
rect 27445 7701 27479 7735
rect 13277 7497 13311 7531
rect 16957 7497 16991 7531
rect 17601 7497 17635 7531
rect 18245 7497 18279 7531
rect 23765 7497 23799 7531
rect 25697 7497 25731 7531
rect 26341 7497 26375 7531
rect 28549 7497 28583 7531
rect 29837 7497 29871 7531
rect 1869 7429 1903 7463
rect 10609 7429 10643 7463
rect 14749 7429 14783 7463
rect 27905 7429 27939 7463
rect 29193 7429 29227 7463
rect 1685 7361 1719 7395
rect 13369 7361 13403 7395
rect 17049 7361 17083 7395
rect 17509 7361 17543 7395
rect 18337 7361 18371 7395
rect 18797 7361 18831 7395
rect 21465 7361 21499 7395
rect 22017 7361 22051 7395
rect 24501 7361 24535 7395
rect 25145 7361 25179 7395
rect 25789 7361 25823 7395
rect 26433 7361 26467 7395
rect 27353 7361 27387 7395
rect 27997 7361 28031 7395
rect 28641 7361 28675 7395
rect 29285 7361 29319 7395
rect 29929 7361 29963 7395
rect 30573 7361 30607 7395
rect 14013 7293 14047 7327
rect 14473 7293 14507 7327
rect 19073 7293 19107 7327
rect 20545 7293 20579 7327
rect 22293 7293 22327 7327
rect 12725 7225 12759 7259
rect 24409 7225 24443 7259
rect 30481 7225 30515 7259
rect 11069 7157 11103 7191
rect 12081 7157 12115 7191
rect 16221 7157 16255 7191
rect 25053 7157 25087 7191
rect 27261 7157 27295 7191
rect 1593 6953 1627 6987
rect 17325 6885 17359 6919
rect 26709 6885 26743 6919
rect 10333 6817 10367 6851
rect 12265 6817 12299 6851
rect 15117 6817 15151 6851
rect 15577 6817 15611 6851
rect 17969 6817 18003 6851
rect 19533 6817 19567 6851
rect 20177 6817 20211 6851
rect 20729 6817 20763 6851
rect 21189 6817 21223 6851
rect 21465 6817 21499 6851
rect 22937 6817 22971 6851
rect 24961 6817 24995 6851
rect 29101 6817 29135 6851
rect 11989 6749 12023 6783
rect 18889 6749 18923 6783
rect 19625 6749 19659 6783
rect 24041 6749 24075 6783
rect 24877 6749 24911 6783
rect 25605 6749 25639 6783
rect 25697 6749 25731 6783
rect 26801 6749 26835 6783
rect 27445 6749 27479 6783
rect 28089 6749 28123 6783
rect 29193 6749 29227 6783
rect 15853 6681 15887 6715
rect 10977 6613 11011 6647
rect 11437 6613 11471 6647
rect 13737 6613 13771 6647
rect 14565 6613 14599 6647
rect 23949 6613 23983 6647
rect 27353 6613 27387 6647
rect 27997 6613 28031 6647
rect 20637 6409 20671 6443
rect 10609 6341 10643 6375
rect 14841 6341 14875 6375
rect 27905 6341 27939 6375
rect 38025 6341 38059 6375
rect 17233 6273 17267 6307
rect 17785 6273 17819 6307
rect 24961 6273 24995 6307
rect 26157 6273 26191 6307
rect 26249 6273 26283 6307
rect 27261 6273 27295 6307
rect 27353 6273 27387 6307
rect 27997 6273 28031 6307
rect 37565 6273 37599 6307
rect 38209 6273 38243 6307
rect 11897 6205 11931 6239
rect 12357 6205 12391 6239
rect 12633 6205 12667 6239
rect 14565 6205 14599 6239
rect 16313 6205 16347 6239
rect 18061 6205 18095 6239
rect 19533 6205 19567 6239
rect 22109 6205 22143 6239
rect 23581 6205 23615 6239
rect 23857 6205 23891 6239
rect 28549 6137 28583 6171
rect 29101 6137 29135 6171
rect 29653 6137 29687 6171
rect 9965 6069 9999 6103
rect 11069 6069 11103 6103
rect 14105 6069 14139 6103
rect 21097 6069 21131 6103
rect 24869 6069 24903 6103
rect 25421 6069 25455 6103
rect 30113 6069 30147 6103
rect 10425 5865 10459 5899
rect 20361 5865 20395 5899
rect 21005 5865 21039 5899
rect 23305 5865 23339 5899
rect 27905 5865 27939 5899
rect 16681 5797 16715 5831
rect 19717 5797 19751 5831
rect 13737 5729 13771 5763
rect 14473 5729 14507 5763
rect 14933 5729 14967 5763
rect 15209 5729 15243 5763
rect 17141 5729 17175 5763
rect 18889 5729 18923 5763
rect 21557 5729 21591 5763
rect 26709 5729 26743 5763
rect 24593 5661 24627 5695
rect 24685 5661 24719 5695
rect 25881 5661 25915 5695
rect 26801 5661 26835 5695
rect 28917 5661 28951 5695
rect 11437 5593 11471 5627
rect 13461 5593 13495 5627
rect 17417 5593 17451 5627
rect 21833 5593 21867 5627
rect 28825 5593 28859 5627
rect 9873 5525 9907 5559
rect 10977 5525 11011 5559
rect 11989 5525 12023 5559
rect 23857 5525 23891 5559
rect 25789 5525 25823 5559
rect 27261 5525 27295 5559
rect 29837 5525 29871 5559
rect 30389 5525 30423 5559
rect 30849 5525 30883 5559
rect 14105 5321 14139 5355
rect 27261 5321 27295 5355
rect 31217 5321 31251 5355
rect 12633 5253 12667 5287
rect 14841 5253 14875 5287
rect 30113 5253 30147 5287
rect 1869 5185 1903 5219
rect 12357 5185 12391 5219
rect 14565 5185 14599 5219
rect 16957 5185 16991 5219
rect 17417 5185 17451 5219
rect 26525 5185 26559 5219
rect 27353 5185 27387 5219
rect 27997 5185 28031 5219
rect 28917 5185 28951 5219
rect 29561 5185 29595 5219
rect 30205 5185 30239 5219
rect 9505 5117 9539 5151
rect 17693 5117 17727 5151
rect 19625 5117 19659 5151
rect 19901 5117 19935 5151
rect 22017 5117 22051 5151
rect 22293 5117 22327 5151
rect 29469 5117 29503 5151
rect 38025 5117 38059 5151
rect 38301 5117 38335 5151
rect 27905 5049 27939 5083
rect 30757 5049 30791 5083
rect 1685 4981 1719 5015
rect 9965 4981 9999 5015
rect 10517 4981 10551 5015
rect 11069 4981 11103 5015
rect 11897 4981 11931 5015
rect 16313 4981 16347 5015
rect 19165 4981 19199 5015
rect 21373 4981 21407 5015
rect 23765 4981 23799 5015
rect 24317 4981 24351 5015
rect 24777 4981 24811 5015
rect 25329 4981 25363 5015
rect 26433 4981 26467 5015
rect 28825 4981 28859 5015
rect 11437 4777 11471 4811
rect 18889 4777 18923 4811
rect 19533 4777 19567 4811
rect 20821 4777 20855 4811
rect 23673 4777 23707 4811
rect 24685 4777 24719 4811
rect 25237 4777 25271 4811
rect 25789 4777 25823 4811
rect 26341 4777 26375 4811
rect 27721 4777 27755 4811
rect 29101 4777 29135 4811
rect 33057 4777 33091 4811
rect 38301 4777 38335 4811
rect 29837 4709 29871 4743
rect 11989 4641 12023 4675
rect 12265 4641 12299 4675
rect 13737 4641 13771 4675
rect 16405 4641 16439 4675
rect 17141 4641 17175 4675
rect 20085 4641 20119 4675
rect 23121 4641 23155 4675
rect 31033 4641 31067 4675
rect 9873 4573 9907 4607
rect 27077 4573 27111 4607
rect 27169 4573 27203 4607
rect 28457 4573 28491 4607
rect 29193 4573 29227 4607
rect 29929 4573 29963 4607
rect 30573 4573 30607 4607
rect 32229 4573 32263 4607
rect 32505 4573 32539 4607
rect 16129 4505 16163 4539
rect 17417 4505 17451 4539
rect 22845 4505 22879 4539
rect 30481 4505 30515 4539
rect 9321 4437 9355 4471
rect 10425 4437 10459 4471
rect 10977 4437 11011 4471
rect 14657 4437 14691 4471
rect 21373 4437 21407 4471
rect 28273 4437 28307 4471
rect 10057 4233 10091 4267
rect 11069 4233 11103 4267
rect 12081 4233 12115 4267
rect 21373 4233 21407 4267
rect 13553 4165 13587 4199
rect 16313 4165 16347 4199
rect 24501 4165 24535 4199
rect 16865 4097 16899 4131
rect 23765 4097 23799 4131
rect 24225 4097 24259 4131
rect 27537 4097 27571 4131
rect 27629 4097 27663 4131
rect 28273 4097 28307 4131
rect 29193 4097 29227 4131
rect 29285 4097 29319 4131
rect 29929 4097 29963 4131
rect 30389 4097 30423 4131
rect 31217 4097 31251 4131
rect 32321 4097 32355 4131
rect 33241 4097 33275 4131
rect 13829 4029 13863 4063
rect 14289 4029 14323 4063
rect 14565 4029 14599 4063
rect 17141 4029 17175 4063
rect 18613 4029 18647 4063
rect 18889 4029 18923 4063
rect 20637 4029 20671 4063
rect 22017 4029 22051 4063
rect 23489 4029 23523 4063
rect 31677 4029 31711 4063
rect 32505 4029 32539 4063
rect 26525 3961 26559 3995
rect 30481 3961 30515 3995
rect 31125 3961 31159 3995
rect 8309 3893 8343 3927
rect 8861 3893 8895 3927
rect 9413 3893 9447 3927
rect 10609 3893 10643 3927
rect 25973 3893 26007 3927
rect 28181 3893 28215 3927
rect 29837 3893 29871 3927
rect 9229 3689 9263 3723
rect 20269 3689 20303 3723
rect 28825 3689 28859 3723
rect 32413 3689 32447 3723
rect 34897 3689 34931 3723
rect 4813 3621 4847 3655
rect 13737 3621 13771 3655
rect 26341 3621 26375 3655
rect 26985 3621 27019 3655
rect 38025 3621 38059 3655
rect 8585 3553 8619 3587
rect 12265 3553 12299 3587
rect 14933 3553 14967 3587
rect 16865 3553 16899 3587
rect 21005 3553 21039 3587
rect 24593 3553 24627 3587
rect 24869 3553 24903 3587
rect 29837 3553 29871 3587
rect 32965 3553 32999 3587
rect 1593 3485 1627 3519
rect 2237 3485 2271 3519
rect 11437 3485 11471 3519
rect 11529 3485 11563 3519
rect 11989 3485 12023 3519
rect 14657 3485 14691 3519
rect 19441 3485 19475 3519
rect 20453 3485 20487 3519
rect 23765 3485 23799 3519
rect 26801 3485 26835 3519
rect 27537 3485 27571 3519
rect 27629 3485 27663 3519
rect 28273 3485 28307 3519
rect 28925 3485 28959 3519
rect 29929 3485 29963 3519
rect 30573 3485 30607 3519
rect 31125 3485 31159 3519
rect 31217 3485 31251 3519
rect 31861 3485 31895 3519
rect 32505 3485 32539 3519
rect 17141 3417 17175 3451
rect 18889 3417 18923 3451
rect 21281 3417 21315 3451
rect 23029 3417 23063 3451
rect 37565 3417 37599 3451
rect 38209 3417 38243 3451
rect 1777 3349 1811 3383
rect 7481 3349 7515 3383
rect 8033 3349 8067 3383
rect 9781 3349 9815 3383
rect 10241 3349 10275 3383
rect 10793 3349 10827 3383
rect 16405 3349 16439 3383
rect 19625 3349 19659 3383
rect 23581 3349 23615 3383
rect 28181 3349 28215 3383
rect 30481 3349 30515 3383
rect 31769 3349 31803 3383
rect 33609 3349 33643 3383
rect 34069 3349 34103 3383
rect 2789 3145 2823 3179
rect 3341 3145 3375 3179
rect 7205 3145 7239 3179
rect 11805 3145 11839 3179
rect 16313 3145 16347 3179
rect 32413 3145 32447 3179
rect 10333 3077 10367 3111
rect 12633 3077 12667 3111
rect 14841 3077 14875 3111
rect 19717 3077 19751 3111
rect 33057 3077 33091 3111
rect 1869 3009 1903 3043
rect 4445 3009 4479 3043
rect 5273 3009 5307 3043
rect 9321 3009 9355 3043
rect 9413 3009 9447 3043
rect 10885 3009 10919 3043
rect 11713 3009 11747 3043
rect 12357 3009 12391 3043
rect 17233 3009 17267 3043
rect 19441 3009 19475 3043
rect 24041 3009 24075 3043
rect 26249 3009 26283 3043
rect 27445 3009 27479 3043
rect 28089 3009 28123 3043
rect 28549 3009 28583 3043
rect 29193 3009 29227 3043
rect 29837 3009 29871 3043
rect 30665 3009 30699 3043
rect 31309 3009 31343 3043
rect 32505 3009 32539 3043
rect 32965 3009 32999 3043
rect 33609 3009 33643 3043
rect 38025 3009 38059 3043
rect 8861 2941 8895 2975
rect 14105 2941 14139 2975
rect 14565 2941 14599 2975
rect 17509 2941 17543 2975
rect 18981 2941 19015 2975
rect 21465 2941 21499 2975
rect 22017 2941 22051 2975
rect 23765 2941 23799 2975
rect 24501 2941 24535 2975
rect 25973 2941 26007 2975
rect 34253 2941 34287 2975
rect 35357 2941 35391 2975
rect 5089 2873 5123 2907
rect 6653 2873 6687 2907
rect 33793 2873 33827 2907
rect 1685 2805 1719 2839
rect 4629 2805 4663 2839
rect 7757 2805 7791 2839
rect 8217 2805 8251 2839
rect 11069 2805 11103 2839
rect 27261 2805 27295 2839
rect 27905 2805 27939 2839
rect 28733 2805 28767 2839
rect 29285 2805 29319 2839
rect 29929 2805 29963 2839
rect 30573 2805 30607 2839
rect 31217 2805 31251 2839
rect 34805 2805 34839 2839
rect 35909 2805 35943 2839
rect 38209 2805 38243 2839
rect 3249 2601 3283 2635
rect 7481 2601 7515 2635
rect 8033 2601 8067 2635
rect 10057 2601 10091 2635
rect 11989 2601 12023 2635
rect 14822 2601 14856 2635
rect 27997 2601 28031 2635
rect 32965 2601 32999 2635
rect 34161 2601 34195 2635
rect 2421 2533 2455 2567
rect 10885 2533 10919 2567
rect 24593 2533 24627 2567
rect 35633 2533 35667 2567
rect 13737 2465 13771 2499
rect 14565 2465 14599 2499
rect 17141 2465 17175 2499
rect 19717 2465 19751 2499
rect 22293 2465 22327 2499
rect 26341 2465 26375 2499
rect 29837 2465 29871 2499
rect 1869 2397 1903 2431
rect 2605 2397 2639 2431
rect 3341 2397 3375 2431
rect 3985 2397 4019 2431
rect 4905 2397 4939 2431
rect 6837 2397 6871 2431
rect 9873 2397 9907 2431
rect 11069 2397 11103 2431
rect 19441 2397 19475 2431
rect 22017 2397 22051 2431
rect 27445 2397 27479 2431
rect 28825 2397 28859 2431
rect 29745 2397 29779 2431
rect 30665 2397 30699 2431
rect 31309 2397 31343 2431
rect 32321 2397 32355 2431
rect 33149 2397 33183 2431
rect 34897 2397 34931 2431
rect 36645 2397 36679 2431
rect 37473 2397 37507 2431
rect 6009 2329 6043 2363
rect 9229 2329 9263 2363
rect 13461 2329 13495 2363
rect 17417 2329 17451 2363
rect 21465 2329 21499 2363
rect 26065 2329 26099 2363
rect 28089 2329 28123 2363
rect 35817 2329 35851 2363
rect 1685 2261 1719 2295
rect 4721 2261 4755 2295
rect 6653 2261 6687 2295
rect 8585 2261 8619 2295
rect 9321 2261 9355 2295
rect 16313 2261 16347 2295
rect 18889 2261 18923 2295
rect 23765 2261 23799 2295
rect 27261 2261 27295 2295
rect 28733 2261 28767 2295
rect 30481 2261 30515 2295
rect 31125 2261 31159 2295
rect 32505 2261 32539 2295
rect 33609 2261 33643 2295
rect 35081 2261 35115 2295
rect 36829 2261 36863 2295
rect 37657 2261 37691 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 17681 37451 17739 37457
rect 17681 37417 17693 37451
rect 17727 37448 17739 37451
rect 18046 37448 18052 37460
rect 17727 37420 18052 37448
rect 17727 37417 17739 37420
rect 17681 37411 17739 37417
rect 18046 37408 18052 37420
rect 18104 37408 18110 37460
rect 12437 37315 12495 37321
rect 12437 37281 12449 37315
rect 12483 37281 12495 37315
rect 12437 37275 12495 37281
rect 14461 37315 14519 37321
rect 14461 37281 14473 37315
rect 14507 37312 14519 37315
rect 14826 37312 14832 37324
rect 14507 37284 14832 37312
rect 14507 37281 14519 37284
rect 14461 37275 14519 37281
rect 1857 37247 1915 37253
rect 1857 37213 1869 37247
rect 1903 37244 1915 37247
rect 2314 37244 2320 37256
rect 1903 37216 2320 37244
rect 1903 37213 1915 37216
rect 1857 37207 1915 37213
rect 2314 37204 2320 37216
rect 2372 37204 2378 37256
rect 2961 37247 3019 37253
rect 2961 37213 2973 37247
rect 3007 37213 3019 37247
rect 2961 37207 3019 37213
rect 4893 37247 4951 37253
rect 4893 37213 4905 37247
rect 4939 37244 4951 37247
rect 5442 37244 5448 37256
rect 4939 37216 5448 37244
rect 4939 37213 4951 37216
rect 4893 37207 4951 37213
rect 2976 37176 3004 37207
rect 5442 37204 5448 37216
rect 5500 37204 5506 37256
rect 6825 37247 6883 37253
rect 6825 37213 6837 37247
rect 6871 37244 6883 37247
rect 7282 37244 7288 37256
rect 6871 37216 7288 37244
rect 6871 37213 6883 37216
rect 6825 37207 6883 37213
rect 7282 37204 7288 37216
rect 7340 37204 7346 37256
rect 7377 37247 7435 37253
rect 7377 37213 7389 37247
rect 7423 37244 7435 37247
rect 7742 37244 7748 37256
rect 7423 37216 7748 37244
rect 7423 37213 7435 37216
rect 7377 37207 7435 37213
rect 7742 37204 7748 37216
rect 7800 37244 7806 37256
rect 7929 37247 7987 37253
rect 7929 37244 7941 37247
rect 7800 37216 7941 37244
rect 7800 37204 7806 37216
rect 7929 37213 7941 37216
rect 7975 37213 7987 37247
rect 7929 37207 7987 37213
rect 10045 37247 10103 37253
rect 10045 37213 10057 37247
rect 10091 37213 10103 37247
rect 10045 37207 10103 37213
rect 11977 37247 12035 37253
rect 11977 37213 11989 37247
rect 12023 37244 12035 37247
rect 12066 37244 12072 37256
rect 12023 37216 12072 37244
rect 12023 37213 12035 37216
rect 11977 37207 12035 37213
rect 6730 37176 6736 37188
rect 2976 37148 6736 37176
rect 6730 37136 6736 37148
rect 6788 37136 6794 37188
rect 10060 37176 10088 37207
rect 12066 37204 12072 37216
rect 12124 37244 12130 37256
rect 12452 37244 12480 37275
rect 14826 37272 14832 37284
rect 14884 37312 14890 37324
rect 14921 37315 14979 37321
rect 14921 37312 14933 37315
rect 14884 37284 14933 37312
rect 14884 37272 14890 37284
rect 14921 37281 14933 37284
rect 14967 37281 14979 37315
rect 14921 37275 14979 37281
rect 16301 37315 16359 37321
rect 16301 37281 16313 37315
rect 16347 37312 16359 37315
rect 16666 37312 16672 37324
rect 16347 37284 16672 37312
rect 16347 37281 16359 37284
rect 16301 37275 16359 37281
rect 16666 37272 16672 37284
rect 16724 37272 16730 37324
rect 16758 37272 16764 37324
rect 16816 37312 16822 37324
rect 17129 37315 17187 37321
rect 17129 37312 17141 37315
rect 16816 37284 17141 37312
rect 16816 37272 16822 37284
rect 17129 37281 17141 37284
rect 17175 37281 17187 37315
rect 18138 37312 18144 37324
rect 18099 37284 18144 37312
rect 17129 37275 17187 37281
rect 18138 37272 18144 37284
rect 18196 37272 18202 37324
rect 21453 37315 21511 37321
rect 21453 37281 21465 37315
rect 21499 37312 21511 37315
rect 21910 37312 21916 37324
rect 21499 37284 21916 37312
rect 21499 37281 21511 37284
rect 21453 37275 21511 37281
rect 21910 37272 21916 37284
rect 21968 37312 21974 37324
rect 22005 37315 22063 37321
rect 22005 37312 22017 37315
rect 21968 37284 22017 37312
rect 21968 37272 21974 37284
rect 22005 37281 22017 37284
rect 22051 37281 22063 37315
rect 22005 37275 22063 37281
rect 35069 37315 35127 37321
rect 35069 37281 35081 37315
rect 35115 37312 35127 37315
rect 35434 37312 35440 37324
rect 35115 37284 35440 37312
rect 35115 37281 35127 37284
rect 35069 37275 35127 37281
rect 35434 37272 35440 37284
rect 35492 37312 35498 37324
rect 35529 37315 35587 37321
rect 35529 37312 35541 37315
rect 35492 37284 35541 37312
rect 35492 37272 35498 37284
rect 35529 37281 35541 37284
rect 35575 37281 35587 37315
rect 35529 37275 35587 37281
rect 36909 37315 36967 37321
rect 36909 37281 36921 37315
rect 36955 37312 36967 37315
rect 38286 37312 38292 37324
rect 36955 37284 38292 37312
rect 36955 37281 36967 37284
rect 36909 37275 36967 37281
rect 38286 37272 38292 37284
rect 38344 37272 38350 37324
rect 13262 37244 13268 37256
rect 12124 37216 12480 37244
rect 13223 37216 13268 37244
rect 12124 37204 12130 37216
rect 13262 37204 13268 37216
rect 13320 37204 13326 37256
rect 13354 37204 13360 37256
rect 13412 37244 13418 37256
rect 15197 37247 15255 37253
rect 15197 37244 15209 37247
rect 13412 37216 15209 37244
rect 13412 37204 13418 37216
rect 15197 37213 15209 37216
rect 15243 37213 15255 37247
rect 16684 37244 16712 37272
rect 16945 37247 17003 37253
rect 16945 37244 16957 37247
rect 16684 37216 16957 37244
rect 15197 37207 15255 37213
rect 16945 37213 16957 37216
rect 16991 37213 17003 37247
rect 16945 37207 17003 37213
rect 18046 37204 18052 37256
rect 18104 37244 18110 37256
rect 18325 37247 18383 37253
rect 18325 37244 18337 37247
rect 18104 37216 18337 37244
rect 18104 37204 18110 37216
rect 18325 37213 18337 37216
rect 18371 37213 18383 37247
rect 20070 37244 20076 37256
rect 20031 37216 20076 37244
rect 18325 37207 18383 37213
rect 20070 37204 20076 37216
rect 20128 37204 20134 37256
rect 20530 37204 20536 37256
rect 20588 37244 20594 37256
rect 22281 37247 22339 37253
rect 22281 37244 22293 37247
rect 20588 37216 22293 37244
rect 20588 37204 20594 37216
rect 22281 37213 22293 37216
rect 22327 37244 22339 37247
rect 23014 37244 23020 37256
rect 22327 37216 23020 37244
rect 22327 37213 22339 37216
rect 22281 37207 22339 37213
rect 23014 37204 23020 37216
rect 23072 37204 23078 37256
rect 23290 37244 23296 37256
rect 23251 37216 23296 37244
rect 23290 37204 23296 37216
rect 23348 37204 23354 37256
rect 25225 37247 25283 37253
rect 25225 37213 25237 37247
rect 25271 37213 25283 37247
rect 25225 37207 25283 37213
rect 13170 37176 13176 37188
rect 10060 37148 13176 37176
rect 13170 37136 13176 37148
rect 13228 37136 13234 37188
rect 20714 37136 20720 37188
rect 20772 37176 20778 37188
rect 25240 37176 25268 37207
rect 25866 37204 25872 37256
rect 25924 37244 25930 37256
rect 27157 37247 27215 37253
rect 27157 37244 27169 37247
rect 25924 37216 27169 37244
rect 25924 37204 25930 37216
rect 27157 37213 27169 37216
rect 27203 37213 27215 37247
rect 27157 37207 27215 37213
rect 27430 37204 27436 37256
rect 27488 37244 27494 37256
rect 28445 37247 28503 37253
rect 28445 37244 28457 37247
rect 27488 37216 28457 37244
rect 27488 37204 27494 37216
rect 28445 37213 28457 37216
rect 28491 37213 28503 37247
rect 28445 37207 28503 37213
rect 30377 37247 30435 37253
rect 30377 37213 30389 37247
rect 30423 37244 30435 37247
rect 30466 37244 30472 37256
rect 30423 37216 30472 37244
rect 30423 37213 30435 37216
rect 30377 37207 30435 37213
rect 30466 37204 30472 37216
rect 30524 37204 30530 37256
rect 30834 37204 30840 37256
rect 30892 37244 30898 37256
rect 32309 37247 32367 37253
rect 32309 37244 32321 37247
rect 30892 37216 32321 37244
rect 30892 37204 30898 37216
rect 32309 37213 32321 37216
rect 32355 37213 32367 37247
rect 33594 37244 33600 37256
rect 33555 37216 33600 37244
rect 32309 37207 32367 37213
rect 33594 37204 33600 37216
rect 33652 37204 33658 37256
rect 35802 37244 35808 37256
rect 35763 37216 35808 37244
rect 35802 37204 35808 37216
rect 35860 37204 35866 37256
rect 37826 37204 37832 37256
rect 37884 37244 37890 37256
rect 38013 37247 38071 37253
rect 38013 37244 38025 37247
rect 37884 37216 38025 37244
rect 37884 37204 37890 37216
rect 38013 37213 38025 37216
rect 38059 37213 38071 37247
rect 38013 37207 38071 37213
rect 20772 37148 25268 37176
rect 20772 37136 20778 37148
rect 1302 37068 1308 37120
rect 1360 37108 1366 37120
rect 1673 37111 1731 37117
rect 1673 37108 1685 37111
rect 1360 37080 1685 37108
rect 1360 37068 1366 37080
rect 1673 37077 1685 37080
rect 1719 37077 1731 37111
rect 2774 37108 2780 37120
rect 2735 37080 2780 37108
rect 1673 37071 1731 37077
rect 2774 37068 2780 37080
rect 2832 37068 2838 37120
rect 4614 37068 4620 37120
rect 4672 37108 4678 37120
rect 4709 37111 4767 37117
rect 4709 37108 4721 37111
rect 4672 37080 4721 37108
rect 4672 37068 4678 37080
rect 4709 37077 4721 37080
rect 4755 37077 4767 37111
rect 5442 37108 5448 37120
rect 5403 37080 5448 37108
rect 4709 37071 4767 37077
rect 5442 37068 5448 37080
rect 5500 37068 5506 37120
rect 6454 37068 6460 37120
rect 6512 37108 6518 37120
rect 6641 37111 6699 37117
rect 6641 37108 6653 37111
rect 6512 37080 6653 37108
rect 6512 37068 6518 37080
rect 6641 37077 6653 37080
rect 6687 37077 6699 37111
rect 8018 37108 8024 37120
rect 7979 37080 8024 37108
rect 6641 37071 6699 37077
rect 8018 37068 8024 37080
rect 8076 37068 8082 37120
rect 9674 37068 9680 37120
rect 9732 37108 9738 37120
rect 9861 37111 9919 37117
rect 9861 37108 9873 37111
rect 9732 37080 9873 37108
rect 9732 37068 9738 37080
rect 9861 37077 9873 37080
rect 9907 37077 9919 37111
rect 9861 37071 9919 37077
rect 11606 37068 11612 37120
rect 11664 37108 11670 37120
rect 11793 37111 11851 37117
rect 11793 37108 11805 37111
rect 11664 37080 11805 37108
rect 11664 37068 11670 37080
rect 11793 37077 11805 37080
rect 11839 37077 11851 37111
rect 11793 37071 11851 37077
rect 12894 37068 12900 37120
rect 12952 37108 12958 37120
rect 13081 37111 13139 37117
rect 13081 37108 13093 37111
rect 12952 37080 13093 37108
rect 12952 37068 12958 37080
rect 13081 37077 13093 37080
rect 13127 37077 13139 37111
rect 13081 37071 13139 37077
rect 19978 37068 19984 37120
rect 20036 37108 20042 37120
rect 20257 37111 20315 37117
rect 20257 37108 20269 37111
rect 20036 37080 20269 37108
rect 20036 37068 20042 37080
rect 20257 37077 20269 37080
rect 20303 37077 20315 37111
rect 20257 37071 20315 37077
rect 23198 37068 23204 37120
rect 23256 37108 23262 37120
rect 23477 37111 23535 37117
rect 23477 37108 23489 37111
rect 23256 37080 23489 37108
rect 23256 37068 23262 37080
rect 23477 37077 23489 37080
rect 23523 37077 23535 37111
rect 23477 37071 23535 37077
rect 25130 37068 25136 37120
rect 25188 37108 25194 37120
rect 25409 37111 25467 37117
rect 25409 37108 25421 37111
rect 25188 37080 25421 37108
rect 25188 37068 25194 37080
rect 25409 37077 25421 37080
rect 25455 37077 25467 37111
rect 25409 37071 25467 37077
rect 27062 37068 27068 37120
rect 27120 37108 27126 37120
rect 27341 37111 27399 37117
rect 27341 37108 27353 37111
rect 27120 37080 27353 37108
rect 27120 37068 27126 37080
rect 27341 37077 27353 37080
rect 27387 37077 27399 37111
rect 27341 37071 27399 37077
rect 28350 37068 28356 37120
rect 28408 37108 28414 37120
rect 28629 37111 28687 37117
rect 28629 37108 28641 37111
rect 28408 37080 28641 37108
rect 28408 37068 28414 37080
rect 28629 37077 28641 37080
rect 28675 37077 28687 37111
rect 28629 37071 28687 37077
rect 30374 37068 30380 37120
rect 30432 37108 30438 37120
rect 30561 37111 30619 37117
rect 30561 37108 30573 37111
rect 30432 37080 30573 37108
rect 30432 37068 30438 37080
rect 30561 37077 30573 37080
rect 30607 37077 30619 37111
rect 30561 37071 30619 37077
rect 32214 37068 32220 37120
rect 32272 37108 32278 37120
rect 32493 37111 32551 37117
rect 32493 37108 32505 37111
rect 32272 37080 32505 37108
rect 32272 37068 32278 37080
rect 32493 37077 32505 37080
rect 32539 37077 32551 37111
rect 32493 37071 32551 37077
rect 33502 37068 33508 37120
rect 33560 37108 33566 37120
rect 33781 37111 33839 37117
rect 33781 37108 33793 37111
rect 33560 37080 33793 37108
rect 33560 37068 33566 37080
rect 33781 37077 33793 37080
rect 33827 37077 33839 37111
rect 33781 37071 33839 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 5442 36864 5448 36916
rect 5500 36904 5506 36916
rect 22094 36904 22100 36916
rect 5500 36876 22100 36904
rect 5500 36864 5506 36876
rect 22094 36864 22100 36876
rect 22152 36864 22158 36916
rect 22189 36907 22247 36913
rect 22189 36873 22201 36907
rect 22235 36904 22247 36907
rect 23290 36904 23296 36916
rect 22235 36876 23296 36904
rect 22235 36873 22247 36876
rect 22189 36867 22247 36873
rect 23290 36864 23296 36876
rect 23348 36864 23354 36916
rect 27985 36907 28043 36913
rect 27985 36873 27997 36907
rect 28031 36904 28043 36907
rect 33594 36904 33600 36916
rect 28031 36876 33600 36904
rect 28031 36873 28043 36876
rect 27985 36867 28043 36873
rect 33594 36864 33600 36876
rect 33652 36864 33658 36916
rect 37366 36864 37372 36916
rect 37424 36904 37430 36916
rect 37553 36907 37611 36913
rect 37553 36904 37565 36907
rect 37424 36876 37565 36904
rect 37424 36864 37430 36876
rect 37553 36873 37565 36876
rect 37599 36873 37611 36907
rect 37553 36867 37611 36873
rect 2409 36839 2467 36845
rect 2409 36805 2421 36839
rect 2455 36836 2467 36839
rect 2866 36836 2872 36848
rect 2455 36808 2872 36836
rect 2455 36805 2467 36808
rect 2409 36799 2467 36805
rect 2866 36796 2872 36808
rect 2924 36796 2930 36848
rect 1673 36771 1731 36777
rect 1673 36737 1685 36771
rect 1719 36768 1731 36771
rect 2958 36768 2964 36780
rect 1719 36740 2964 36768
rect 1719 36737 1731 36740
rect 1673 36731 1731 36737
rect 2958 36728 2964 36740
rect 3016 36768 3022 36780
rect 3053 36771 3111 36777
rect 3053 36768 3065 36771
rect 3016 36740 3065 36768
rect 3016 36728 3022 36740
rect 3053 36737 3065 36740
rect 3099 36737 3111 36771
rect 3053 36731 3111 36737
rect 10597 36771 10655 36777
rect 10597 36737 10609 36771
rect 10643 36768 10655 36771
rect 13354 36768 13360 36780
rect 10643 36740 13360 36768
rect 10643 36737 10655 36740
rect 10597 36731 10655 36737
rect 13354 36728 13360 36740
rect 13412 36728 13418 36780
rect 22005 36771 22063 36777
rect 22005 36737 22017 36771
rect 22051 36768 22063 36771
rect 22278 36768 22284 36780
rect 22051 36740 22284 36768
rect 22051 36737 22063 36740
rect 22005 36731 22063 36737
rect 22278 36728 22284 36740
rect 22336 36768 22342 36780
rect 22738 36768 22744 36780
rect 22336 36740 22744 36768
rect 22336 36728 22342 36740
rect 22738 36728 22744 36740
rect 22796 36728 22802 36780
rect 23014 36728 23020 36780
rect 23072 36768 23078 36780
rect 27801 36771 27859 36777
rect 27801 36768 27813 36771
rect 23072 36740 27813 36768
rect 23072 36728 23078 36740
rect 27801 36737 27813 36740
rect 27847 36737 27859 36771
rect 27801 36731 27859 36737
rect 36725 36771 36783 36777
rect 36725 36737 36737 36771
rect 36771 36737 36783 36771
rect 37734 36768 37740 36780
rect 37647 36740 37740 36768
rect 36725 36731 36783 36737
rect 36740 36700 36768 36731
rect 37734 36728 37740 36740
rect 37792 36768 37798 36780
rect 38197 36771 38255 36777
rect 38197 36768 38209 36771
rect 37792 36740 38209 36768
rect 37792 36728 37798 36740
rect 38197 36737 38209 36740
rect 38243 36737 38255 36771
rect 38197 36731 38255 36737
rect 37918 36700 37924 36712
rect 36740 36672 37924 36700
rect 37918 36660 37924 36672
rect 37976 36660 37982 36712
rect 1857 36635 1915 36641
rect 1857 36601 1869 36635
rect 1903 36632 1915 36635
rect 16298 36632 16304 36644
rect 1903 36604 16304 36632
rect 1903 36601 1915 36604
rect 1857 36595 1915 36601
rect 16298 36592 16304 36604
rect 16356 36592 16362 36644
rect 2498 36564 2504 36576
rect 2459 36536 2504 36564
rect 2498 36524 2504 36536
rect 2556 36524 2562 36576
rect 7282 36524 7288 36576
rect 7340 36564 7346 36576
rect 10413 36567 10471 36573
rect 10413 36564 10425 36567
rect 7340 36536 10425 36564
rect 7340 36524 7346 36536
rect 10413 36533 10425 36536
rect 10459 36533 10471 36567
rect 22738 36564 22744 36576
rect 22699 36536 22744 36564
rect 10413 36527 10471 36533
rect 22738 36524 22744 36536
rect 22796 36524 22802 36576
rect 36909 36567 36967 36573
rect 36909 36533 36921 36567
rect 36955 36564 36967 36567
rect 38010 36564 38016 36576
rect 36955 36536 38016 36564
rect 36955 36533 36967 36536
rect 36909 36527 36967 36533
rect 38010 36524 38016 36536
rect 38068 36524 38074 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 2409 36363 2467 36369
rect 2409 36329 2421 36363
rect 2455 36360 2467 36363
rect 2866 36360 2872 36372
rect 2455 36332 2872 36360
rect 2455 36329 2467 36332
rect 2409 36323 2467 36329
rect 2866 36320 2872 36332
rect 2924 36320 2930 36372
rect 22738 36320 22744 36372
rect 22796 36360 22802 36372
rect 35802 36360 35808 36372
rect 22796 36332 35808 36360
rect 22796 36320 22802 36332
rect 35802 36320 35808 36332
rect 35860 36320 35866 36372
rect 37182 36320 37188 36372
rect 37240 36360 37246 36372
rect 37461 36363 37519 36369
rect 37461 36360 37473 36363
rect 37240 36332 37473 36360
rect 37240 36320 37246 36332
rect 37461 36329 37473 36332
rect 37507 36329 37519 36363
rect 37461 36323 37519 36329
rect 38197 36363 38255 36369
rect 38197 36329 38209 36363
rect 38243 36360 38255 36363
rect 38654 36360 38660 36372
rect 38243 36332 38660 36360
rect 38243 36329 38255 36332
rect 38197 36323 38255 36329
rect 38654 36320 38660 36332
rect 38712 36320 38718 36372
rect 1854 36156 1860 36168
rect 1815 36128 1860 36156
rect 1854 36116 1860 36128
rect 1912 36116 1918 36168
rect 37277 36159 37335 36165
rect 37277 36156 37289 36159
rect 36740 36128 37289 36156
rect 36740 36032 36768 36128
rect 37277 36125 37289 36128
rect 37323 36125 37335 36159
rect 38010 36156 38016 36168
rect 37971 36128 38016 36156
rect 37277 36119 37335 36125
rect 38010 36116 38016 36128
rect 38068 36116 38074 36168
rect 1670 36020 1676 36032
rect 1631 35992 1676 36020
rect 1670 35980 1676 35992
rect 1728 35980 1734 36032
rect 36722 36020 36728 36032
rect 36683 35992 36728 36020
rect 36722 35980 36728 35992
rect 36780 35980 36786 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 1854 35776 1860 35828
rect 1912 35816 1918 35828
rect 2133 35819 2191 35825
rect 2133 35816 2145 35819
rect 1912 35788 2145 35816
rect 1912 35776 1918 35788
rect 2133 35785 2145 35788
rect 2179 35785 2191 35819
rect 2133 35779 2191 35785
rect 2225 35683 2283 35689
rect 2225 35649 2237 35683
rect 2271 35680 2283 35683
rect 2271 35652 2820 35680
rect 2271 35649 2283 35652
rect 2225 35643 2283 35649
rect 2792 35485 2820 35652
rect 37918 35572 37924 35624
rect 37976 35612 37982 35624
rect 38013 35615 38071 35621
rect 38013 35612 38025 35615
rect 37976 35584 38025 35612
rect 37976 35572 37982 35584
rect 38013 35581 38025 35584
rect 38059 35581 38071 35615
rect 38286 35612 38292 35624
rect 38247 35584 38292 35612
rect 38013 35575 38071 35581
rect 38286 35572 38292 35584
rect 38344 35572 38350 35624
rect 2777 35479 2835 35485
rect 2777 35445 2789 35479
rect 2823 35476 2835 35479
rect 3418 35476 3424 35488
rect 2823 35448 3424 35476
rect 2823 35445 2835 35448
rect 2777 35439 2835 35445
rect 3418 35436 3424 35448
rect 3476 35436 3482 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 20257 35275 20315 35281
rect 20257 35241 20269 35275
rect 20303 35272 20315 35275
rect 20714 35272 20720 35284
rect 20303 35244 20720 35272
rect 20303 35241 20315 35244
rect 20257 35235 20315 35241
rect 20714 35232 20720 35244
rect 20772 35232 20778 35284
rect 29917 35275 29975 35281
rect 29917 35241 29929 35275
rect 29963 35272 29975 35275
rect 30466 35272 30472 35284
rect 29963 35244 30472 35272
rect 29963 35241 29975 35244
rect 29917 35235 29975 35241
rect 30466 35232 30472 35244
rect 30524 35232 30530 35284
rect 38286 35272 38292 35284
rect 38247 35244 38292 35272
rect 38286 35232 38292 35244
rect 38344 35232 38350 35284
rect 19978 35028 19984 35080
rect 20036 35068 20042 35080
rect 20073 35071 20131 35077
rect 20073 35068 20085 35071
rect 20036 35040 20085 35068
rect 20036 35028 20042 35040
rect 20073 35037 20085 35040
rect 20119 35068 20131 35071
rect 20717 35071 20775 35077
rect 20717 35068 20729 35071
rect 20119 35040 20729 35068
rect 20119 35037 20131 35040
rect 20073 35031 20131 35037
rect 20717 35037 20729 35040
rect 20763 35037 20775 35071
rect 20717 35031 20775 35037
rect 29638 35028 29644 35080
rect 29696 35068 29702 35080
rect 29733 35071 29791 35077
rect 29733 35068 29745 35071
rect 29696 35040 29745 35068
rect 29696 35028 29702 35040
rect 29733 35037 29745 35040
rect 29779 35068 29791 35071
rect 30377 35071 30435 35077
rect 30377 35068 30389 35071
rect 29779 35040 30389 35068
rect 29779 35037 29791 35040
rect 29733 35031 29791 35037
rect 30377 35037 30389 35040
rect 30423 35037 30435 35071
rect 30377 35031 30435 35037
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1857 34595 1915 34601
rect 1857 34561 1869 34595
rect 1903 34592 1915 34595
rect 1903 34564 2268 34592
rect 1903 34561 1915 34564
rect 1857 34555 1915 34561
rect 2240 34536 2268 34564
rect 2222 34484 2228 34536
rect 2280 34524 2286 34536
rect 2317 34527 2375 34533
rect 2317 34524 2329 34527
rect 2280 34496 2329 34524
rect 2280 34484 2286 34496
rect 2317 34493 2329 34496
rect 2363 34493 2375 34527
rect 2317 34487 2375 34493
rect 1670 34388 1676 34400
rect 1631 34360 1676 34388
rect 1670 34348 1676 34360
rect 1728 34348 1734 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 6730 34144 6736 34196
rect 6788 34184 6794 34196
rect 7009 34187 7067 34193
rect 7009 34184 7021 34187
rect 6788 34156 7021 34184
rect 6788 34144 6794 34156
rect 7009 34153 7021 34156
rect 7055 34153 7067 34187
rect 7009 34147 7067 34153
rect 7098 33980 7104 33992
rect 7059 33952 7104 33980
rect 7098 33940 7104 33952
rect 7156 33980 7162 33992
rect 7561 33983 7619 33989
rect 7561 33980 7573 33983
rect 7156 33952 7573 33980
rect 7156 33940 7162 33952
rect 7561 33949 7573 33952
rect 7607 33949 7619 33983
rect 7561 33943 7619 33949
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 12710 33464 12716 33516
rect 12768 33504 12774 33516
rect 37461 33507 37519 33513
rect 37461 33504 37473 33507
rect 12768 33476 37473 33504
rect 12768 33464 12774 33476
rect 37461 33473 37473 33476
rect 37507 33504 37519 33507
rect 38013 33507 38071 33513
rect 38013 33504 38025 33507
rect 37507 33476 38025 33504
rect 37507 33473 37519 33476
rect 37461 33467 37519 33473
rect 38013 33473 38025 33476
rect 38059 33473 38071 33507
rect 38013 33467 38071 33473
rect 38194 33368 38200 33380
rect 38155 33340 38200 33368
rect 38194 33328 38200 33340
rect 38252 33328 38258 33380
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 1578 32376 1584 32428
rect 1636 32416 1642 32428
rect 1673 32419 1731 32425
rect 1673 32416 1685 32419
rect 1636 32388 1685 32416
rect 1636 32376 1642 32388
rect 1673 32385 1685 32388
rect 1719 32385 1731 32419
rect 19978 32416 19984 32428
rect 1673 32379 1731 32385
rect 16546 32388 19984 32416
rect 1765 32215 1823 32221
rect 1765 32181 1777 32215
rect 1811 32212 1823 32215
rect 12986 32212 12992 32224
rect 1811 32184 12992 32212
rect 1811 32181 1823 32184
rect 1765 32175 1823 32181
rect 12986 32172 12992 32184
rect 13044 32212 13050 32224
rect 16546 32212 16574 32388
rect 19978 32376 19984 32388
rect 20036 32376 20042 32428
rect 29638 32376 29644 32428
rect 29696 32416 29702 32428
rect 38013 32419 38071 32425
rect 38013 32416 38025 32419
rect 29696 32388 38025 32416
rect 29696 32376 29702 32388
rect 38013 32385 38025 32388
rect 38059 32385 38071 32419
rect 38013 32379 38071 32385
rect 38286 32348 38292 32360
rect 38247 32320 38292 32348
rect 38286 32308 38292 32320
rect 38344 32308 38350 32360
rect 13044 32184 16574 32212
rect 13044 32172 13050 32184
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 1578 32008 1584 32020
rect 1539 31980 1584 32008
rect 1578 31968 1584 31980
rect 1636 31968 1642 32020
rect 38286 32008 38292 32020
rect 38247 31980 38292 32008
rect 38286 31968 38292 31980
rect 38344 31968 38350 32020
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 27430 30920 27436 30932
rect 27391 30892 27436 30920
rect 27430 30880 27436 30892
rect 27488 30880 27494 30932
rect 30834 30920 30840 30932
rect 30795 30892 30840 30920
rect 30834 30880 30840 30892
rect 30892 30880 30898 30932
rect 27249 30719 27307 30725
rect 27249 30685 27261 30719
rect 27295 30716 27307 30719
rect 27295 30688 28028 30716
rect 27295 30685 27307 30688
rect 27249 30679 27307 30685
rect 1670 30648 1676 30660
rect 1631 30620 1676 30648
rect 1670 30608 1676 30620
rect 1728 30608 1734 30660
rect 1762 30580 1768 30592
rect 1723 30552 1768 30580
rect 1762 30540 1768 30552
rect 1820 30540 1826 30592
rect 28000 30589 28028 30688
rect 30558 30676 30564 30728
rect 30616 30716 30622 30728
rect 30745 30719 30803 30725
rect 30745 30716 30757 30719
rect 30616 30688 30757 30716
rect 30616 30676 30622 30688
rect 30745 30685 30757 30688
rect 30791 30716 30803 30719
rect 31389 30719 31447 30725
rect 31389 30716 31401 30719
rect 30791 30688 31401 30716
rect 30791 30685 30803 30688
rect 30745 30679 30803 30685
rect 31389 30685 31401 30688
rect 31435 30685 31447 30719
rect 31389 30679 31447 30685
rect 27985 30583 28043 30589
rect 27985 30549 27997 30583
rect 28031 30580 28043 30583
rect 29270 30580 29276 30592
rect 28031 30552 29276 30580
rect 28031 30549 28043 30552
rect 27985 30543 28043 30549
rect 29270 30540 29276 30552
rect 29328 30540 29334 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 1670 30376 1676 30388
rect 1631 30348 1676 30376
rect 1670 30336 1676 30348
rect 1728 30336 1734 30388
rect 14734 30200 14740 30252
rect 14792 30240 14798 30252
rect 15381 30243 15439 30249
rect 15381 30240 15393 30243
rect 14792 30212 15393 30240
rect 14792 30200 14798 30212
rect 15381 30209 15393 30212
rect 15427 30209 15439 30243
rect 38010 30240 38016 30252
rect 37971 30212 38016 30240
rect 15381 30203 15439 30209
rect 38010 30200 38016 30212
rect 38068 30200 38074 30252
rect 14734 30036 14740 30048
rect 14695 30008 14740 30036
rect 14734 29996 14740 30008
rect 14792 29996 14798 30048
rect 15473 30039 15531 30045
rect 15473 30005 15485 30039
rect 15519 30036 15531 30039
rect 36722 30036 36728 30048
rect 15519 30008 36728 30036
rect 15519 30005 15531 30008
rect 15473 29999 15531 30005
rect 36722 29996 36728 30008
rect 36780 29996 36786 30048
rect 38194 30036 38200 30048
rect 38155 30008 38200 30036
rect 38194 29996 38200 30008
rect 38252 29996 38258 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 38010 29832 38016 29844
rect 37971 29804 38016 29832
rect 38010 29792 38016 29804
rect 38068 29792 38074 29844
rect 37826 29628 37832 29640
rect 37787 29600 37832 29628
rect 37826 29588 37832 29600
rect 37884 29588 37890 29640
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 37826 29248 37832 29300
rect 37884 29288 37890 29300
rect 38102 29288 38108 29300
rect 37884 29260 38108 29288
rect 37884 29248 37890 29260
rect 38102 29248 38108 29260
rect 38160 29248 38166 29300
rect 20530 29152 20536 29164
rect 20491 29124 20536 29152
rect 20530 29112 20536 29124
rect 20588 29112 20594 29164
rect 1578 29084 1584 29096
rect 1539 29056 1584 29084
rect 1578 29044 1584 29056
rect 1636 29044 1642 29096
rect 1857 29087 1915 29093
rect 1857 29053 1869 29087
rect 1903 29084 1915 29087
rect 14734 29084 14740 29096
rect 1903 29056 14740 29084
rect 1903 29053 1915 29056
rect 1857 29047 1915 29053
rect 14734 29044 14740 29056
rect 14792 29044 14798 29096
rect 20254 28976 20260 29028
rect 20312 29016 20318 29028
rect 20441 29019 20499 29025
rect 20441 29016 20453 29019
rect 20312 28988 20453 29016
rect 20312 28976 20318 28988
rect 20441 28985 20453 28988
rect 20487 28985 20499 29019
rect 20441 28979 20499 28985
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 22278 28744 22284 28756
rect 22239 28716 22284 28744
rect 22278 28704 22284 28716
rect 22336 28704 22342 28756
rect 1578 28676 1584 28688
rect 1539 28648 1584 28676
rect 1578 28636 1584 28648
rect 1636 28636 1642 28688
rect 13265 28543 13323 28549
rect 13265 28509 13277 28543
rect 13311 28540 13323 28543
rect 13354 28540 13360 28552
rect 13311 28512 13360 28540
rect 13311 28509 13323 28512
rect 13265 28503 13323 28509
rect 13354 28500 13360 28512
rect 13412 28500 13418 28552
rect 21821 28543 21879 28549
rect 21821 28509 21833 28543
rect 21867 28540 21879 28543
rect 22278 28540 22284 28552
rect 21867 28512 22284 28540
rect 21867 28509 21879 28512
rect 21821 28503 21879 28509
rect 22278 28500 22284 28512
rect 22336 28500 22342 28552
rect 13357 28407 13415 28413
rect 13357 28373 13369 28407
rect 13403 28404 13415 28407
rect 14274 28404 14280 28416
rect 13403 28376 14280 28404
rect 13403 28373 13415 28376
rect 13357 28367 13415 28373
rect 14274 28364 14280 28376
rect 14332 28364 14338 28416
rect 21729 28407 21787 28413
rect 21729 28373 21741 28407
rect 21775 28404 21787 28407
rect 22646 28404 22652 28416
rect 21775 28376 22652 28404
rect 21775 28373 21787 28376
rect 21729 28367 21787 28373
rect 22646 28364 22652 28376
rect 22704 28364 22710 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 13170 28160 13176 28212
rect 13228 28200 13234 28212
rect 14461 28203 14519 28209
rect 14461 28200 14473 28203
rect 13228 28172 14473 28200
rect 13228 28160 13234 28172
rect 14461 28169 14473 28172
rect 14507 28169 14519 28203
rect 14461 28163 14519 28169
rect 14553 28067 14611 28073
rect 14553 28033 14565 28067
rect 14599 28064 14611 28067
rect 14599 28036 15148 28064
rect 14599 28033 14611 28036
rect 14553 28027 14611 28033
rect 15120 27869 15148 28036
rect 16482 28024 16488 28076
rect 16540 28064 16546 28076
rect 37461 28067 37519 28073
rect 37461 28064 37473 28067
rect 16540 28036 37473 28064
rect 16540 28024 16546 28036
rect 37461 28033 37473 28036
rect 37507 28064 37519 28067
rect 38013 28067 38071 28073
rect 38013 28064 38025 28067
rect 37507 28036 38025 28064
rect 37507 28033 37519 28036
rect 37461 28027 37519 28033
rect 38013 28033 38025 28036
rect 38059 28033 38071 28067
rect 38013 28027 38071 28033
rect 38194 27928 38200 27940
rect 38155 27900 38200 27928
rect 38194 27888 38200 27900
rect 38252 27888 38258 27940
rect 15105 27863 15163 27869
rect 15105 27829 15117 27863
rect 15151 27860 15163 27863
rect 17586 27860 17592 27872
rect 15151 27832 17592 27860
rect 15151 27829 15163 27832
rect 15105 27823 15163 27829
rect 17586 27820 17592 27832
rect 17644 27820 17650 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 22094 27044 22100 27056
rect 22055 27016 22100 27044
rect 22094 27004 22100 27016
rect 22152 27004 22158 27056
rect 1857 26979 1915 26985
rect 1857 26945 1869 26979
rect 1903 26976 1915 26979
rect 6546 26976 6552 26988
rect 1903 26948 6552 26976
rect 1903 26945 1915 26948
rect 1857 26939 1915 26945
rect 6546 26936 6552 26948
rect 6604 26936 6610 26988
rect 22281 26979 22339 26985
rect 22281 26945 22293 26979
rect 22327 26976 22339 26979
rect 30653 26979 30711 26985
rect 22327 26948 22968 26976
rect 22327 26945 22339 26948
rect 22281 26939 22339 26945
rect 1670 26772 1676 26784
rect 1631 26744 1676 26772
rect 1670 26732 1676 26744
rect 1728 26732 1734 26784
rect 22940 26781 22968 26948
rect 30653 26945 30665 26979
rect 30699 26976 30711 26979
rect 37918 26976 37924 26988
rect 30699 26948 37924 26976
rect 30699 26945 30711 26948
rect 30653 26939 30711 26945
rect 37918 26936 37924 26948
rect 37976 26936 37982 26988
rect 38010 26908 38016 26920
rect 37971 26880 38016 26908
rect 38010 26868 38016 26880
rect 38068 26868 38074 26920
rect 38286 26908 38292 26920
rect 38247 26880 38292 26908
rect 38286 26868 38292 26880
rect 38344 26868 38350 26920
rect 22925 26775 22983 26781
rect 22925 26741 22937 26775
rect 22971 26772 22983 26775
rect 23382 26772 23388 26784
rect 22971 26744 23388 26772
rect 22971 26741 22983 26744
rect 22925 26735 22983 26741
rect 23382 26732 23388 26744
rect 23440 26732 23446 26784
rect 26418 26732 26424 26784
rect 26476 26772 26482 26784
rect 30561 26775 30619 26781
rect 30561 26772 30573 26775
rect 26476 26744 30573 26772
rect 26476 26732 26482 26744
rect 30561 26741 30573 26744
rect 30607 26741 30619 26775
rect 30561 26735 30619 26741
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 23382 26528 23388 26580
rect 23440 26568 23446 26580
rect 38010 26568 38016 26580
rect 23440 26540 38016 26568
rect 23440 26528 23446 26540
rect 38010 26528 38016 26540
rect 38068 26528 38074 26580
rect 38286 26568 38292 26580
rect 38247 26540 38292 26568
rect 38286 26528 38292 26540
rect 38344 26528 38350 26580
rect 16482 26500 16488 26512
rect 16443 26472 16488 26500
rect 16482 26460 16488 26472
rect 16540 26460 16546 26512
rect 15749 26367 15807 26373
rect 15749 26333 15761 26367
rect 15795 26364 15807 26367
rect 16298 26364 16304 26376
rect 15795 26336 16304 26364
rect 15795 26333 15807 26336
rect 15749 26327 15807 26333
rect 16298 26324 16304 26336
rect 16356 26324 16362 26376
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 13262 25984 13268 26036
rect 13320 26024 13326 26036
rect 18877 26027 18935 26033
rect 18877 26024 18889 26027
rect 13320 25996 18889 26024
rect 13320 25984 13326 25996
rect 18877 25993 18889 25996
rect 18923 25993 18935 26027
rect 18877 25987 18935 25993
rect 18230 25848 18236 25900
rect 18288 25888 18294 25900
rect 19061 25891 19119 25897
rect 19061 25888 19073 25891
rect 18288 25860 19073 25888
rect 18288 25848 18294 25860
rect 19061 25857 19073 25860
rect 19107 25888 19119 25891
rect 19521 25891 19579 25897
rect 19521 25888 19533 25891
rect 19107 25860 19533 25888
rect 19107 25857 19119 25860
rect 19061 25851 19119 25857
rect 19521 25857 19533 25860
rect 19567 25857 19579 25891
rect 19521 25851 19579 25857
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 12986 25480 12992 25492
rect 12947 25452 12992 25480
rect 12986 25440 12992 25452
rect 13044 25440 13050 25492
rect 28445 25483 28503 25489
rect 28445 25449 28457 25483
rect 28491 25480 28503 25483
rect 29638 25480 29644 25492
rect 28491 25452 29644 25480
rect 28491 25449 28503 25452
rect 28445 25443 28503 25449
rect 1578 25276 1584 25288
rect 1539 25248 1584 25276
rect 1578 25236 1584 25248
rect 1636 25236 1642 25288
rect 1857 25279 1915 25285
rect 1857 25245 1869 25279
rect 1903 25276 1915 25279
rect 2038 25276 2044 25288
rect 1903 25248 2044 25276
rect 1903 25245 1915 25248
rect 1857 25239 1915 25245
rect 2038 25236 2044 25248
rect 2096 25236 2102 25288
rect 12986 25236 12992 25288
rect 13044 25276 13050 25288
rect 13725 25279 13783 25285
rect 13725 25276 13737 25279
rect 13044 25248 13737 25276
rect 13044 25236 13050 25248
rect 13725 25245 13737 25248
rect 13771 25245 13783 25279
rect 13725 25239 13783 25245
rect 16117 25279 16175 25285
rect 16117 25245 16129 25279
rect 16163 25276 16175 25279
rect 16298 25276 16304 25288
rect 16163 25248 16304 25276
rect 16163 25245 16175 25248
rect 16117 25239 16175 25245
rect 16298 25236 16304 25248
rect 16356 25276 16362 25288
rect 16761 25279 16819 25285
rect 16761 25276 16773 25279
rect 16356 25248 16773 25276
rect 16356 25236 16362 25248
rect 16761 25245 16773 25248
rect 16807 25245 16819 25279
rect 16761 25239 16819 25245
rect 27893 25279 27951 25285
rect 27893 25245 27905 25279
rect 27939 25276 27951 25279
rect 28460 25276 28488 25443
rect 29638 25440 29644 25452
rect 29696 25440 29702 25492
rect 27939 25248 28488 25276
rect 27939 25245 27951 25248
rect 27893 25239 27951 25245
rect 16209 25211 16267 25217
rect 16209 25177 16221 25211
rect 16255 25208 16267 25211
rect 16942 25208 16948 25220
rect 16255 25180 16948 25208
rect 16255 25177 16267 25180
rect 16209 25171 16267 25177
rect 16942 25168 16948 25180
rect 17000 25168 17006 25220
rect 12894 25100 12900 25152
rect 12952 25140 12958 25152
rect 13633 25143 13691 25149
rect 13633 25140 13645 25143
rect 12952 25112 13645 25140
rect 12952 25100 12958 25112
rect 13633 25109 13645 25112
rect 13679 25109 13691 25143
rect 13633 25103 13691 25109
rect 25222 25100 25228 25152
rect 25280 25140 25286 25152
rect 27801 25143 27859 25149
rect 27801 25140 27813 25143
rect 25280 25112 27813 25140
rect 25280 25100 25286 25112
rect 27801 25109 27813 25112
rect 27847 25109 27859 25143
rect 27801 25103 27859 25109
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 1578 24936 1584 24948
rect 1539 24908 1584 24936
rect 1578 24896 1584 24908
rect 1636 24896 1642 24948
rect 37553 24803 37611 24809
rect 37553 24769 37565 24803
rect 37599 24800 37611 24803
rect 38010 24800 38016 24812
rect 37599 24772 38016 24800
rect 37599 24769 37611 24772
rect 37553 24763 37611 24769
rect 38010 24760 38016 24772
rect 38068 24760 38074 24812
rect 38194 24596 38200 24608
rect 38155 24568 38200 24596
rect 38194 24556 38200 24568
rect 38252 24556 38258 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 31297 24395 31355 24401
rect 31297 24361 31309 24395
rect 31343 24392 31355 24395
rect 38102 24392 38108 24404
rect 31343 24364 38108 24392
rect 31343 24361 31355 24364
rect 31297 24355 31355 24361
rect 30745 24191 30803 24197
rect 30745 24157 30757 24191
rect 30791 24188 30803 24191
rect 31312 24188 31340 24355
rect 38102 24352 38108 24364
rect 38160 24352 38166 24404
rect 30791 24160 31340 24188
rect 30791 24157 30803 24160
rect 30745 24151 30803 24157
rect 7098 24080 7104 24132
rect 7156 24120 7162 24132
rect 17770 24120 17776 24132
rect 7156 24092 17776 24120
rect 7156 24080 7162 24092
rect 17770 24080 17776 24092
rect 17828 24080 17834 24132
rect 24118 24080 24124 24132
rect 24176 24120 24182 24132
rect 30558 24120 30564 24132
rect 24176 24092 30564 24120
rect 24176 24080 24182 24092
rect 30558 24080 30564 24092
rect 30616 24080 30622 24132
rect 24854 24012 24860 24064
rect 24912 24052 24918 24064
rect 30653 24055 30711 24061
rect 30653 24052 30665 24055
rect 24912 24024 30665 24052
rect 24912 24012 24918 24024
rect 30653 24021 30665 24024
rect 30699 24021 30711 24055
rect 30653 24015 30711 24021
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 1854 23712 1860 23724
rect 1815 23684 1860 23712
rect 1854 23672 1860 23684
rect 1912 23672 1918 23724
rect 1670 23508 1676 23520
rect 1631 23480 1676 23508
rect 1670 23468 1676 23480
rect 1728 23468 1734 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 14826 22624 14832 22636
rect 14787 22596 14832 22624
rect 14826 22584 14832 22596
rect 14884 22624 14890 22636
rect 15289 22627 15347 22633
rect 15289 22624 15301 22627
rect 14884 22596 15301 22624
rect 14884 22584 14890 22596
rect 15289 22593 15301 22596
rect 15335 22593 15347 22627
rect 15289 22587 15347 22593
rect 37553 22627 37611 22633
rect 37553 22593 37565 22627
rect 37599 22624 37611 22627
rect 38194 22624 38200 22636
rect 37599 22596 38200 22624
rect 37599 22593 37611 22596
rect 37553 22587 37611 22593
rect 38194 22584 38200 22596
rect 38252 22584 38258 22636
rect 37918 22448 37924 22500
rect 37976 22488 37982 22500
rect 38013 22491 38071 22497
rect 38013 22488 38025 22491
rect 37976 22460 38025 22488
rect 37976 22448 37982 22460
rect 38013 22457 38025 22460
rect 38059 22457 38071 22491
rect 38013 22451 38071 22457
rect 14366 22380 14372 22432
rect 14424 22420 14430 22432
rect 14737 22423 14795 22429
rect 14737 22420 14749 22423
rect 14424 22392 14749 22420
rect 14424 22380 14430 22392
rect 14737 22389 14749 22392
rect 14783 22389 14795 22423
rect 14737 22383 14795 22389
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 6546 21672 6552 21684
rect 6507 21644 6552 21672
rect 6546 21632 6552 21644
rect 6604 21632 6610 21684
rect 19978 21672 19984 21684
rect 19939 21644 19984 21672
rect 19978 21632 19984 21644
rect 20036 21632 20042 21684
rect 25866 21672 25872 21684
rect 25827 21644 25872 21672
rect 25866 21632 25872 21644
rect 25924 21632 25930 21684
rect 1762 21496 1768 21548
rect 1820 21536 1826 21548
rect 1857 21539 1915 21545
rect 1857 21536 1869 21539
rect 1820 21508 1869 21536
rect 1820 21496 1826 21508
rect 1857 21505 1869 21508
rect 1903 21505 1915 21539
rect 1857 21499 1915 21505
rect 6733 21539 6791 21545
rect 6733 21505 6745 21539
rect 6779 21536 6791 21539
rect 6779 21508 7328 21536
rect 6779 21505 6791 21508
rect 6733 21499 6791 21505
rect 1670 21332 1676 21344
rect 1631 21304 1676 21332
rect 1670 21292 1676 21304
rect 1728 21292 1734 21344
rect 7300 21341 7328 21508
rect 17770 21496 17776 21548
rect 17828 21536 17834 21548
rect 19797 21539 19855 21545
rect 19797 21536 19809 21539
rect 17828 21508 19809 21536
rect 17828 21496 17834 21508
rect 19797 21505 19809 21508
rect 19843 21536 19855 21539
rect 20441 21539 20499 21545
rect 20441 21536 20453 21539
rect 19843 21508 20453 21536
rect 19843 21505 19855 21508
rect 19797 21499 19855 21505
rect 20441 21505 20453 21508
rect 20487 21505 20499 21539
rect 20441 21499 20499 21505
rect 25685 21539 25743 21545
rect 25685 21505 25697 21539
rect 25731 21536 25743 21539
rect 26329 21539 26387 21545
rect 26329 21536 26341 21539
rect 25731 21508 26341 21536
rect 25731 21505 25743 21508
rect 25685 21499 25743 21505
rect 26329 21505 26341 21508
rect 26375 21536 26387 21539
rect 28626 21536 28632 21548
rect 26375 21508 28632 21536
rect 26375 21505 26387 21508
rect 26329 21499 26387 21505
rect 28626 21496 28632 21508
rect 28684 21496 28690 21548
rect 37458 21496 37464 21548
rect 37516 21536 37522 21548
rect 38013 21539 38071 21545
rect 38013 21536 38025 21539
rect 37516 21508 38025 21536
rect 37516 21496 37522 21508
rect 38013 21505 38025 21508
rect 38059 21505 38071 21539
rect 38013 21499 38071 21505
rect 7285 21335 7343 21341
rect 7285 21301 7297 21335
rect 7331 21332 7343 21335
rect 10042 21332 10048 21344
rect 7331 21304 10048 21332
rect 7331 21301 7343 21304
rect 7285 21295 7343 21301
rect 10042 21292 10048 21304
rect 10100 21292 10106 21344
rect 37458 21332 37464 21344
rect 37419 21304 37464 21332
rect 37458 21292 37464 21304
rect 37516 21292 37522 21344
rect 38194 21332 38200 21344
rect 38155 21304 38200 21332
rect 38194 21292 38200 21304
rect 38252 21292 38258 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 1762 21128 1768 21140
rect 1723 21100 1768 21128
rect 1762 21088 1768 21100
rect 1820 21088 1826 21140
rect 1949 20927 2007 20933
rect 1949 20893 1961 20927
rect 1995 20924 2007 20927
rect 2038 20924 2044 20936
rect 1995 20896 2044 20924
rect 1995 20893 2007 20896
rect 1949 20887 2007 20893
rect 2038 20884 2044 20896
rect 2096 20884 2102 20936
rect 19426 20788 19432 20800
rect 19387 20760 19432 20788
rect 19426 20748 19432 20760
rect 19484 20748 19490 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 19334 20516 19340 20528
rect 19295 20488 19340 20516
rect 19334 20476 19340 20488
rect 19392 20476 19398 20528
rect 19426 20476 19432 20528
rect 19484 20516 19490 20528
rect 19484 20488 19529 20516
rect 19484 20476 19490 20488
rect 19150 20380 19156 20392
rect 19111 20352 19156 20380
rect 19150 20340 19156 20352
rect 19208 20340 19214 20392
rect 19610 20204 19616 20256
rect 19668 20244 19674 20256
rect 19981 20247 20039 20253
rect 19981 20244 19993 20247
rect 19668 20216 19993 20244
rect 19668 20204 19674 20216
rect 19981 20213 19993 20216
rect 20027 20213 20039 20247
rect 19981 20207 20039 20213
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 2314 20040 2320 20052
rect 2275 20012 2320 20040
rect 2314 20000 2320 20012
rect 2372 20000 2378 20052
rect 19334 20000 19340 20052
rect 19392 20040 19398 20052
rect 19521 20043 19579 20049
rect 19521 20040 19533 20043
rect 19392 20012 19533 20040
rect 19392 20000 19398 20012
rect 19521 20009 19533 20012
rect 19567 20009 19579 20043
rect 19521 20003 19579 20009
rect 23382 20000 23388 20052
rect 23440 20040 23446 20052
rect 23661 20043 23719 20049
rect 23661 20040 23673 20043
rect 23440 20012 23673 20040
rect 23440 20000 23446 20012
rect 23661 20009 23673 20012
rect 23707 20009 23719 20043
rect 23661 20003 23719 20009
rect 1946 19864 1952 19916
rect 2004 19904 2010 19916
rect 2004 19876 20300 19904
rect 2004 19864 2010 19876
rect 1857 19839 1915 19845
rect 1857 19805 1869 19839
rect 1903 19805 1915 19839
rect 1857 19799 1915 19805
rect 2501 19839 2559 19845
rect 2501 19805 2513 19839
rect 2547 19836 2559 19839
rect 2590 19836 2596 19848
rect 2547 19808 2596 19836
rect 2547 19805 2559 19808
rect 2501 19799 2559 19805
rect 1872 19768 1900 19799
rect 2590 19796 2596 19808
rect 2648 19836 2654 19848
rect 2961 19839 3019 19845
rect 2961 19836 2973 19839
rect 2648 19808 2973 19836
rect 2648 19796 2654 19808
rect 2961 19805 2973 19808
rect 3007 19805 3019 19839
rect 18693 19839 18751 19845
rect 18693 19836 18705 19839
rect 2961 19799 3019 19805
rect 18156 19808 18705 19836
rect 4614 19768 4620 19780
rect 1872 19740 4620 19768
rect 4614 19728 4620 19740
rect 4672 19728 4678 19780
rect 1670 19700 1676 19712
rect 1631 19672 1676 19700
rect 1670 19660 1676 19672
rect 1728 19660 1734 19712
rect 16114 19660 16120 19712
rect 16172 19700 16178 19712
rect 18156 19709 18184 19808
rect 18693 19805 18705 19808
rect 18739 19836 18751 19839
rect 19610 19836 19616 19848
rect 18739 19808 19616 19836
rect 18739 19805 18751 19808
rect 18693 19799 18751 19805
rect 19610 19796 19616 19808
rect 19668 19796 19674 19848
rect 20272 19845 20300 19876
rect 20257 19839 20315 19845
rect 20257 19805 20269 19839
rect 20303 19836 20315 19839
rect 20717 19839 20775 19845
rect 20717 19836 20729 19839
rect 20303 19808 20729 19836
rect 20303 19805 20315 19808
rect 20257 19799 20315 19805
rect 20717 19805 20729 19808
rect 20763 19836 20775 19839
rect 22094 19836 22100 19848
rect 20763 19808 22100 19836
rect 20763 19805 20775 19808
rect 20717 19799 20775 19805
rect 22094 19796 22100 19808
rect 22152 19796 22158 19848
rect 23201 19839 23259 19845
rect 23201 19805 23213 19839
rect 23247 19836 23259 19839
rect 23382 19836 23388 19848
rect 23247 19808 23388 19836
rect 23247 19805 23259 19808
rect 23201 19799 23259 19805
rect 23382 19796 23388 19808
rect 23440 19796 23446 19848
rect 19978 19728 19984 19780
rect 20036 19768 20042 19780
rect 20165 19771 20223 19777
rect 20165 19768 20177 19771
rect 20036 19740 20177 19768
rect 20036 19728 20042 19740
rect 20165 19737 20177 19740
rect 20211 19737 20223 19771
rect 20165 19731 20223 19737
rect 18141 19703 18199 19709
rect 18141 19700 18153 19703
rect 16172 19672 18153 19700
rect 16172 19660 16178 19672
rect 18141 19669 18153 19672
rect 18187 19669 18199 19703
rect 18141 19663 18199 19669
rect 18785 19703 18843 19709
rect 18785 19669 18797 19703
rect 18831 19700 18843 19703
rect 20070 19700 20076 19712
rect 18831 19672 20076 19700
rect 18831 19669 18843 19672
rect 18785 19663 18843 19669
rect 20070 19660 20076 19672
rect 20128 19660 20134 19712
rect 23106 19700 23112 19712
rect 23067 19672 23112 19700
rect 23106 19660 23112 19672
rect 23164 19660 23170 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 1854 19456 1860 19508
rect 1912 19496 1918 19508
rect 1949 19499 2007 19505
rect 1949 19496 1961 19499
rect 1912 19468 1961 19496
rect 1912 19456 1918 19468
rect 1949 19465 1961 19468
rect 1995 19465 2007 19499
rect 1949 19459 2007 19465
rect 2498 19456 2504 19508
rect 2556 19496 2562 19508
rect 2556 19468 12204 19496
rect 2556 19456 2562 19468
rect 2038 19388 2044 19440
rect 2096 19428 2102 19440
rect 12176 19428 12204 19468
rect 12250 19456 12256 19508
rect 12308 19496 12314 19508
rect 15470 19496 15476 19508
rect 12308 19468 15476 19496
rect 12308 19456 12314 19468
rect 15470 19456 15476 19468
rect 15528 19456 15534 19508
rect 2096 19400 9720 19428
rect 12176 19400 20484 19428
rect 2096 19388 2102 19400
rect 2130 19360 2136 19372
rect 2043 19332 2136 19360
rect 2130 19320 2136 19332
rect 2188 19360 2194 19372
rect 9692 19369 9720 19400
rect 9677 19363 9735 19369
rect 2188 19332 2728 19360
rect 2188 19320 2194 19332
rect 2700 19165 2728 19332
rect 9677 19329 9689 19363
rect 9723 19329 9735 19363
rect 9677 19323 9735 19329
rect 9769 19363 9827 19369
rect 9769 19329 9781 19363
rect 9815 19360 9827 19363
rect 12250 19360 12256 19372
rect 9815 19332 12256 19360
rect 9815 19329 9827 19332
rect 9769 19323 9827 19329
rect 12250 19320 12256 19332
rect 12308 19320 12314 19372
rect 12621 19363 12679 19369
rect 12621 19360 12633 19363
rect 12406 19332 12633 19360
rect 2685 19159 2743 19165
rect 2685 19125 2697 19159
rect 2731 19156 2743 19159
rect 9674 19156 9680 19168
rect 2731 19128 9680 19156
rect 2731 19125 2743 19128
rect 2685 19119 2743 19125
rect 9674 19116 9680 19128
rect 9732 19116 9738 19168
rect 11514 19116 11520 19168
rect 11572 19156 11578 19168
rect 11977 19159 12035 19165
rect 11977 19156 11989 19159
rect 11572 19128 11989 19156
rect 11572 19116 11578 19128
rect 11977 19125 11989 19128
rect 12023 19156 12035 19159
rect 12406 19156 12434 19332
rect 12621 19329 12633 19332
rect 12667 19329 12679 19363
rect 12621 19323 12679 19329
rect 19613 19363 19671 19369
rect 19613 19329 19625 19363
rect 19659 19329 19671 19363
rect 20346 19360 20352 19372
rect 20307 19332 20352 19360
rect 19613 19323 19671 19329
rect 12710 19252 12716 19304
rect 12768 19292 12774 19304
rect 12805 19295 12863 19301
rect 12805 19292 12817 19295
rect 12768 19264 12817 19292
rect 12768 19252 12774 19264
rect 12805 19261 12817 19264
rect 12851 19261 12863 19295
rect 12805 19255 12863 19261
rect 19153 19227 19211 19233
rect 19153 19193 19165 19227
rect 19199 19224 19211 19227
rect 19628 19224 19656 19323
rect 20346 19320 20352 19332
rect 20404 19320 20410 19372
rect 20456 19369 20484 19400
rect 20441 19363 20499 19369
rect 20441 19329 20453 19363
rect 20487 19360 20499 19363
rect 20487 19332 20944 19360
rect 20487 19329 20499 19332
rect 20441 19323 20499 19329
rect 20916 19301 20944 19332
rect 36630 19320 36636 19372
rect 36688 19360 36694 19372
rect 38013 19363 38071 19369
rect 38013 19360 38025 19363
rect 36688 19332 38025 19360
rect 36688 19320 36694 19332
rect 38013 19329 38025 19332
rect 38059 19329 38071 19363
rect 38013 19323 38071 19329
rect 20901 19295 20959 19301
rect 20901 19261 20913 19295
rect 20947 19292 20959 19295
rect 24486 19292 24492 19304
rect 20947 19264 24492 19292
rect 20947 19261 20959 19264
rect 20901 19255 20959 19261
rect 24486 19252 24492 19264
rect 24544 19252 24550 19304
rect 19886 19224 19892 19236
rect 19199 19196 19892 19224
rect 19199 19193 19211 19196
rect 19153 19187 19211 19193
rect 19886 19184 19892 19196
rect 19944 19184 19950 19236
rect 21082 19184 21088 19236
rect 21140 19224 21146 19236
rect 22097 19227 22155 19233
rect 22097 19224 22109 19227
rect 21140 19196 22109 19224
rect 21140 19184 21146 19196
rect 22097 19193 22109 19196
rect 22143 19224 22155 19227
rect 24394 19224 24400 19236
rect 22143 19196 24400 19224
rect 22143 19193 22155 19196
rect 22097 19187 22155 19193
rect 24394 19184 24400 19196
rect 24452 19184 24458 19236
rect 12023 19128 12434 19156
rect 19705 19159 19763 19165
rect 12023 19125 12035 19128
rect 11977 19119 12035 19125
rect 19705 19125 19717 19159
rect 19751 19156 19763 19159
rect 20162 19156 20168 19168
rect 19751 19128 20168 19156
rect 19751 19125 19763 19128
rect 19705 19119 19763 19125
rect 20162 19116 20168 19128
rect 20220 19116 20226 19168
rect 23014 19156 23020 19168
rect 22975 19128 23020 19156
rect 23014 19116 23020 19128
rect 23072 19116 23078 19168
rect 23661 19159 23719 19165
rect 23661 19125 23673 19159
rect 23707 19156 23719 19159
rect 23750 19156 23756 19168
rect 23707 19128 23756 19156
rect 23707 19125 23719 19128
rect 23661 19119 23719 19125
rect 23750 19116 23756 19128
rect 23808 19116 23814 19168
rect 38194 19156 38200 19168
rect 38155 19128 38200 19156
rect 38194 19116 38200 19128
rect 38252 19116 38258 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 18230 18952 18236 18964
rect 18191 18924 18236 18952
rect 18230 18912 18236 18924
rect 18288 18952 18294 18964
rect 18506 18952 18512 18964
rect 18288 18924 18512 18952
rect 18288 18912 18294 18924
rect 18506 18912 18512 18924
rect 18564 18912 18570 18964
rect 17126 18844 17132 18896
rect 17184 18884 17190 18896
rect 26878 18884 26884 18896
rect 17184 18856 26884 18884
rect 17184 18844 17190 18856
rect 26878 18844 26884 18856
rect 26936 18844 26942 18896
rect 1762 18776 1768 18828
rect 1820 18816 1826 18828
rect 19426 18816 19432 18828
rect 1820 18788 19432 18816
rect 1820 18776 1826 18788
rect 19426 18776 19432 18788
rect 19484 18776 19490 18828
rect 20165 18819 20223 18825
rect 20165 18785 20177 18819
rect 20211 18816 20223 18819
rect 20438 18816 20444 18828
rect 20211 18788 20444 18816
rect 20211 18785 20223 18788
rect 20165 18779 20223 18785
rect 20438 18776 20444 18788
rect 20496 18776 20502 18828
rect 16853 18751 16911 18757
rect 16853 18717 16865 18751
rect 16899 18748 16911 18751
rect 18230 18748 18236 18760
rect 16899 18720 18236 18748
rect 16899 18717 16911 18720
rect 16853 18711 16911 18717
rect 18230 18708 18236 18720
rect 18288 18708 18294 18760
rect 22094 18708 22100 18760
rect 22152 18748 22158 18760
rect 22741 18751 22799 18757
rect 22741 18748 22753 18751
rect 22152 18720 22753 18748
rect 22152 18708 22158 18720
rect 22741 18717 22753 18720
rect 22787 18717 22799 18751
rect 22741 18711 22799 18717
rect 23661 18751 23719 18757
rect 23661 18717 23673 18751
rect 23707 18748 23719 18751
rect 24210 18748 24216 18760
rect 23707 18720 24216 18748
rect 23707 18717 23719 18720
rect 23661 18711 23719 18717
rect 24210 18708 24216 18720
rect 24268 18708 24274 18760
rect 16206 18680 16212 18692
rect 16119 18652 16212 18680
rect 16206 18640 16212 18652
rect 16264 18680 16270 18692
rect 16264 18652 18828 18680
rect 16264 18640 16270 18652
rect 18800 18624 18828 18652
rect 20162 18640 20168 18692
rect 20220 18680 20226 18692
rect 20349 18683 20407 18689
rect 20349 18680 20361 18683
rect 20220 18652 20361 18680
rect 20220 18640 20226 18652
rect 20349 18649 20361 18652
rect 20395 18649 20407 18683
rect 20349 18643 20407 18649
rect 20441 18683 20499 18689
rect 20441 18649 20453 18683
rect 20487 18680 20499 18683
rect 20993 18683 21051 18689
rect 20993 18680 21005 18683
rect 20487 18652 21005 18680
rect 20487 18649 20499 18652
rect 20441 18643 20499 18649
rect 20993 18649 21005 18652
rect 21039 18649 21051 18683
rect 37458 18680 37464 18692
rect 20993 18643 21051 18649
rect 22296 18652 37464 18680
rect 17126 18572 17132 18624
rect 17184 18612 17190 18624
rect 17405 18615 17463 18621
rect 17405 18612 17417 18615
rect 17184 18584 17417 18612
rect 17184 18572 17190 18584
rect 17405 18581 17417 18584
rect 17451 18581 17463 18615
rect 18782 18612 18788 18624
rect 18743 18584 18788 18612
rect 17405 18575 17463 18581
rect 18782 18572 18788 18584
rect 18840 18572 18846 18624
rect 22296 18621 22324 18652
rect 37458 18640 37464 18652
rect 37516 18640 37522 18692
rect 22281 18615 22339 18621
rect 22281 18581 22293 18615
rect 22327 18581 22339 18615
rect 22281 18575 22339 18581
rect 23474 18572 23480 18624
rect 23532 18612 23538 18624
rect 23569 18615 23627 18621
rect 23569 18612 23581 18615
rect 23532 18584 23581 18612
rect 23532 18572 23538 18584
rect 23569 18581 23581 18584
rect 23615 18581 23627 18615
rect 24578 18612 24584 18624
rect 24539 18584 24584 18612
rect 23569 18575 23627 18581
rect 24578 18572 24584 18584
rect 24636 18572 24642 18624
rect 25225 18615 25283 18621
rect 25225 18581 25237 18615
rect 25271 18612 25283 18615
rect 25958 18612 25964 18624
rect 25271 18584 25964 18612
rect 25271 18581 25283 18584
rect 25225 18575 25283 18581
rect 25958 18572 25964 18584
rect 26016 18572 26022 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 1762 18408 1768 18420
rect 1723 18380 1768 18408
rect 1762 18368 1768 18380
rect 1820 18368 1826 18420
rect 4614 18408 4620 18420
rect 4575 18380 4620 18408
rect 4614 18368 4620 18380
rect 4672 18368 4678 18420
rect 20990 18408 20996 18420
rect 18892 18380 20996 18408
rect 18892 18349 18920 18380
rect 20990 18368 20996 18380
rect 21048 18368 21054 18420
rect 24210 18408 24216 18420
rect 21284 18380 24216 18408
rect 16209 18343 16267 18349
rect 16209 18309 16221 18343
rect 16255 18340 16267 18343
rect 17037 18343 17095 18349
rect 17037 18340 17049 18343
rect 16255 18312 17049 18340
rect 16255 18309 16267 18312
rect 16209 18303 16267 18309
rect 17037 18309 17049 18312
rect 17083 18309 17095 18343
rect 17037 18303 17095 18309
rect 18877 18343 18935 18349
rect 18877 18309 18889 18343
rect 18923 18309 18935 18343
rect 20070 18340 20076 18352
rect 20031 18312 20076 18340
rect 18877 18303 18935 18309
rect 20070 18300 20076 18312
rect 20128 18300 20134 18352
rect 1578 18232 1584 18284
rect 1636 18272 1642 18284
rect 1673 18275 1731 18281
rect 1673 18272 1685 18275
rect 1636 18244 1685 18272
rect 1636 18232 1642 18244
rect 1673 18241 1685 18244
rect 1719 18241 1731 18275
rect 1673 18235 1731 18241
rect 4801 18275 4859 18281
rect 4801 18241 4813 18275
rect 4847 18272 4859 18275
rect 15657 18275 15715 18281
rect 4847 18244 5396 18272
rect 4847 18241 4859 18244
rect 4801 18235 4859 18241
rect 5368 18077 5396 18244
rect 15657 18241 15669 18275
rect 15703 18272 15715 18275
rect 16114 18272 16120 18284
rect 15703 18244 16120 18272
rect 15703 18241 15715 18244
rect 15657 18235 15715 18241
rect 16114 18232 16120 18244
rect 16172 18232 16178 18284
rect 21284 18281 21312 18380
rect 24210 18368 24216 18380
rect 24268 18368 24274 18420
rect 26878 18368 26884 18420
rect 26936 18408 26942 18420
rect 37734 18408 37740 18420
rect 26936 18380 37740 18408
rect 26936 18368 26942 18380
rect 37734 18368 37740 18380
rect 37792 18368 37798 18420
rect 22554 18340 22560 18352
rect 22515 18312 22560 18340
rect 22554 18300 22560 18312
rect 22612 18300 22618 18352
rect 22646 18300 22652 18352
rect 22704 18340 22710 18352
rect 22704 18312 22749 18340
rect 22704 18300 22710 18312
rect 21269 18275 21327 18281
rect 21269 18241 21281 18275
rect 21315 18241 21327 18275
rect 23750 18272 23756 18284
rect 23711 18244 23756 18272
rect 21269 18235 21327 18241
rect 23750 18232 23756 18244
rect 23808 18232 23814 18284
rect 24578 18272 24584 18284
rect 24491 18244 24584 18272
rect 24578 18232 24584 18244
rect 24636 18272 24642 18284
rect 25041 18275 25099 18281
rect 25041 18272 25053 18275
rect 24636 18244 25053 18272
rect 24636 18232 24642 18244
rect 25041 18241 25053 18244
rect 25087 18272 25099 18275
rect 25685 18275 25743 18281
rect 25685 18272 25697 18275
rect 25087 18244 25697 18272
rect 25087 18241 25099 18244
rect 25041 18235 25099 18241
rect 25685 18241 25697 18244
rect 25731 18241 25743 18275
rect 25685 18235 25743 18241
rect 16942 18204 16948 18216
rect 16903 18176 16948 18204
rect 16942 18164 16948 18176
rect 17000 18204 17006 18216
rect 18785 18207 18843 18213
rect 18785 18204 18797 18207
rect 17000 18176 18797 18204
rect 17000 18164 17006 18176
rect 18785 18173 18797 18176
rect 18831 18173 18843 18207
rect 19978 18204 19984 18216
rect 19939 18176 19984 18204
rect 18785 18167 18843 18173
rect 19978 18164 19984 18176
rect 20036 18164 20042 18216
rect 23382 18164 23388 18216
rect 23440 18204 23446 18216
rect 24596 18204 24624 18232
rect 23440 18176 24624 18204
rect 23440 18164 23446 18176
rect 17402 18096 17408 18148
rect 17460 18136 17466 18148
rect 17497 18139 17555 18145
rect 17497 18136 17509 18139
rect 17460 18108 17509 18136
rect 17460 18096 17466 18108
rect 17497 18105 17509 18108
rect 17543 18105 17555 18139
rect 19334 18136 19340 18148
rect 19295 18108 19340 18136
rect 17497 18099 17555 18105
rect 19334 18096 19340 18108
rect 19392 18096 19398 18148
rect 20530 18136 20536 18148
rect 20491 18108 20536 18136
rect 20530 18096 20536 18108
rect 20588 18096 20594 18148
rect 22097 18139 22155 18145
rect 22097 18136 22109 18139
rect 20640 18108 22109 18136
rect 5353 18071 5411 18077
rect 5353 18037 5365 18071
rect 5399 18068 5411 18071
rect 8018 18068 8024 18080
rect 5399 18040 8024 18068
rect 5399 18037 5411 18040
rect 5353 18031 5411 18037
rect 8018 18028 8024 18040
rect 8076 18068 8082 18080
rect 11146 18068 11152 18080
rect 8076 18040 11152 18068
rect 8076 18028 8082 18040
rect 11146 18028 11152 18040
rect 11204 18028 11210 18080
rect 18230 18068 18236 18080
rect 18191 18040 18236 18068
rect 18230 18028 18236 18040
rect 18288 18028 18294 18080
rect 19150 18028 19156 18080
rect 19208 18068 19214 18080
rect 20640 18068 20668 18108
rect 22097 18105 22109 18108
rect 22143 18105 22155 18139
rect 22097 18099 22155 18105
rect 23845 18139 23903 18145
rect 23845 18105 23857 18139
rect 23891 18136 23903 18139
rect 25038 18136 25044 18148
rect 23891 18108 25044 18136
rect 23891 18105 23903 18108
rect 23845 18099 23903 18105
rect 25038 18096 25044 18108
rect 25096 18096 25102 18148
rect 21174 18068 21180 18080
rect 19208 18040 20668 18068
rect 21135 18040 21180 18068
rect 19208 18028 19214 18040
rect 21174 18028 21180 18040
rect 21232 18028 21238 18080
rect 22278 18028 22284 18080
rect 22336 18068 22342 18080
rect 23290 18068 23296 18080
rect 22336 18040 23296 18068
rect 22336 18028 22342 18040
rect 23290 18028 23296 18040
rect 23348 18028 23354 18080
rect 24026 18028 24032 18080
rect 24084 18068 24090 18080
rect 24489 18071 24547 18077
rect 24489 18068 24501 18071
rect 24084 18040 24501 18068
rect 24084 18028 24090 18040
rect 24489 18037 24501 18040
rect 24535 18037 24547 18071
rect 25130 18068 25136 18080
rect 25091 18040 25136 18068
rect 24489 18031 24547 18037
rect 25130 18028 25136 18040
rect 25188 18028 25194 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 22373 17867 22431 17873
rect 15672 17836 21588 17864
rect 1578 17796 1584 17808
rect 1539 17768 1584 17796
rect 1578 17756 1584 17768
rect 1636 17756 1642 17808
rect 14461 17663 14519 17669
rect 14461 17629 14473 17663
rect 14507 17660 14519 17663
rect 14918 17660 14924 17672
rect 14507 17632 14924 17660
rect 14507 17629 14519 17632
rect 14461 17623 14519 17629
rect 14918 17620 14924 17632
rect 14976 17620 14982 17672
rect 15672 17669 15700 17836
rect 15930 17756 15936 17808
rect 15988 17796 15994 17808
rect 15988 17768 20944 17796
rect 15988 17756 15994 17768
rect 16684 17700 18276 17728
rect 16684 17669 16712 17700
rect 18248 17672 18276 17700
rect 18414 17688 18420 17740
rect 18472 17728 18478 17740
rect 19886 17728 19892 17740
rect 18472 17700 19892 17728
rect 18472 17688 18478 17700
rect 19886 17688 19892 17700
rect 19944 17688 19950 17740
rect 20254 17688 20260 17740
rect 20312 17728 20318 17740
rect 20622 17728 20628 17740
rect 20312 17700 20357 17728
rect 20583 17700 20628 17728
rect 20312 17688 20318 17700
rect 20622 17688 20628 17700
rect 20680 17688 20686 17740
rect 15013 17663 15071 17669
rect 15013 17629 15025 17663
rect 15059 17660 15071 17663
rect 15657 17663 15715 17669
rect 15657 17660 15669 17663
rect 15059 17632 15669 17660
rect 15059 17629 15071 17632
rect 15013 17623 15071 17629
rect 15657 17629 15669 17632
rect 15703 17629 15715 17663
rect 15657 17623 15715 17629
rect 16669 17663 16727 17669
rect 16669 17629 16681 17663
rect 16715 17629 16727 17663
rect 16669 17623 16727 17629
rect 17126 17620 17132 17672
rect 17184 17660 17190 17672
rect 17313 17663 17371 17669
rect 17313 17660 17325 17663
rect 17184 17632 17325 17660
rect 17184 17620 17190 17632
rect 17313 17629 17325 17632
rect 17359 17629 17371 17663
rect 17313 17623 17371 17629
rect 18230 17620 18236 17672
rect 18288 17660 18294 17672
rect 18325 17663 18383 17669
rect 18325 17660 18337 17663
rect 18288 17632 18337 17660
rect 18288 17620 18294 17632
rect 18325 17629 18337 17632
rect 18371 17660 18383 17663
rect 18690 17660 18696 17672
rect 18371 17632 18696 17660
rect 18371 17629 18383 17632
rect 18325 17623 18383 17629
rect 18690 17620 18696 17632
rect 18748 17620 18754 17672
rect 19521 17663 19579 17669
rect 19521 17629 19533 17663
rect 19567 17660 19579 17663
rect 20070 17660 20076 17672
rect 19567 17632 20076 17660
rect 19567 17629 19579 17632
rect 19521 17623 19579 17629
rect 11238 17552 11244 17604
rect 11296 17592 11302 17604
rect 16758 17592 16764 17604
rect 11296 17564 16764 17592
rect 11296 17552 11302 17564
rect 16758 17552 16764 17564
rect 16816 17552 16822 17604
rect 17865 17595 17923 17601
rect 17865 17561 17877 17595
rect 17911 17592 17923 17595
rect 19536 17592 19564 17623
rect 20070 17620 20076 17632
rect 20128 17620 20134 17672
rect 17911 17564 19564 17592
rect 19613 17595 19671 17601
rect 17911 17561 17923 17564
rect 17865 17555 17923 17561
rect 19613 17561 19625 17595
rect 19659 17561 19671 17595
rect 19613 17555 19671 17561
rect 20349 17595 20407 17601
rect 20349 17561 20361 17595
rect 20395 17561 20407 17595
rect 20916 17592 20944 17768
rect 21560 17728 21588 17836
rect 22373 17833 22385 17867
rect 22419 17864 22431 17867
rect 22554 17864 22560 17876
rect 22419 17836 22560 17864
rect 22419 17833 22431 17836
rect 22373 17827 22431 17833
rect 22554 17824 22560 17836
rect 22612 17824 22618 17876
rect 23290 17824 23296 17876
rect 23348 17864 23354 17876
rect 27062 17864 27068 17876
rect 23348 17836 27068 17864
rect 23348 17824 23354 17836
rect 27062 17824 27068 17836
rect 27120 17824 27126 17876
rect 24673 17799 24731 17805
rect 24673 17796 24685 17799
rect 22572 17768 24685 17796
rect 22370 17728 22376 17740
rect 21560 17700 22376 17728
rect 21560 17669 21588 17700
rect 22370 17688 22376 17700
rect 22428 17688 22434 17740
rect 21545 17663 21603 17669
rect 21545 17629 21557 17663
rect 21591 17629 21603 17663
rect 21545 17623 21603 17629
rect 21634 17620 21640 17672
rect 21692 17660 21698 17672
rect 22278 17660 22284 17672
rect 21692 17632 22284 17660
rect 21692 17620 21698 17632
rect 22278 17620 22284 17632
rect 22336 17620 22342 17672
rect 22572 17592 22600 17768
rect 24673 17765 24685 17768
rect 24719 17796 24731 17799
rect 25866 17796 25872 17808
rect 24719 17768 25872 17796
rect 24719 17765 24731 17768
rect 24673 17759 24731 17765
rect 25866 17756 25872 17768
rect 25924 17756 25930 17808
rect 22646 17688 22652 17740
rect 22704 17728 22710 17740
rect 23017 17731 23075 17737
rect 23017 17728 23029 17731
rect 22704 17700 23029 17728
rect 22704 17688 22710 17700
rect 23017 17697 23029 17700
rect 23063 17697 23075 17731
rect 23017 17691 23075 17697
rect 23198 17688 23204 17740
rect 23256 17728 23262 17740
rect 23750 17728 23756 17740
rect 23256 17700 23756 17728
rect 23256 17688 23262 17700
rect 23750 17688 23756 17700
rect 23808 17728 23814 17740
rect 26878 17728 26884 17740
rect 23808 17700 26884 17728
rect 23808 17688 23814 17700
rect 26878 17688 26884 17700
rect 26936 17688 26942 17740
rect 25958 17660 25964 17672
rect 25919 17632 25964 17660
rect 25958 17620 25964 17632
rect 26016 17660 26022 17672
rect 26421 17663 26479 17669
rect 26421 17660 26433 17663
rect 26016 17632 26433 17660
rect 26016 17620 26022 17632
rect 26421 17629 26433 17632
rect 26467 17629 26479 17663
rect 26421 17623 26479 17629
rect 20916 17564 22600 17592
rect 23109 17595 23167 17601
rect 20349 17555 20407 17561
rect 23109 17561 23121 17595
rect 23155 17592 23167 17595
rect 23474 17592 23480 17604
rect 23155 17564 23480 17592
rect 23155 17561 23167 17564
rect 23109 17555 23167 17561
rect 15378 17484 15384 17536
rect 15436 17524 15442 17536
rect 15565 17527 15623 17533
rect 15565 17524 15577 17527
rect 15436 17496 15577 17524
rect 15436 17484 15442 17496
rect 15565 17493 15577 17496
rect 15611 17493 15623 17527
rect 15565 17487 15623 17493
rect 16577 17527 16635 17533
rect 16577 17493 16589 17527
rect 16623 17524 16635 17527
rect 16666 17524 16672 17536
rect 16623 17496 16672 17524
rect 16623 17493 16635 17496
rect 16577 17487 16635 17493
rect 16666 17484 16672 17496
rect 16724 17484 16730 17536
rect 17221 17527 17279 17533
rect 17221 17493 17233 17527
rect 17267 17524 17279 17527
rect 17494 17524 17500 17536
rect 17267 17496 17500 17524
rect 17267 17493 17279 17496
rect 17221 17487 17279 17493
rect 17494 17484 17500 17496
rect 17552 17484 17558 17536
rect 18417 17527 18475 17533
rect 18417 17493 18429 17527
rect 18463 17524 18475 17527
rect 18598 17524 18604 17536
rect 18463 17496 18604 17524
rect 18463 17493 18475 17496
rect 18417 17487 18475 17493
rect 18598 17484 18604 17496
rect 18656 17484 18662 17536
rect 19628 17524 19656 17555
rect 20364 17524 20392 17555
rect 23474 17552 23480 17564
rect 23532 17552 23538 17604
rect 23661 17595 23719 17601
rect 23661 17561 23673 17595
rect 23707 17592 23719 17595
rect 24302 17592 24308 17604
rect 23707 17564 24308 17592
rect 23707 17561 23719 17564
rect 23661 17555 23719 17561
rect 24302 17552 24308 17564
rect 24360 17552 24366 17604
rect 25038 17552 25044 17604
rect 25096 17592 25102 17604
rect 25133 17595 25191 17601
rect 25133 17592 25145 17595
rect 25096 17564 25145 17592
rect 25096 17552 25102 17564
rect 25133 17561 25145 17564
rect 25179 17561 25191 17595
rect 25133 17555 25191 17561
rect 25222 17552 25228 17604
rect 25280 17592 25286 17604
rect 25280 17564 25325 17592
rect 25280 17552 25286 17564
rect 19628 17496 20392 17524
rect 20714 17484 20720 17536
rect 20772 17524 20778 17536
rect 21453 17527 21511 17533
rect 21453 17524 21465 17527
rect 20772 17496 21465 17524
rect 20772 17484 20778 17496
rect 21453 17493 21465 17496
rect 21499 17493 21511 17527
rect 21453 17487 21511 17493
rect 25406 17484 25412 17536
rect 25464 17524 25470 17536
rect 25869 17527 25927 17533
rect 25869 17524 25881 17527
rect 25464 17496 25881 17524
rect 25464 17484 25470 17496
rect 25869 17493 25881 17496
rect 25915 17493 25927 17527
rect 27062 17524 27068 17536
rect 27023 17496 27068 17524
rect 25869 17487 25927 17493
rect 27062 17484 27068 17496
rect 27120 17484 27126 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 19886 17320 19892 17332
rect 16684 17292 19892 17320
rect 12802 17212 12808 17264
rect 12860 17252 12866 17264
rect 16022 17252 16028 17264
rect 12860 17224 16028 17252
rect 12860 17212 12866 17224
rect 16022 17212 16028 17224
rect 16080 17212 16086 17264
rect 16117 17255 16175 17261
rect 16117 17221 16129 17255
rect 16163 17252 16175 17255
rect 16574 17252 16580 17264
rect 16163 17224 16580 17252
rect 16163 17221 16175 17224
rect 16117 17215 16175 17221
rect 16574 17212 16580 17224
rect 16632 17212 16638 17264
rect 14461 17187 14519 17193
rect 14461 17153 14473 17187
rect 14507 17153 14519 17187
rect 14918 17184 14924 17196
rect 14879 17156 14924 17184
rect 14461 17147 14519 17153
rect 14476 17116 14504 17147
rect 14918 17144 14924 17156
rect 14976 17144 14982 17196
rect 15838 17116 15844 17128
rect 14476 17088 15844 17116
rect 15838 17076 15844 17088
rect 15896 17076 15902 17128
rect 15930 17076 15936 17128
rect 15988 17116 15994 17128
rect 16209 17119 16267 17125
rect 15988 17088 16033 17116
rect 15988 17076 15994 17088
rect 16209 17085 16221 17119
rect 16255 17116 16267 17119
rect 16684 17116 16712 17292
rect 19886 17280 19892 17292
rect 19944 17320 19950 17332
rect 20346 17320 20352 17332
rect 19944 17292 20352 17320
rect 19944 17280 19950 17292
rect 20346 17280 20352 17292
rect 20404 17280 20410 17332
rect 20990 17320 20996 17332
rect 20951 17292 20996 17320
rect 20990 17280 20996 17292
rect 21048 17280 21054 17332
rect 27338 17320 27344 17332
rect 23216 17292 27344 17320
rect 17037 17255 17095 17261
rect 17037 17221 17049 17255
rect 17083 17252 17095 17255
rect 18322 17252 18328 17264
rect 17083 17224 18328 17252
rect 17083 17221 17095 17224
rect 17037 17215 17095 17221
rect 18322 17212 18328 17224
rect 18380 17212 18386 17264
rect 18782 17252 18788 17264
rect 18616 17224 18788 17252
rect 18414 17184 18420 17196
rect 17604 17156 18420 17184
rect 16255 17088 16712 17116
rect 16255 17085 16267 17088
rect 16209 17079 16267 17085
rect 16758 17076 16764 17128
rect 16816 17116 16822 17128
rect 16945 17119 17003 17125
rect 16945 17116 16957 17119
rect 16816 17088 16957 17116
rect 16816 17076 16822 17088
rect 16945 17085 16957 17088
rect 16991 17085 17003 17119
rect 17604 17116 17632 17156
rect 18414 17144 18420 17156
rect 18472 17144 18478 17196
rect 18616 17193 18644 17224
rect 18782 17212 18788 17224
rect 18840 17252 18846 17264
rect 19702 17252 19708 17264
rect 18840 17224 19708 17252
rect 18840 17212 18846 17224
rect 19702 17212 19708 17224
rect 19760 17212 19766 17264
rect 19797 17255 19855 17261
rect 19797 17221 19809 17255
rect 19843 17252 19855 17255
rect 21174 17252 21180 17264
rect 19843 17224 21180 17252
rect 19843 17221 19855 17224
rect 19797 17215 19855 17221
rect 21174 17212 21180 17224
rect 21232 17212 21238 17264
rect 18601 17187 18659 17193
rect 18601 17153 18613 17187
rect 18647 17153 18659 17187
rect 21082 17184 21088 17196
rect 21043 17156 21088 17184
rect 18601 17147 18659 17153
rect 21082 17144 21088 17156
rect 21140 17144 21146 17196
rect 22281 17187 22339 17193
rect 22281 17153 22293 17187
rect 22327 17184 22339 17187
rect 23216 17184 23244 17292
rect 27338 17280 27344 17292
rect 27396 17280 27402 17332
rect 23477 17255 23535 17261
rect 23477 17221 23489 17255
rect 23523 17252 23535 17255
rect 24581 17255 24639 17261
rect 24581 17252 24593 17255
rect 23523 17224 24593 17252
rect 23523 17221 23535 17224
rect 23477 17215 23535 17221
rect 24581 17221 24593 17224
rect 24627 17221 24639 17255
rect 25406 17252 25412 17264
rect 25367 17224 25412 17252
rect 24581 17215 24639 17221
rect 25406 17212 25412 17224
rect 25464 17212 25470 17264
rect 27154 17252 27160 17264
rect 25976 17224 27160 17252
rect 22327 17156 23244 17184
rect 22327 17153 22339 17156
rect 22281 17147 22339 17153
rect 16945 17079 17003 17085
rect 17052 17088 17632 17116
rect 18141 17119 18199 17125
rect 15654 17008 15660 17060
rect 15712 17048 15718 17060
rect 15948 17048 15976 17076
rect 15712 17020 15976 17048
rect 15712 17008 15718 17020
rect 16022 17008 16028 17060
rect 16080 17048 16086 17060
rect 17052 17048 17080 17088
rect 18141 17085 18153 17119
rect 18187 17116 18199 17119
rect 19610 17116 19616 17128
rect 18187 17088 19616 17116
rect 18187 17085 18199 17088
rect 18141 17079 18199 17085
rect 19610 17076 19616 17088
rect 19668 17076 19674 17128
rect 19886 17116 19892 17128
rect 19847 17088 19892 17116
rect 19886 17076 19892 17088
rect 19944 17076 19950 17128
rect 16080 17020 17080 17048
rect 17497 17051 17555 17057
rect 16080 17008 16086 17020
rect 17497 17017 17509 17051
rect 17543 17048 17555 17051
rect 17862 17048 17868 17060
rect 17543 17020 17868 17048
rect 17543 17017 17555 17020
rect 17497 17011 17555 17017
rect 17862 17008 17868 17020
rect 17920 17008 17926 17060
rect 19334 17048 19340 17060
rect 19295 17020 19340 17048
rect 19334 17008 19340 17020
rect 19392 17008 19398 17060
rect 21450 17008 21456 17060
rect 21508 17048 21514 17060
rect 22296 17048 22324 17147
rect 24394 17144 24400 17196
rect 24452 17184 24458 17196
rect 24673 17187 24731 17193
rect 24673 17184 24685 17187
rect 24452 17156 24685 17184
rect 24452 17144 24458 17156
rect 24673 17153 24685 17156
rect 24719 17153 24731 17187
rect 24673 17147 24731 17153
rect 22370 17076 22376 17128
rect 22428 17116 22434 17128
rect 22830 17116 22836 17128
rect 22428 17088 22836 17116
rect 22428 17076 22434 17088
rect 22830 17076 22836 17088
rect 22888 17076 22894 17128
rect 23382 17116 23388 17128
rect 23343 17088 23388 17116
rect 23382 17076 23388 17088
rect 23440 17076 23446 17128
rect 24029 17119 24087 17125
rect 24029 17085 24041 17119
rect 24075 17116 24087 17119
rect 24302 17116 24308 17128
rect 24075 17088 24308 17116
rect 24075 17085 24087 17088
rect 24029 17079 24087 17085
rect 24302 17076 24308 17088
rect 24360 17076 24366 17128
rect 25314 17116 25320 17128
rect 25275 17088 25320 17116
rect 25314 17076 25320 17088
rect 25372 17076 25378 17128
rect 25976 17116 26004 17224
rect 27154 17212 27160 17224
rect 27212 17212 27218 17264
rect 26605 17187 26663 17193
rect 26605 17153 26617 17187
rect 26651 17184 26663 17187
rect 27062 17184 27068 17196
rect 26651 17156 27068 17184
rect 26651 17153 26663 17156
rect 26605 17147 26663 17153
rect 27062 17144 27068 17156
rect 27120 17144 27126 17196
rect 37553 17187 37611 17193
rect 37553 17153 37565 17187
rect 37599 17184 37611 17187
rect 38194 17184 38200 17196
rect 37599 17156 38200 17184
rect 37599 17153 37611 17156
rect 37553 17147 37611 17153
rect 38194 17144 38200 17156
rect 38252 17144 38258 17196
rect 25424 17088 26004 17116
rect 21508 17020 22324 17048
rect 21508 17008 21514 17020
rect 13170 16980 13176 16992
rect 13131 16952 13176 16980
rect 13170 16940 13176 16952
rect 13228 16940 13234 16992
rect 13814 16980 13820 16992
rect 13775 16952 13820 16980
rect 13814 16940 13820 16952
rect 13872 16940 13878 16992
rect 14182 16940 14188 16992
rect 14240 16980 14246 16992
rect 14369 16983 14427 16989
rect 14369 16980 14381 16983
rect 14240 16952 14381 16980
rect 14240 16940 14246 16952
rect 14369 16949 14381 16952
rect 14415 16949 14427 16983
rect 14369 16943 14427 16949
rect 15013 16983 15071 16989
rect 15013 16949 15025 16983
rect 15059 16980 15071 16983
rect 16390 16980 16396 16992
rect 15059 16952 16396 16980
rect 15059 16949 15071 16952
rect 15013 16943 15071 16949
rect 16390 16940 16396 16952
rect 16448 16940 16454 16992
rect 18693 16983 18751 16989
rect 18693 16949 18705 16983
rect 18739 16980 18751 16983
rect 20990 16980 20996 16992
rect 18739 16952 20996 16980
rect 18739 16949 18751 16952
rect 18693 16943 18751 16949
rect 20990 16940 20996 16952
rect 21048 16940 21054 16992
rect 22186 16940 22192 16992
rect 22244 16980 22250 16992
rect 22244 16952 22289 16980
rect 22244 16940 22250 16952
rect 22646 16940 22652 16992
rect 22704 16980 22710 16992
rect 25424 16980 25452 17088
rect 26234 17076 26240 17128
rect 26292 17116 26298 17128
rect 27157 17119 27215 17125
rect 27157 17116 27169 17119
rect 26292 17088 27169 17116
rect 26292 17076 26298 17088
rect 27157 17085 27169 17088
rect 27203 17085 27215 17119
rect 27157 17079 27215 17085
rect 25869 17051 25927 17057
rect 25869 17017 25881 17051
rect 25915 17048 25927 17051
rect 26050 17048 26056 17060
rect 25915 17020 26056 17048
rect 25915 17017 25927 17020
rect 25869 17011 25927 17017
rect 26050 17008 26056 17020
rect 26108 17048 26114 17060
rect 27798 17048 27804 17060
rect 26108 17020 27804 17048
rect 26108 17008 26114 17020
rect 27798 17008 27804 17020
rect 27856 17008 27862 17060
rect 35894 17008 35900 17060
rect 35952 17048 35958 17060
rect 38013 17051 38071 17057
rect 38013 17048 38025 17051
rect 35952 17020 38025 17048
rect 35952 17008 35958 17020
rect 38013 17017 38025 17020
rect 38059 17017 38071 17051
rect 38013 17011 38071 17017
rect 22704 16952 25452 16980
rect 22704 16940 22710 16952
rect 26142 16940 26148 16992
rect 26200 16980 26206 16992
rect 26513 16983 26571 16989
rect 26513 16980 26525 16983
rect 26200 16952 26525 16980
rect 26200 16940 26206 16952
rect 26513 16949 26525 16952
rect 26559 16949 26571 16983
rect 26513 16943 26571 16949
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 2222 16736 2228 16788
rect 2280 16776 2286 16788
rect 19521 16779 19579 16785
rect 19521 16776 19533 16779
rect 2280 16748 19533 16776
rect 2280 16736 2286 16748
rect 19521 16745 19533 16748
rect 19567 16745 19579 16779
rect 19521 16739 19579 16745
rect 20162 16736 20168 16788
rect 20220 16776 20226 16788
rect 23198 16776 23204 16788
rect 20220 16748 23204 16776
rect 20220 16736 20226 16748
rect 23198 16736 23204 16748
rect 23256 16736 23262 16788
rect 25148 16748 27200 16776
rect 13648 16680 15332 16708
rect 13648 16640 13676 16680
rect 15304 16652 15332 16680
rect 15838 16668 15844 16720
rect 15896 16708 15902 16720
rect 15896 16680 17172 16708
rect 15896 16668 15902 16680
rect 14366 16640 14372 16652
rect 13556 16612 13676 16640
rect 14327 16612 14372 16640
rect 13081 16575 13139 16581
rect 13081 16572 13093 16575
rect 12728 16544 13093 16572
rect 8202 16464 8208 16516
rect 8260 16504 8266 16516
rect 12618 16504 12624 16516
rect 8260 16476 12624 16504
rect 8260 16464 8266 16476
rect 12618 16464 12624 16476
rect 12676 16464 12682 16516
rect 12728 16448 12756 16544
rect 13081 16541 13093 16544
rect 13127 16572 13139 16575
rect 13170 16572 13176 16584
rect 13127 16544 13176 16572
rect 13127 16541 13139 16544
rect 13081 16535 13139 16541
rect 13170 16532 13176 16544
rect 13228 16532 13234 16584
rect 13556 16581 13584 16612
rect 14366 16600 14372 16612
rect 14424 16600 14430 16652
rect 15286 16600 15292 16652
rect 15344 16640 15350 16652
rect 16206 16640 16212 16652
rect 15344 16612 15976 16640
rect 15344 16600 15350 16612
rect 13541 16575 13599 16581
rect 13541 16541 13553 16575
rect 13587 16541 13599 16575
rect 13541 16535 13599 16541
rect 14458 16464 14464 16516
rect 14516 16504 14522 16516
rect 15010 16504 15016 16516
rect 14516 16476 14561 16504
rect 14971 16476 15016 16504
rect 14516 16464 14522 16476
rect 15010 16464 15016 16476
rect 15068 16464 15074 16516
rect 15948 16504 15976 16612
rect 16040 16612 16212 16640
rect 16040 16581 16068 16612
rect 16206 16600 16212 16612
rect 16264 16600 16270 16652
rect 16025 16575 16083 16581
rect 16025 16541 16037 16575
rect 16071 16541 16083 16575
rect 16574 16572 16580 16584
rect 16535 16544 16580 16572
rect 16025 16535 16083 16541
rect 16574 16532 16580 16544
rect 16632 16532 16638 16584
rect 17144 16581 17172 16680
rect 17586 16668 17592 16720
rect 17644 16708 17650 16720
rect 18046 16708 18052 16720
rect 17644 16680 18052 16708
rect 17644 16668 17650 16680
rect 18046 16668 18052 16680
rect 18104 16668 18110 16720
rect 19702 16668 19708 16720
rect 19760 16708 19766 16720
rect 20809 16711 20867 16717
rect 19760 16680 20576 16708
rect 19760 16668 19766 16680
rect 17862 16640 17868 16652
rect 17775 16612 17868 16640
rect 17862 16600 17868 16612
rect 17920 16640 17926 16652
rect 20438 16640 20444 16652
rect 17920 16612 20444 16640
rect 17920 16600 17926 16612
rect 20438 16600 20444 16612
rect 20496 16600 20502 16652
rect 20548 16640 20576 16680
rect 20809 16677 20821 16711
rect 20855 16708 20867 16711
rect 20898 16708 20904 16720
rect 20855 16680 20904 16708
rect 20855 16677 20867 16680
rect 20809 16671 20867 16677
rect 20898 16668 20904 16680
rect 20956 16708 20962 16720
rect 22281 16711 22339 16717
rect 22281 16708 22293 16711
rect 20956 16680 22293 16708
rect 20956 16668 20962 16680
rect 22281 16677 22293 16680
rect 22327 16677 22339 16711
rect 25148 16708 25176 16748
rect 25774 16708 25780 16720
rect 22281 16671 22339 16677
rect 22572 16680 25176 16708
rect 25240 16680 25780 16708
rect 22572 16652 22600 16680
rect 22554 16640 22560 16652
rect 20548 16612 22560 16640
rect 22554 16600 22560 16612
rect 22612 16600 22618 16652
rect 24854 16640 24860 16652
rect 23492 16612 24860 16640
rect 16669 16575 16727 16581
rect 16669 16541 16681 16575
rect 16715 16541 16727 16575
rect 16669 16535 16727 16541
rect 17129 16575 17187 16581
rect 17129 16541 17141 16575
rect 17175 16541 17187 16575
rect 21542 16572 21548 16584
rect 21503 16544 21548 16572
rect 17129 16535 17187 16541
rect 16684 16504 16712 16535
rect 21542 16532 21548 16544
rect 21600 16572 21606 16584
rect 21600 16544 22232 16572
rect 21600 16532 21606 16544
rect 15948 16476 16712 16504
rect 17957 16507 18015 16513
rect 17957 16473 17969 16507
rect 18003 16473 18015 16507
rect 17957 16467 18015 16473
rect 11238 16396 11244 16448
rect 11296 16436 11302 16448
rect 11425 16439 11483 16445
rect 11425 16436 11437 16439
rect 11296 16408 11437 16436
rect 11296 16396 11302 16408
rect 11425 16405 11437 16408
rect 11471 16405 11483 16439
rect 11425 16399 11483 16405
rect 12437 16439 12495 16445
rect 12437 16405 12449 16439
rect 12483 16436 12495 16439
rect 12710 16436 12716 16448
rect 12483 16408 12716 16436
rect 12483 16405 12495 16408
rect 12437 16399 12495 16405
rect 12710 16396 12716 16408
rect 12768 16396 12774 16448
rect 12986 16436 12992 16448
rect 12947 16408 12992 16436
rect 12986 16396 12992 16408
rect 13044 16396 13050 16448
rect 13633 16439 13691 16445
rect 13633 16405 13645 16439
rect 13679 16436 13691 16439
rect 14550 16436 14556 16448
rect 13679 16408 14556 16436
rect 13679 16405 13691 16408
rect 13633 16399 13691 16405
rect 14550 16396 14556 16408
rect 14608 16396 14614 16448
rect 15746 16396 15752 16448
rect 15804 16436 15810 16448
rect 15933 16439 15991 16445
rect 15933 16436 15945 16439
rect 15804 16408 15945 16436
rect 15804 16396 15810 16408
rect 15933 16405 15945 16408
rect 15979 16405 15991 16439
rect 17218 16436 17224 16448
rect 17179 16408 17224 16436
rect 15933 16399 15991 16405
rect 17218 16396 17224 16408
rect 17276 16396 17282 16448
rect 17678 16396 17684 16448
rect 17736 16436 17742 16448
rect 17972 16436 18000 16467
rect 18046 16464 18052 16516
rect 18104 16504 18110 16516
rect 18877 16507 18935 16513
rect 18877 16504 18889 16507
rect 18104 16476 18889 16504
rect 18104 16464 18110 16476
rect 18877 16473 18889 16476
rect 18923 16473 18935 16507
rect 19610 16504 19616 16516
rect 19523 16476 19616 16504
rect 18877 16467 18935 16473
rect 17736 16408 18000 16436
rect 18892 16436 18920 16467
rect 19610 16464 19616 16476
rect 19668 16504 19674 16516
rect 20070 16504 20076 16516
rect 19668 16476 20076 16504
rect 19668 16464 19674 16476
rect 20070 16464 20076 16476
rect 20128 16464 20134 16516
rect 20254 16504 20260 16516
rect 20215 16476 20260 16504
rect 20254 16464 20260 16476
rect 20312 16464 20318 16516
rect 20349 16507 20407 16513
rect 20349 16473 20361 16507
rect 20395 16504 20407 16507
rect 20714 16504 20720 16516
rect 20395 16476 20720 16504
rect 20395 16473 20407 16476
rect 20349 16467 20407 16473
rect 20714 16464 20720 16476
rect 20772 16464 20778 16516
rect 21358 16464 21364 16516
rect 21416 16504 21422 16516
rect 22204 16504 22232 16544
rect 22646 16504 22652 16516
rect 21416 16476 22094 16504
rect 22204 16476 22652 16504
rect 21416 16464 21422 16476
rect 20622 16436 20628 16448
rect 18892 16408 20628 16436
rect 17736 16396 17742 16408
rect 20622 16396 20628 16408
rect 20680 16396 20686 16448
rect 20806 16396 20812 16448
rect 20864 16436 20870 16448
rect 21453 16439 21511 16445
rect 21453 16436 21465 16439
rect 20864 16408 21465 16436
rect 20864 16396 20870 16408
rect 21453 16405 21465 16408
rect 21499 16405 21511 16439
rect 22066 16436 22094 16476
rect 22646 16464 22652 16476
rect 22704 16464 22710 16516
rect 22741 16507 22799 16513
rect 22741 16473 22753 16507
rect 22787 16473 22799 16507
rect 22741 16467 22799 16473
rect 22833 16507 22891 16513
rect 22833 16473 22845 16507
rect 22879 16504 22891 16507
rect 23014 16504 23020 16516
rect 22879 16476 23020 16504
rect 22879 16473 22891 16476
rect 22833 16467 22891 16473
rect 22756 16436 22784 16467
rect 23014 16464 23020 16476
rect 23072 16504 23078 16516
rect 23492 16504 23520 16612
rect 24854 16600 24860 16612
rect 24912 16640 24918 16652
rect 25038 16640 25044 16652
rect 24912 16612 25044 16640
rect 24912 16600 24918 16612
rect 25038 16600 25044 16612
rect 25096 16600 25102 16652
rect 25240 16649 25268 16680
rect 25774 16668 25780 16680
rect 25832 16708 25838 16720
rect 27172 16708 27200 16748
rect 28261 16711 28319 16717
rect 28261 16708 28273 16711
rect 25832 16680 26464 16708
rect 25832 16668 25838 16680
rect 26436 16652 26464 16680
rect 27172 16680 28273 16708
rect 25225 16643 25283 16649
rect 25225 16609 25237 16643
rect 25271 16609 25283 16643
rect 26050 16640 26056 16652
rect 26011 16612 26056 16640
rect 25225 16603 25283 16609
rect 26050 16600 26056 16612
rect 26108 16600 26114 16652
rect 26418 16640 26424 16652
rect 26379 16612 26424 16640
rect 26418 16600 26424 16612
rect 26476 16600 26482 16652
rect 26786 16532 26792 16584
rect 26844 16572 26850 16584
rect 27172 16581 27200 16680
rect 28261 16677 28273 16680
rect 28307 16677 28319 16711
rect 28261 16671 28319 16677
rect 27338 16600 27344 16652
rect 27396 16640 27402 16652
rect 27396 16612 27660 16640
rect 27396 16600 27402 16612
rect 27632 16581 27660 16612
rect 27065 16575 27123 16581
rect 27065 16572 27077 16575
rect 26844 16544 27077 16572
rect 26844 16532 26850 16544
rect 27065 16541 27077 16544
rect 27111 16541 27123 16575
rect 27065 16535 27123 16541
rect 27157 16575 27215 16581
rect 27157 16541 27169 16575
rect 27203 16541 27215 16575
rect 27157 16535 27215 16541
rect 27617 16575 27675 16581
rect 27617 16541 27629 16575
rect 27663 16541 27675 16575
rect 27617 16535 27675 16541
rect 24578 16504 24584 16516
rect 23072 16476 23520 16504
rect 24539 16476 24584 16504
rect 23072 16464 23078 16476
rect 24578 16464 24584 16476
rect 24636 16464 24642 16516
rect 25133 16507 25191 16513
rect 25133 16473 25145 16507
rect 25179 16473 25191 16507
rect 26326 16504 26332 16516
rect 26287 16476 26332 16504
rect 25133 16467 25191 16473
rect 23382 16436 23388 16448
rect 22066 16408 22784 16436
rect 23343 16408 23388 16436
rect 21453 16399 21511 16405
rect 23382 16396 23388 16408
rect 23440 16396 23446 16448
rect 25148 16436 25176 16467
rect 26326 16464 26332 16476
rect 26384 16464 26390 16516
rect 26418 16464 26424 16516
rect 26476 16504 26482 16516
rect 30282 16504 30288 16516
rect 26476 16476 30288 16504
rect 26476 16464 26482 16476
rect 30282 16464 30288 16476
rect 30340 16464 30346 16516
rect 26142 16436 26148 16448
rect 25148 16408 26148 16436
rect 26142 16396 26148 16408
rect 26200 16396 26206 16448
rect 26602 16396 26608 16448
rect 26660 16436 26666 16448
rect 27709 16439 27767 16445
rect 27709 16436 27721 16439
rect 26660 16408 27721 16436
rect 26660 16396 26666 16408
rect 27709 16405 27721 16408
rect 27755 16405 27767 16439
rect 27709 16399 27767 16405
rect 28442 16396 28448 16448
rect 28500 16436 28506 16448
rect 28813 16439 28871 16445
rect 28813 16436 28825 16439
rect 28500 16408 28825 16436
rect 28500 16396 28506 16408
rect 28813 16405 28825 16408
rect 28859 16405 28871 16439
rect 28813 16399 28871 16405
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 11054 16192 11060 16244
rect 11112 16232 11118 16244
rect 17310 16232 17316 16244
rect 11112 16204 14228 16232
rect 11112 16192 11118 16204
rect 12986 16164 12992 16176
rect 12947 16136 12992 16164
rect 12986 16124 12992 16136
rect 13044 16124 13050 16176
rect 14200 16173 14228 16204
rect 14752 16204 17316 16232
rect 14752 16173 14780 16204
rect 17310 16192 17316 16204
rect 17368 16192 17374 16244
rect 18322 16232 18328 16244
rect 18283 16204 18328 16232
rect 18322 16192 18328 16204
rect 18380 16192 18386 16244
rect 21542 16232 21548 16244
rect 18432 16204 21548 16232
rect 14185 16167 14243 16173
rect 14185 16133 14197 16167
rect 14231 16133 14243 16167
rect 14185 16127 14243 16133
rect 14737 16167 14795 16173
rect 14737 16133 14749 16167
rect 14783 16133 14795 16167
rect 15746 16164 15752 16176
rect 15707 16136 15752 16164
rect 14737 16127 14795 16133
rect 15746 16124 15752 16136
rect 15804 16124 15810 16176
rect 16390 16124 16396 16176
rect 16448 16164 16454 16176
rect 17037 16167 17095 16173
rect 17037 16164 17049 16167
rect 16448 16136 17049 16164
rect 16448 16124 16454 16136
rect 17037 16133 17049 16136
rect 17083 16133 17095 16167
rect 17037 16127 17095 16133
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16096 1915 16099
rect 8110 16096 8116 16108
rect 1903 16068 8116 16096
rect 1903 16065 1915 16068
rect 1857 16059 1915 16065
rect 8110 16056 8116 16068
rect 8168 16056 8174 16108
rect 11146 16096 11152 16108
rect 11059 16068 11152 16096
rect 11146 16056 11152 16068
rect 11204 16096 11210 16108
rect 18432 16105 18460 16204
rect 21542 16192 21548 16204
rect 21600 16192 21606 16244
rect 22186 16232 22192 16244
rect 22066 16204 22192 16232
rect 19613 16167 19671 16173
rect 19613 16133 19625 16167
rect 19659 16164 19671 16167
rect 20346 16164 20352 16176
rect 19659 16136 20352 16164
rect 19659 16133 19671 16136
rect 19613 16127 19671 16133
rect 20346 16124 20352 16136
rect 20404 16124 20410 16176
rect 20901 16167 20959 16173
rect 20901 16133 20913 16167
rect 20947 16164 20959 16167
rect 22066 16164 22094 16204
rect 22186 16192 22192 16204
rect 22244 16192 22250 16244
rect 26234 16232 26240 16244
rect 24504 16204 26240 16232
rect 24504 16176 24532 16204
rect 26234 16192 26240 16204
rect 26292 16192 26298 16244
rect 26326 16192 26332 16244
rect 26384 16232 26390 16244
rect 26421 16235 26479 16241
rect 26421 16232 26433 16235
rect 26384 16204 26433 16232
rect 26384 16192 26390 16204
rect 26421 16201 26433 16204
rect 26467 16201 26479 16235
rect 26421 16195 26479 16201
rect 28629 16235 28687 16241
rect 28629 16201 28641 16235
rect 28675 16232 28687 16235
rect 28675 16204 35894 16232
rect 28675 16201 28687 16204
rect 28629 16195 28687 16201
rect 23566 16164 23572 16176
rect 20947 16136 22094 16164
rect 22204 16136 23572 16164
rect 20947 16133 20959 16136
rect 20901 16127 20959 16133
rect 12161 16099 12219 16105
rect 12161 16096 12173 16099
rect 11204 16068 12173 16096
rect 11204 16056 11210 16068
rect 12161 16065 12173 16068
rect 12207 16065 12219 16099
rect 12161 16059 12219 16065
rect 18417 16099 18475 16105
rect 18417 16065 18429 16099
rect 18463 16065 18475 16099
rect 19058 16096 19064 16108
rect 18417 16059 18475 16065
rect 18524 16068 19064 16096
rect 12894 16028 12900 16040
rect 12855 16000 12900 16028
rect 12894 15988 12900 16000
rect 12952 15988 12958 16040
rect 14093 16031 14151 16037
rect 13280 16000 14044 16028
rect 9766 15920 9772 15972
rect 9824 15960 9830 15972
rect 10137 15963 10195 15969
rect 10137 15960 10149 15963
rect 9824 15932 10149 15960
rect 9824 15920 9830 15932
rect 10137 15929 10149 15932
rect 10183 15960 10195 15963
rect 12526 15960 12532 15972
rect 10183 15932 12532 15960
rect 10183 15929 10195 15932
rect 10137 15923 10195 15929
rect 12526 15920 12532 15932
rect 12584 15920 12590 15972
rect 12618 15920 12624 15972
rect 12676 15960 12682 15972
rect 13280 15960 13308 16000
rect 12676 15932 13308 15960
rect 13449 15963 13507 15969
rect 12676 15920 12682 15932
rect 13449 15929 13461 15963
rect 13495 15960 13507 15963
rect 13538 15960 13544 15972
rect 13495 15932 13544 15960
rect 13495 15929 13507 15932
rect 13449 15923 13507 15929
rect 13538 15920 13544 15932
rect 13596 15920 13602 15972
rect 14016 15960 14044 16000
rect 14093 15997 14105 16031
rect 14139 16028 14151 16031
rect 14366 16028 14372 16040
rect 14139 16000 14372 16028
rect 14139 15997 14151 16000
rect 14093 15991 14151 15997
rect 14366 15988 14372 16000
rect 14424 16028 14430 16040
rect 15102 16028 15108 16040
rect 14424 16000 15108 16028
rect 14424 15988 14430 16000
rect 15102 15988 15108 16000
rect 15160 15988 15166 16040
rect 15657 16031 15715 16037
rect 15657 15997 15669 16031
rect 15703 16016 15715 16031
rect 16758 16028 16764 16040
rect 15764 16016 16764 16028
rect 15703 16000 16764 16016
rect 15703 15997 15792 16000
rect 15657 15991 15792 15997
rect 15672 15988 15792 15991
rect 16758 15988 16764 16000
rect 16816 15988 16822 16040
rect 16942 16028 16948 16040
rect 16903 16000 16948 16028
rect 16942 15988 16948 16000
rect 17000 15988 17006 16040
rect 18524 16028 18552 16068
rect 19058 16056 19064 16068
rect 19116 16056 19122 16108
rect 22002 16096 22008 16108
rect 21963 16068 22008 16096
rect 22002 16056 22008 16068
rect 22060 16056 22066 16108
rect 22204 16105 22232 16136
rect 23566 16124 23572 16136
rect 23624 16124 23630 16176
rect 23753 16167 23811 16173
rect 23753 16133 23765 16167
rect 23799 16164 23811 16167
rect 24026 16164 24032 16176
rect 23799 16136 24032 16164
rect 23799 16133 23811 16136
rect 23753 16127 23811 16133
rect 24026 16124 24032 16136
rect 24084 16124 24090 16176
rect 24486 16164 24492 16176
rect 24447 16136 24492 16164
rect 24486 16124 24492 16136
rect 24544 16124 24550 16176
rect 25685 16167 25743 16173
rect 25685 16133 25697 16167
rect 25731 16164 25743 16167
rect 27893 16167 27951 16173
rect 27893 16164 27905 16167
rect 25731 16136 27905 16164
rect 25731 16133 25743 16136
rect 25685 16127 25743 16133
rect 27893 16133 27905 16136
rect 27939 16133 27951 16167
rect 29089 16167 29147 16173
rect 29089 16164 29101 16167
rect 27893 16127 27951 16133
rect 28000 16136 29101 16164
rect 28000 16108 28028 16136
rect 29089 16133 29101 16136
rect 29135 16133 29147 16167
rect 35866 16164 35894 16204
rect 38010 16164 38016 16176
rect 35866 16136 38016 16164
rect 29089 16127 29147 16133
rect 38010 16124 38016 16136
rect 38068 16124 38074 16176
rect 22189 16099 22247 16105
rect 22189 16065 22201 16099
rect 22235 16065 22247 16099
rect 22189 16059 22247 16065
rect 24673 16099 24731 16105
rect 24673 16065 24685 16099
rect 24719 16096 24731 16099
rect 26329 16099 26387 16105
rect 24719 16068 25176 16096
rect 24719 16065 24731 16068
rect 24673 16059 24731 16065
rect 17420 16000 18552 16028
rect 15562 15960 15568 15972
rect 14016 15932 15568 15960
rect 15562 15920 15568 15932
rect 15620 15920 15626 15972
rect 15764 15960 15792 15988
rect 15672 15932 15792 15960
rect 16209 15963 16267 15969
rect 1670 15892 1676 15904
rect 1631 15864 1676 15892
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 12253 15895 12311 15901
rect 12253 15861 12265 15895
rect 12299 15892 12311 15895
rect 15672 15892 15700 15932
rect 16209 15929 16221 15963
rect 16255 15960 16267 15963
rect 17420 15960 17448 16000
rect 18782 15988 18788 16040
rect 18840 16028 18846 16040
rect 19705 16031 19763 16037
rect 19705 16028 19717 16031
rect 18840 16000 19717 16028
rect 18840 15988 18846 16000
rect 19705 15997 19717 16000
rect 19751 16028 19763 16031
rect 20993 16031 21051 16037
rect 20993 16028 21005 16031
rect 19751 16000 21005 16028
rect 19751 15997 19763 16000
rect 19705 15991 19763 15997
rect 20993 15997 21005 16000
rect 21039 15997 21051 16031
rect 23198 16028 23204 16040
rect 23159 16000 23204 16028
rect 20993 15991 21051 15997
rect 23198 15988 23204 16000
rect 23256 15988 23262 16040
rect 23750 16028 23756 16040
rect 23308 16000 23756 16028
rect 16255 15932 17448 15960
rect 17497 15963 17555 15969
rect 16255 15929 16267 15932
rect 16209 15923 16267 15929
rect 17497 15929 17509 15963
rect 17543 15960 17555 15963
rect 17954 15960 17960 15972
rect 17543 15932 17960 15960
rect 17543 15929 17555 15932
rect 17497 15923 17555 15929
rect 17954 15920 17960 15932
rect 18012 15960 18018 15972
rect 19150 15960 19156 15972
rect 18012 15932 19156 15960
rect 18012 15920 18018 15932
rect 19150 15920 19156 15932
rect 19208 15920 19214 15972
rect 20438 15960 20444 15972
rect 20399 15932 20444 15960
rect 20438 15920 20444 15932
rect 20496 15920 20502 15972
rect 20622 15920 20628 15972
rect 20680 15960 20686 15972
rect 22094 15960 22100 15972
rect 20680 15932 22100 15960
rect 20680 15920 20686 15932
rect 22094 15920 22100 15932
rect 22152 15920 22158 15972
rect 23308 15960 23336 16000
rect 23750 15988 23756 16000
rect 23808 15988 23814 16040
rect 23845 16031 23903 16037
rect 23845 15997 23857 16031
rect 23891 16028 23903 16031
rect 24762 16028 24768 16040
rect 23891 16000 24768 16028
rect 23891 15997 23903 16000
rect 23845 15991 23903 15997
rect 24762 15988 24768 16000
rect 24820 15988 24826 16040
rect 25148 16028 25176 16068
rect 26329 16065 26341 16099
rect 26375 16096 26387 16099
rect 26510 16096 26516 16108
rect 26375 16068 26516 16096
rect 26375 16065 26387 16068
rect 26329 16059 26387 16065
rect 26510 16056 26516 16068
rect 26568 16056 26574 16108
rect 26786 16096 26792 16108
rect 26620 16068 26792 16096
rect 25774 16028 25780 16040
rect 25148 16000 25636 16028
rect 25735 16000 25780 16028
rect 22388 15932 23336 15960
rect 12299 15864 15700 15892
rect 12299 15861 12311 15864
rect 12253 15855 12311 15861
rect 15746 15852 15752 15904
rect 15804 15892 15810 15904
rect 18138 15892 18144 15904
rect 15804 15864 18144 15892
rect 15804 15852 15810 15864
rect 18138 15852 18144 15864
rect 18196 15852 18202 15904
rect 20070 15852 20076 15904
rect 20128 15892 20134 15904
rect 22388 15892 22416 15932
rect 23474 15920 23480 15972
rect 23532 15960 23538 15972
rect 25225 15963 25283 15969
rect 25225 15960 25237 15963
rect 23532 15932 25237 15960
rect 23532 15920 23538 15932
rect 25225 15929 25237 15932
rect 25271 15960 25283 15963
rect 25498 15960 25504 15972
rect 25271 15932 25504 15960
rect 25271 15929 25283 15932
rect 25225 15923 25283 15929
rect 25498 15920 25504 15932
rect 25556 15920 25562 15972
rect 25608 15960 25636 16000
rect 25774 15988 25780 16000
rect 25832 15988 25838 16040
rect 25958 15988 25964 16040
rect 26016 16028 26022 16040
rect 26620 16028 26648 16068
rect 26786 16056 26792 16068
rect 26844 16056 26850 16108
rect 27154 16096 27160 16108
rect 27115 16068 27160 16096
rect 27154 16056 27160 16068
rect 27212 16056 27218 16108
rect 27982 16096 27988 16108
rect 27943 16068 27988 16096
rect 27982 16056 27988 16068
rect 28040 16056 28046 16108
rect 28442 16096 28448 16108
rect 28403 16068 28448 16096
rect 28442 16056 28448 16068
rect 28500 16056 28506 16108
rect 37553 16099 37611 16105
rect 37553 16065 37565 16099
rect 37599 16096 37611 16099
rect 38194 16096 38200 16108
rect 37599 16068 38200 16096
rect 37599 16065 37611 16068
rect 37553 16059 37611 16065
rect 38194 16056 38200 16068
rect 38252 16056 38258 16108
rect 26016 16000 26648 16028
rect 26016 15988 26022 16000
rect 30190 15960 30196 15972
rect 25608 15932 30196 15960
rect 30190 15920 30196 15932
rect 30248 15920 30254 15972
rect 38010 15960 38016 15972
rect 37971 15932 38016 15960
rect 38010 15920 38016 15932
rect 38068 15920 38074 15972
rect 20128 15864 22416 15892
rect 20128 15852 20134 15864
rect 23198 15852 23204 15904
rect 23256 15892 23262 15904
rect 23658 15892 23664 15904
rect 23256 15864 23664 15892
rect 23256 15852 23262 15864
rect 23658 15852 23664 15864
rect 23716 15852 23722 15904
rect 26326 15852 26332 15904
rect 26384 15892 26390 15904
rect 27249 15895 27307 15901
rect 27249 15892 27261 15895
rect 26384 15864 27261 15892
rect 26384 15852 26390 15864
rect 27249 15861 27261 15864
rect 27295 15861 27307 15895
rect 27249 15855 27307 15861
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 8110 15688 8116 15700
rect 8071 15660 8116 15688
rect 8110 15648 8116 15660
rect 8168 15648 8174 15700
rect 9674 15688 9680 15700
rect 9635 15660 9680 15688
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 12529 15691 12587 15697
rect 12529 15657 12541 15691
rect 12575 15688 12587 15691
rect 14458 15688 14464 15700
rect 12575 15660 14464 15688
rect 12575 15657 12587 15660
rect 12529 15651 12587 15657
rect 14458 15648 14464 15660
rect 14516 15648 14522 15700
rect 15102 15648 15108 15700
rect 15160 15688 15166 15700
rect 17862 15688 17868 15700
rect 15160 15660 17868 15688
rect 15160 15648 15166 15660
rect 17862 15648 17868 15660
rect 17920 15648 17926 15700
rect 18782 15688 18788 15700
rect 18743 15660 18788 15688
rect 18782 15648 18788 15660
rect 18840 15648 18846 15700
rect 20530 15688 20536 15700
rect 19628 15660 20536 15688
rect 14274 15580 14280 15632
rect 14332 15580 14338 15632
rect 15562 15580 15568 15632
rect 15620 15620 15626 15632
rect 15841 15623 15899 15629
rect 15841 15620 15853 15623
rect 15620 15592 15853 15620
rect 15620 15580 15626 15592
rect 15841 15589 15853 15592
rect 15887 15620 15899 15623
rect 16942 15620 16948 15632
rect 15887 15592 16948 15620
rect 15887 15589 15899 15592
rect 15841 15583 15899 15589
rect 16942 15580 16948 15592
rect 17000 15620 17006 15632
rect 17037 15623 17095 15629
rect 17037 15620 17049 15623
rect 17000 15592 17049 15620
rect 17000 15580 17006 15592
rect 17037 15589 17049 15592
rect 17083 15589 17095 15623
rect 17037 15583 17095 15589
rect 17218 15580 17224 15632
rect 17276 15620 17282 15632
rect 19518 15620 19524 15632
rect 17276 15592 19524 15620
rect 17276 15580 17282 15592
rect 19518 15580 19524 15592
rect 19576 15580 19582 15632
rect 10962 15512 10968 15564
rect 11020 15552 11026 15564
rect 11885 15555 11943 15561
rect 11020 15524 11836 15552
rect 11020 15512 11026 15524
rect 8202 15484 8208 15496
rect 8163 15456 8208 15484
rect 8202 15444 8208 15456
rect 8260 15444 8266 15496
rect 9674 15444 9680 15496
rect 9732 15484 9738 15496
rect 10229 15487 10287 15493
rect 10229 15484 10241 15487
rect 9732 15456 10241 15484
rect 9732 15444 9738 15456
rect 10229 15453 10241 15456
rect 10275 15453 10287 15487
rect 11146 15484 11152 15496
rect 11107 15456 11152 15484
rect 10229 15447 10287 15453
rect 11146 15444 11152 15456
rect 11204 15444 11210 15496
rect 11808 15493 11836 15524
rect 11885 15521 11897 15555
rect 11931 15552 11943 15555
rect 13265 15555 13323 15561
rect 13265 15552 13277 15555
rect 11931 15524 13277 15552
rect 11931 15521 11943 15524
rect 11885 15515 11943 15521
rect 13265 15521 13277 15524
rect 13311 15521 13323 15555
rect 14292 15552 14320 15580
rect 14369 15555 14427 15561
rect 14369 15552 14381 15555
rect 14292 15524 14381 15552
rect 13265 15515 13323 15521
rect 14369 15521 14381 15524
rect 14415 15521 14427 15555
rect 19628 15552 19656 15660
rect 20530 15648 20536 15660
rect 20588 15648 20594 15700
rect 23934 15648 23940 15700
rect 23992 15688 23998 15700
rect 27430 15688 27436 15700
rect 23992 15660 27436 15688
rect 23992 15648 23998 15660
rect 27430 15648 27436 15660
rect 27488 15648 27494 15700
rect 30929 15691 30987 15697
rect 30929 15657 30941 15691
rect 30975 15688 30987 15691
rect 36630 15688 36636 15700
rect 30975 15660 36636 15688
rect 30975 15657 30987 15660
rect 30929 15651 30987 15657
rect 36630 15648 36636 15660
rect 36688 15648 36694 15700
rect 19978 15580 19984 15632
rect 20036 15620 20042 15632
rect 20438 15620 20444 15632
rect 20036 15592 20444 15620
rect 20036 15580 20042 15592
rect 20438 15580 20444 15592
rect 20496 15580 20502 15632
rect 20548 15620 20576 15648
rect 24578 15620 24584 15632
rect 20548 15592 24584 15620
rect 24578 15580 24584 15592
rect 24636 15620 24642 15632
rect 24673 15623 24731 15629
rect 24673 15620 24685 15623
rect 24636 15592 24685 15620
rect 24636 15580 24642 15592
rect 24673 15589 24685 15592
rect 24719 15589 24731 15623
rect 24673 15583 24731 15589
rect 25148 15592 27200 15620
rect 14369 15515 14427 15521
rect 16960 15524 19656 15552
rect 19705 15555 19763 15561
rect 11793 15487 11851 15493
rect 11793 15453 11805 15487
rect 11839 15453 11851 15487
rect 11793 15447 11851 15453
rect 12437 15487 12495 15493
rect 12437 15453 12449 15487
rect 12483 15484 12495 15487
rect 12710 15484 12716 15496
rect 12483 15456 12716 15484
rect 12483 15453 12495 15456
rect 12437 15447 12495 15453
rect 12710 15444 12716 15456
rect 12768 15444 12774 15496
rect 12894 15444 12900 15496
rect 12952 15484 12958 15496
rect 13081 15487 13139 15493
rect 13081 15484 13093 15487
rect 12952 15456 13093 15484
rect 12952 15444 12958 15456
rect 13081 15453 13093 15456
rect 13127 15453 13139 15487
rect 13081 15447 13139 15453
rect 10321 15419 10379 15425
rect 10321 15385 10333 15419
rect 10367 15416 10379 15419
rect 14461 15419 14519 15425
rect 10367 15388 14412 15416
rect 10367 15385 10379 15388
rect 10321 15379 10379 15385
rect 11241 15351 11299 15357
rect 11241 15317 11253 15351
rect 11287 15348 11299 15351
rect 11790 15348 11796 15360
rect 11287 15320 11796 15348
rect 11287 15317 11299 15320
rect 11241 15311 11299 15317
rect 11790 15308 11796 15320
rect 11848 15348 11854 15360
rect 12434 15348 12440 15360
rect 11848 15320 12440 15348
rect 11848 15308 11854 15320
rect 12434 15308 12440 15320
rect 12492 15308 12498 15360
rect 13630 15308 13636 15360
rect 13688 15348 13694 15360
rect 13725 15351 13783 15357
rect 13725 15348 13737 15351
rect 13688 15320 13737 15348
rect 13688 15308 13694 15320
rect 13725 15317 13737 15320
rect 13771 15317 13783 15351
rect 14384 15348 14412 15388
rect 14461 15385 14473 15419
rect 14507 15416 14519 15419
rect 14550 15416 14556 15428
rect 14507 15388 14556 15416
rect 14507 15385 14519 15388
rect 14461 15379 14519 15385
rect 14550 15376 14556 15388
rect 14608 15376 14614 15428
rect 15013 15419 15071 15425
rect 15013 15385 15025 15419
rect 15059 15416 15071 15419
rect 15102 15416 15108 15428
rect 15059 15388 15108 15416
rect 15059 15385 15071 15388
rect 15013 15379 15071 15385
rect 15102 15376 15108 15388
rect 15160 15376 15166 15428
rect 16298 15416 16304 15428
rect 16259 15388 16304 15416
rect 16298 15376 16304 15388
rect 16356 15376 16362 15428
rect 16393 15419 16451 15425
rect 16393 15385 16405 15419
rect 16439 15416 16451 15419
rect 16960 15416 16988 15524
rect 19705 15521 19717 15555
rect 19751 15552 19763 15555
rect 20254 15552 20260 15564
rect 19751 15524 20260 15552
rect 19751 15521 19763 15524
rect 19705 15515 19763 15521
rect 20254 15512 20260 15524
rect 20312 15512 20318 15564
rect 23106 15552 23112 15564
rect 23067 15524 23112 15552
rect 23106 15512 23112 15524
rect 23164 15512 23170 15564
rect 23382 15552 23388 15564
rect 23343 15524 23388 15552
rect 23382 15512 23388 15524
rect 23440 15512 23446 15564
rect 23566 15512 23572 15564
rect 23624 15552 23630 15564
rect 25148 15552 25176 15592
rect 23624 15524 25176 15552
rect 25225 15555 25283 15561
rect 23624 15512 23630 15524
rect 25225 15521 25237 15555
rect 25271 15552 25283 15555
rect 26970 15552 26976 15564
rect 25271 15524 26976 15552
rect 25271 15521 25283 15524
rect 25225 15515 25283 15521
rect 26970 15512 26976 15524
rect 27028 15512 27034 15564
rect 27172 15552 27200 15592
rect 28534 15552 28540 15564
rect 27172 15524 28540 15552
rect 18506 15444 18512 15496
rect 18564 15484 18570 15496
rect 18693 15487 18751 15493
rect 18693 15484 18705 15487
rect 18564 15456 18705 15484
rect 18564 15444 18570 15456
rect 18693 15453 18705 15456
rect 18739 15484 18751 15487
rect 19886 15484 19892 15496
rect 18739 15456 19892 15484
rect 18739 15453 18751 15456
rect 18693 15447 18751 15453
rect 19886 15444 19892 15456
rect 19944 15444 19950 15496
rect 20349 15487 20407 15493
rect 20349 15453 20361 15487
rect 20395 15484 20407 15487
rect 20530 15484 20536 15496
rect 20395 15456 20536 15484
rect 20395 15453 20407 15456
rect 20349 15447 20407 15453
rect 20530 15444 20536 15456
rect 20588 15444 20594 15496
rect 21910 15444 21916 15496
rect 21968 15484 21974 15496
rect 22373 15487 22431 15493
rect 22373 15484 22385 15487
rect 21968 15456 22385 15484
rect 21968 15444 21974 15456
rect 22373 15453 22385 15456
rect 22419 15484 22431 15487
rect 22922 15484 22928 15496
rect 22419 15456 22928 15484
rect 22419 15453 22431 15456
rect 22373 15447 22431 15453
rect 22922 15444 22928 15456
rect 22980 15444 22986 15496
rect 25498 15444 25504 15496
rect 25556 15484 25562 15496
rect 27172 15493 27200 15524
rect 28534 15512 28540 15524
rect 28592 15512 28598 15564
rect 25777 15487 25835 15493
rect 25777 15484 25789 15487
rect 25556 15456 25789 15484
rect 25556 15444 25562 15456
rect 25777 15453 25789 15456
rect 25823 15453 25835 15487
rect 25777 15447 25835 15453
rect 27157 15487 27215 15493
rect 27157 15453 27169 15487
rect 27203 15453 27215 15487
rect 27157 15447 27215 15453
rect 27246 15444 27252 15496
rect 27304 15484 27310 15496
rect 27617 15487 27675 15493
rect 27617 15484 27629 15487
rect 27304 15456 27629 15484
rect 27304 15444 27310 15456
rect 27617 15453 27629 15456
rect 27663 15453 27675 15487
rect 27617 15447 27675 15453
rect 28445 15487 28503 15493
rect 28445 15453 28457 15487
rect 28491 15484 28503 15487
rect 28994 15484 29000 15496
rect 28491 15456 29000 15484
rect 28491 15453 28503 15456
rect 28445 15447 28503 15453
rect 28994 15444 29000 15456
rect 29052 15484 29058 15496
rect 29733 15487 29791 15493
rect 29733 15484 29745 15487
rect 29052 15456 29745 15484
rect 29052 15444 29058 15456
rect 29733 15453 29745 15456
rect 29779 15453 29791 15487
rect 29733 15447 29791 15453
rect 30837 15487 30895 15493
rect 30837 15453 30849 15487
rect 30883 15453 30895 15487
rect 30837 15447 30895 15453
rect 17494 15416 17500 15428
rect 16439 15388 16988 15416
rect 17455 15388 17500 15416
rect 16439 15385 16451 15388
rect 16393 15379 16451 15385
rect 17494 15376 17500 15388
rect 17552 15376 17558 15428
rect 17589 15419 17647 15425
rect 17589 15385 17601 15419
rect 17635 15416 17647 15419
rect 17954 15416 17960 15428
rect 17635 15388 17960 15416
rect 17635 15385 17647 15388
rect 17589 15379 17647 15385
rect 17954 15376 17960 15388
rect 18012 15376 18018 15428
rect 20070 15416 20076 15428
rect 18064 15388 20076 15416
rect 16850 15348 16856 15360
rect 14384 15320 16856 15348
rect 13725 15311 13783 15317
rect 16850 15308 16856 15320
rect 16908 15308 16914 15360
rect 17402 15308 17408 15360
rect 17460 15348 17466 15360
rect 18064 15348 18092 15388
rect 20070 15376 20076 15388
rect 20128 15376 20134 15428
rect 20438 15376 20444 15428
rect 20496 15416 20502 15428
rect 20901 15419 20959 15425
rect 20901 15416 20913 15419
rect 20496 15388 20913 15416
rect 20496 15376 20502 15388
rect 20901 15385 20913 15388
rect 20947 15385 20959 15419
rect 20901 15379 20959 15385
rect 20990 15376 20996 15428
rect 21048 15416 21054 15428
rect 21542 15416 21548 15428
rect 21048 15388 21093 15416
rect 21503 15388 21548 15416
rect 21048 15376 21054 15388
rect 21542 15376 21548 15388
rect 21600 15376 21606 15428
rect 23201 15419 23259 15425
rect 23201 15385 23213 15419
rect 23247 15416 23259 15419
rect 24946 15416 24952 15428
rect 23247 15388 23704 15416
rect 23247 15385 23259 15388
rect 23201 15379 23259 15385
rect 17460 15320 18092 15348
rect 17460 15308 17466 15320
rect 18138 15308 18144 15360
rect 18196 15348 18202 15360
rect 20254 15348 20260 15360
rect 18196 15320 18241 15348
rect 20215 15320 20260 15348
rect 18196 15308 18202 15320
rect 20254 15308 20260 15320
rect 20312 15308 20318 15360
rect 22465 15351 22523 15357
rect 22465 15317 22477 15351
rect 22511 15348 22523 15351
rect 22922 15348 22928 15360
rect 22511 15320 22928 15348
rect 22511 15317 22523 15320
rect 22465 15311 22523 15317
rect 22922 15308 22928 15320
rect 22980 15308 22986 15360
rect 23676 15348 23704 15388
rect 24688 15388 24952 15416
rect 24688 15348 24716 15388
rect 24946 15376 24952 15388
rect 25004 15376 25010 15428
rect 25130 15416 25136 15428
rect 25091 15388 25136 15416
rect 25130 15376 25136 15388
rect 25188 15376 25194 15428
rect 26326 15416 26332 15428
rect 26287 15388 26332 15416
rect 26326 15376 26332 15388
rect 26384 15376 26390 15428
rect 26418 15376 26424 15428
rect 26476 15416 26482 15428
rect 26476 15388 26521 15416
rect 26476 15376 26482 15388
rect 26786 15376 26792 15428
rect 26844 15416 26850 15428
rect 30852 15416 30880 15447
rect 26844 15388 30880 15416
rect 26844 15376 26850 15388
rect 23676 15320 24716 15348
rect 24762 15308 24768 15360
rect 24820 15348 24826 15360
rect 27065 15351 27123 15357
rect 27065 15348 27077 15351
rect 24820 15320 27077 15348
rect 24820 15308 24826 15320
rect 27065 15317 27077 15320
rect 27111 15317 27123 15351
rect 27706 15348 27712 15360
rect 27667 15320 27712 15348
rect 27065 15311 27123 15317
rect 27706 15308 27712 15320
rect 27764 15308 27770 15360
rect 28166 15308 28172 15360
rect 28224 15348 28230 15360
rect 28353 15351 28411 15357
rect 28353 15348 28365 15351
rect 28224 15320 28365 15348
rect 28224 15308 28230 15320
rect 28353 15317 28365 15320
rect 28399 15317 28411 15351
rect 28353 15311 28411 15317
rect 28534 15308 28540 15360
rect 28592 15348 28598 15360
rect 28997 15351 29055 15357
rect 28997 15348 29009 15351
rect 28592 15320 29009 15348
rect 28592 15308 28598 15320
rect 28997 15317 29009 15320
rect 29043 15348 29055 15351
rect 30926 15348 30932 15360
rect 29043 15320 30932 15348
rect 29043 15317 29055 15320
rect 28997 15311 29055 15317
rect 30926 15308 30932 15320
rect 30984 15308 30990 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 11054 15144 11060 15156
rect 11015 15116 11060 15144
rect 11054 15104 11060 15116
rect 11112 15104 11118 15156
rect 15010 15104 15016 15156
rect 15068 15144 15074 15156
rect 17954 15144 17960 15156
rect 15068 15116 17960 15144
rect 15068 15104 15074 15116
rect 17954 15104 17960 15116
rect 18012 15104 18018 15156
rect 20346 15144 20352 15156
rect 18432 15116 20024 15144
rect 20307 15116 20352 15144
rect 9861 15079 9919 15085
rect 9861 15045 9873 15079
rect 9907 15076 9919 15079
rect 12989 15079 13047 15085
rect 12989 15076 13001 15079
rect 9907 15048 12204 15076
rect 9907 15045 9919 15048
rect 9861 15039 9919 15045
rect 12176 15020 12204 15048
rect 12268 15048 13001 15076
rect 9309 15011 9367 15017
rect 9309 14977 9321 15011
rect 9355 15008 9367 15011
rect 10226 15008 10232 15020
rect 9355 14980 10232 15008
rect 9355 14977 9367 14980
rect 9309 14971 9367 14977
rect 10226 14968 10232 14980
rect 10284 15008 10290 15020
rect 10321 15011 10379 15017
rect 10321 15008 10333 15011
rect 10284 14980 10333 15008
rect 10284 14968 10290 14980
rect 10321 14977 10333 14980
rect 10367 14977 10379 15011
rect 10321 14971 10379 14977
rect 10410 14968 10416 15020
rect 10468 15008 10474 15020
rect 10962 15008 10968 15020
rect 10468 14980 10968 15008
rect 10468 14968 10474 14980
rect 10962 14968 10968 14980
rect 11020 14968 11026 15020
rect 12158 15008 12164 15020
rect 12071 14980 12164 15008
rect 12158 14968 12164 14980
rect 12216 14968 12222 15020
rect 12268 14940 12296 15048
rect 12989 15045 13001 15048
rect 13035 15045 13047 15079
rect 12989 15039 13047 15045
rect 13078 15036 13084 15088
rect 13136 15076 13142 15088
rect 13538 15076 13544 15088
rect 13136 15048 13544 15076
rect 13136 15036 13142 15048
rect 13538 15036 13544 15048
rect 13596 15036 13602 15088
rect 14182 15076 14188 15088
rect 14143 15048 14188 15076
rect 14182 15036 14188 15048
rect 14240 15036 14246 15088
rect 15378 15076 15384 15088
rect 15339 15048 15384 15076
rect 15378 15036 15384 15048
rect 15436 15036 15442 15088
rect 16022 15036 16028 15088
rect 16080 15076 16086 15088
rect 17037 15079 17095 15085
rect 17037 15076 17049 15079
rect 16080 15048 17049 15076
rect 16080 15036 16086 15048
rect 17037 15045 17049 15048
rect 17083 15045 17095 15079
rect 17037 15039 17095 15045
rect 18138 15036 18144 15088
rect 18196 15076 18202 15088
rect 18432 15076 18460 15116
rect 18598 15076 18604 15088
rect 18196 15048 18460 15076
rect 18559 15048 18604 15076
rect 18196 15036 18202 15048
rect 18598 15036 18604 15048
rect 18656 15036 18662 15088
rect 18874 15036 18880 15088
rect 18932 15076 18938 15088
rect 19153 15079 19211 15085
rect 19153 15076 19165 15079
rect 18932 15048 19165 15076
rect 18932 15036 18938 15048
rect 19153 15045 19165 15048
rect 19199 15045 19211 15079
rect 19153 15039 19211 15045
rect 19334 15036 19340 15088
rect 19392 15076 19398 15088
rect 19886 15076 19892 15088
rect 19392 15048 19892 15076
rect 19392 15036 19398 15048
rect 19886 15036 19892 15048
rect 19944 15036 19950 15088
rect 17862 14968 17868 15020
rect 17920 15008 17926 15020
rect 17920 14980 18092 15008
rect 17920 14968 17926 14980
rect 10336 14912 12296 14940
rect 10336 14884 10364 14912
rect 12434 14900 12440 14952
rect 12492 14940 12498 14952
rect 12897 14943 12955 14949
rect 12897 14940 12909 14943
rect 12492 14912 12909 14940
rect 12492 14900 12498 14912
rect 12897 14909 12909 14912
rect 12943 14909 12955 14943
rect 12897 14903 12955 14909
rect 13078 14900 13084 14952
rect 13136 14940 13142 14952
rect 14093 14943 14151 14949
rect 14093 14940 14105 14943
rect 13136 14912 14105 14940
rect 13136 14900 13142 14912
rect 14093 14909 14105 14912
rect 14139 14909 14151 14943
rect 14826 14940 14832 14952
rect 14093 14903 14151 14909
rect 14568 14912 14832 14940
rect 8757 14875 8815 14881
rect 8757 14841 8769 14875
rect 8803 14872 8815 14875
rect 9306 14872 9312 14884
rect 8803 14844 9312 14872
rect 8803 14841 8815 14844
rect 8757 14835 8815 14841
rect 9306 14832 9312 14844
rect 9364 14832 9370 14884
rect 10318 14832 10324 14884
rect 10376 14832 10382 14884
rect 10413 14875 10471 14881
rect 10413 14841 10425 14875
rect 10459 14872 10471 14875
rect 12066 14872 12072 14884
rect 10459 14844 12072 14872
rect 10459 14841 10471 14844
rect 10413 14835 10471 14841
rect 12066 14832 12072 14844
rect 12124 14832 12130 14884
rect 14568 14872 14596 14912
rect 14826 14900 14832 14912
rect 14884 14940 14890 14952
rect 15289 14943 15347 14949
rect 14884 14912 15240 14940
rect 14884 14900 14890 14912
rect 12176 14844 14596 14872
rect 11422 14764 11428 14816
rect 11480 14804 11486 14816
rect 12176 14804 12204 14844
rect 14642 14832 14648 14884
rect 14700 14872 14706 14884
rect 15212 14872 15240 14912
rect 15289 14909 15301 14943
rect 15335 14940 15347 14943
rect 15470 14940 15476 14952
rect 15335 14912 15476 14940
rect 15335 14909 15347 14912
rect 15289 14903 15347 14909
rect 15470 14900 15476 14912
rect 15528 14900 15534 14952
rect 15933 14943 15991 14949
rect 15933 14909 15945 14943
rect 15979 14940 15991 14943
rect 16945 14943 17003 14949
rect 16945 14940 16957 14943
rect 15979 14912 16957 14940
rect 15979 14909 15991 14912
rect 15933 14903 15991 14909
rect 16945 14909 16957 14912
rect 16991 14909 17003 14943
rect 17586 14940 17592 14952
rect 17547 14912 17592 14940
rect 16945 14903 17003 14909
rect 16298 14872 16304 14884
rect 14700 14844 14745 14872
rect 15212 14844 16304 14872
rect 14700 14832 14706 14844
rect 16298 14832 16304 14844
rect 16356 14832 16362 14884
rect 16960 14872 16988 14903
rect 17586 14900 17592 14912
rect 17644 14900 17650 14952
rect 18064 14940 18092 14980
rect 19426 14968 19432 15020
rect 19484 15008 19490 15020
rect 19794 15008 19800 15020
rect 19484 14980 19800 15008
rect 19484 14968 19490 14980
rect 19794 14968 19800 14980
rect 19852 14968 19858 15020
rect 19996 15008 20024 15116
rect 20346 15104 20352 15116
rect 20404 15104 20410 15156
rect 21358 15144 21364 15156
rect 21319 15116 21364 15144
rect 21358 15104 21364 15116
rect 21416 15104 21422 15156
rect 24394 15144 24400 15156
rect 22066 15116 24400 15144
rect 20070 15036 20076 15088
rect 20128 15076 20134 15088
rect 22066 15076 22094 15116
rect 24394 15104 24400 15116
rect 24452 15104 24458 15156
rect 24946 15104 24952 15156
rect 25004 15144 25010 15156
rect 25004 15116 26280 15144
rect 25004 15104 25010 15116
rect 22370 15076 22376 15088
rect 20128 15048 22094 15076
rect 22204 15048 22376 15076
rect 20128 15036 20134 15048
rect 20441 15011 20499 15017
rect 20441 15008 20453 15011
rect 19996 14980 20453 15008
rect 20441 14977 20453 14980
rect 20487 15008 20499 15011
rect 20530 15008 20536 15020
rect 20487 14980 20536 15008
rect 20487 14977 20499 14980
rect 20441 14971 20499 14977
rect 20530 14968 20536 14980
rect 20588 14968 20594 15020
rect 21266 15008 21272 15020
rect 21227 14980 21272 15008
rect 21266 14968 21272 14980
rect 21324 14968 21330 15020
rect 21358 14968 21364 15020
rect 21416 15008 21422 15020
rect 22204 15008 22232 15048
rect 22370 15036 22376 15048
rect 22428 15036 22434 15088
rect 22462 15036 22468 15088
rect 22520 15076 22526 15088
rect 22925 15079 22983 15085
rect 22925 15076 22937 15079
rect 22520 15048 22937 15076
rect 22520 15036 22526 15048
rect 22925 15045 22937 15048
rect 22971 15045 22983 15079
rect 23566 15076 23572 15088
rect 23527 15048 23572 15076
rect 22925 15039 22983 15045
rect 23566 15036 23572 15048
rect 23624 15036 23630 15088
rect 24670 15076 24676 15088
rect 24631 15048 24676 15076
rect 24670 15036 24676 15048
rect 24728 15036 24734 15088
rect 24762 15036 24768 15088
rect 24820 15076 24826 15088
rect 25869 15079 25927 15085
rect 24820 15048 24865 15076
rect 24820 15036 24826 15048
rect 25869 15045 25881 15079
rect 25915 15076 25927 15079
rect 25958 15076 25964 15088
rect 25915 15048 25964 15076
rect 25915 15045 25927 15048
rect 25869 15039 25927 15045
rect 25958 15036 25964 15048
rect 26016 15036 26022 15088
rect 26252 15076 26280 15116
rect 26418 15104 26424 15156
rect 26476 15144 26482 15156
rect 28537 15147 28595 15153
rect 28537 15144 28549 15147
rect 26476 15116 28549 15144
rect 26476 15104 26482 15116
rect 28537 15113 28549 15116
rect 28583 15113 28595 15147
rect 28537 15107 28595 15113
rect 27893 15079 27951 15085
rect 27893 15076 27905 15079
rect 26252 15048 27905 15076
rect 27893 15045 27905 15048
rect 27939 15045 27951 15079
rect 27893 15039 27951 15045
rect 27338 15008 27344 15020
rect 21416 14980 22232 15008
rect 27299 14980 27344 15008
rect 21416 14968 21422 14980
rect 27338 14968 27344 14980
rect 27396 14968 27402 15020
rect 27522 14968 27528 15020
rect 27580 15008 27586 15020
rect 27801 15011 27859 15017
rect 27801 15008 27813 15011
rect 27580 14980 27813 15008
rect 27580 14968 27586 14980
rect 27801 14977 27813 14980
rect 27847 14977 27859 15011
rect 28626 15008 28632 15020
rect 28587 14980 28632 15008
rect 27801 14971 27859 14977
rect 28626 14968 28632 14980
rect 28684 15008 28690 15020
rect 29638 15008 29644 15020
rect 28684 14980 29644 15008
rect 28684 14968 28690 14980
rect 29638 14968 29644 14980
rect 29696 14968 29702 15020
rect 18509 14943 18567 14949
rect 18509 14940 18521 14943
rect 18064 14912 18521 14940
rect 18509 14909 18521 14912
rect 18555 14909 18567 14943
rect 18509 14903 18567 14909
rect 19242 14900 19248 14952
rect 19300 14940 19306 14952
rect 21910 14940 21916 14952
rect 19300 14912 21916 14940
rect 19300 14900 19306 14912
rect 21910 14900 21916 14912
rect 21968 14900 21974 14952
rect 22186 14900 22192 14952
rect 22244 14940 22250 14952
rect 22244 14912 22289 14940
rect 22244 14900 22250 14912
rect 22370 14900 22376 14952
rect 22428 14940 22434 14952
rect 22830 14940 22836 14952
rect 22428 14912 22836 14940
rect 22428 14900 22434 14912
rect 22830 14900 22836 14912
rect 22888 14900 22894 14952
rect 23017 14943 23075 14949
rect 23017 14909 23029 14943
rect 23063 14909 23075 14943
rect 23017 14903 23075 14909
rect 20714 14872 20720 14884
rect 16960 14844 20720 14872
rect 20714 14832 20720 14844
rect 20772 14832 20778 14884
rect 22002 14832 22008 14884
rect 22060 14872 22066 14884
rect 23032 14872 23060 14903
rect 24946 14900 24952 14952
rect 25004 14940 25010 14952
rect 25317 14943 25375 14949
rect 25317 14940 25329 14943
rect 25004 14912 25329 14940
rect 25004 14900 25010 14912
rect 25317 14909 25329 14912
rect 25363 14909 25375 14943
rect 25317 14903 25375 14909
rect 25498 14900 25504 14952
rect 25556 14940 25562 14952
rect 25961 14943 26019 14949
rect 25961 14940 25973 14943
rect 25556 14912 25973 14940
rect 25556 14900 25562 14912
rect 25961 14909 25973 14912
rect 26007 14940 26019 14943
rect 26418 14940 26424 14952
rect 26007 14912 26424 14940
rect 26007 14909 26019 14912
rect 25961 14903 26019 14909
rect 26418 14900 26424 14912
rect 26476 14900 26482 14952
rect 24213 14875 24271 14881
rect 22060 14844 24164 14872
rect 22060 14832 22066 14844
rect 11480 14776 12204 14804
rect 12253 14807 12311 14813
rect 11480 14764 11486 14776
rect 12253 14773 12265 14807
rect 12299 14804 12311 14807
rect 17034 14804 17040 14816
rect 12299 14776 17040 14804
rect 12299 14773 12311 14776
rect 12253 14767 12311 14773
rect 17034 14764 17040 14776
rect 17092 14764 17098 14816
rect 19426 14764 19432 14816
rect 19484 14804 19490 14816
rect 19705 14807 19763 14813
rect 19705 14804 19717 14807
rect 19484 14776 19717 14804
rect 19484 14764 19490 14776
rect 19705 14773 19717 14776
rect 19751 14773 19763 14807
rect 19705 14767 19763 14773
rect 23014 14764 23020 14816
rect 23072 14804 23078 14816
rect 23842 14804 23848 14816
rect 23072 14776 23848 14804
rect 23072 14764 23078 14776
rect 23842 14764 23848 14776
rect 23900 14764 23906 14816
rect 24136 14804 24164 14844
rect 24213 14841 24225 14875
rect 24259 14872 24271 14875
rect 24394 14872 24400 14884
rect 24259 14844 24400 14872
rect 24259 14841 24271 14844
rect 24213 14835 24271 14841
rect 24394 14832 24400 14844
rect 24452 14832 24458 14884
rect 28442 14872 28448 14884
rect 26528 14844 28448 14872
rect 26528 14816 26556 14844
rect 28442 14832 28448 14844
rect 28500 14832 28506 14884
rect 25406 14804 25412 14816
rect 24136 14776 25412 14804
rect 25406 14764 25412 14776
rect 25464 14764 25470 14816
rect 26510 14804 26516 14816
rect 26471 14776 26516 14804
rect 26510 14764 26516 14776
rect 26568 14764 26574 14816
rect 26694 14764 26700 14816
rect 26752 14804 26758 14816
rect 27249 14807 27307 14813
rect 27249 14804 27261 14807
rect 26752 14776 27261 14804
rect 26752 14764 26758 14776
rect 27249 14773 27261 14776
rect 27295 14773 27307 14807
rect 27249 14767 27307 14773
rect 28994 14764 29000 14816
rect 29052 14804 29058 14816
rect 29089 14807 29147 14813
rect 29089 14804 29101 14807
rect 29052 14776 29101 14804
rect 29052 14764 29058 14776
rect 29089 14773 29101 14776
rect 29135 14773 29147 14807
rect 29089 14767 29147 14773
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 3418 14560 3424 14612
rect 3476 14600 3482 14612
rect 11974 14600 11980 14612
rect 3476 14572 11980 14600
rect 3476 14560 3482 14572
rect 11974 14560 11980 14572
rect 12032 14560 12038 14612
rect 12158 14560 12164 14612
rect 12216 14600 12222 14612
rect 21358 14600 21364 14612
rect 12216 14572 21364 14600
rect 12216 14560 12222 14572
rect 21358 14560 21364 14572
rect 21416 14560 21422 14612
rect 21910 14560 21916 14612
rect 21968 14600 21974 14612
rect 23934 14600 23940 14612
rect 21968 14572 23940 14600
rect 21968 14560 21974 14572
rect 23934 14560 23940 14572
rect 23992 14560 23998 14612
rect 24670 14560 24676 14612
rect 24728 14600 24734 14612
rect 27985 14603 28043 14609
rect 27985 14600 27997 14603
rect 24728 14572 27997 14600
rect 24728 14560 24734 14572
rect 27985 14569 27997 14572
rect 28031 14569 28043 14603
rect 27985 14563 28043 14569
rect 9125 14535 9183 14541
rect 9125 14532 9137 14535
rect 1872 14504 9137 14532
rect 1872 14405 1900 14504
rect 9125 14501 9137 14504
rect 9171 14501 9183 14535
rect 9125 14495 9183 14501
rect 11149 14535 11207 14541
rect 11149 14501 11161 14535
rect 11195 14532 11207 14535
rect 12250 14532 12256 14544
rect 11195 14504 12256 14532
rect 11195 14501 11207 14504
rect 11149 14495 11207 14501
rect 12250 14492 12256 14504
rect 12308 14492 12314 14544
rect 12437 14535 12495 14541
rect 12437 14501 12449 14535
rect 12483 14532 12495 14535
rect 17494 14532 17500 14544
rect 12483 14504 17500 14532
rect 12483 14501 12495 14504
rect 12437 14495 12495 14501
rect 17494 14492 17500 14504
rect 17552 14492 17558 14544
rect 18690 14492 18696 14544
rect 18748 14532 18754 14544
rect 20714 14532 20720 14544
rect 18748 14504 20720 14532
rect 18748 14492 18754 14504
rect 20714 14492 20720 14504
rect 20772 14532 20778 14544
rect 20901 14535 20959 14541
rect 20772 14504 20852 14532
rect 20772 14492 20778 14504
rect 8573 14467 8631 14473
rect 8573 14433 8585 14467
rect 8619 14464 8631 14467
rect 9398 14464 9404 14476
rect 8619 14436 9404 14464
rect 8619 14433 8631 14436
rect 8573 14427 8631 14433
rect 9398 14424 9404 14436
rect 9456 14464 9462 14476
rect 14553 14467 14611 14473
rect 9456 14436 10456 14464
rect 9456 14424 9462 14436
rect 1857 14399 1915 14405
rect 1857 14365 1869 14399
rect 1903 14365 1915 14399
rect 9306 14396 9312 14408
rect 9267 14368 9312 14396
rect 1857 14359 1915 14365
rect 9306 14356 9312 14368
rect 9364 14356 9370 14408
rect 9766 14396 9772 14408
rect 9727 14368 9772 14396
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 10428 14405 10456 14436
rect 14553 14433 14565 14467
rect 14599 14464 14611 14467
rect 16758 14464 16764 14476
rect 14599 14436 16764 14464
rect 14599 14433 14611 14436
rect 14553 14427 14611 14433
rect 16758 14424 16764 14436
rect 16816 14424 16822 14476
rect 16942 14464 16948 14476
rect 16903 14436 16948 14464
rect 16942 14424 16948 14436
rect 17000 14424 17006 14476
rect 17402 14424 17408 14476
rect 17460 14464 17466 14476
rect 17589 14467 17647 14473
rect 17589 14464 17601 14467
rect 17460 14436 17601 14464
rect 17460 14424 17466 14436
rect 17589 14433 17601 14436
rect 17635 14433 17647 14467
rect 17589 14427 17647 14433
rect 18785 14467 18843 14473
rect 18785 14433 18797 14467
rect 18831 14464 18843 14467
rect 19426 14464 19432 14476
rect 18831 14436 19432 14464
rect 18831 14433 18843 14436
rect 18785 14427 18843 14433
rect 19426 14424 19432 14436
rect 19484 14424 19490 14476
rect 20346 14464 20352 14476
rect 20307 14436 20352 14464
rect 20346 14424 20352 14436
rect 20404 14424 20410 14476
rect 20824 14464 20852 14504
rect 20901 14501 20913 14535
rect 20947 14532 20959 14535
rect 22002 14532 22008 14544
rect 20947 14504 22008 14532
rect 20947 14501 20959 14504
rect 20901 14495 20959 14501
rect 22002 14492 22008 14504
rect 22060 14492 22066 14544
rect 23661 14535 23719 14541
rect 23661 14532 23673 14535
rect 22480 14504 23673 14532
rect 22480 14473 22508 14504
rect 23661 14501 23673 14504
rect 23707 14532 23719 14535
rect 24946 14532 24952 14544
rect 23707 14504 24952 14532
rect 23707 14501 23719 14504
rect 23661 14495 23719 14501
rect 24946 14492 24952 14504
rect 25004 14492 25010 14544
rect 25038 14492 25044 14544
rect 25096 14532 25102 14544
rect 29733 14535 29791 14541
rect 29733 14532 29745 14535
rect 25096 14504 29745 14532
rect 25096 14492 25102 14504
rect 22465 14467 22523 14473
rect 20824 14436 21588 14464
rect 10413 14399 10471 14405
rect 10413 14365 10425 14399
rect 10459 14365 10471 14399
rect 10413 14359 10471 14365
rect 10502 14356 10508 14408
rect 10560 14396 10566 14408
rect 11241 14399 11299 14405
rect 10560 14368 10605 14396
rect 10560 14356 10566 14368
rect 11241 14365 11253 14399
rect 11287 14396 11299 14399
rect 11974 14396 11980 14408
rect 11287 14368 11980 14396
rect 11287 14365 11299 14368
rect 11241 14359 11299 14365
rect 11974 14356 11980 14368
rect 12032 14356 12038 14408
rect 12526 14396 12532 14408
rect 12487 14368 12532 14396
rect 12526 14356 12532 14368
rect 12584 14356 12590 14408
rect 13814 14356 13820 14408
rect 13872 14396 13878 14408
rect 14366 14396 14372 14408
rect 13872 14368 14372 14396
rect 13872 14356 13878 14368
rect 14366 14356 14372 14368
rect 14424 14396 14430 14408
rect 14461 14399 14519 14405
rect 14461 14396 14473 14399
rect 14424 14368 14473 14396
rect 14424 14356 14430 14368
rect 14461 14365 14473 14368
rect 14507 14396 14519 14399
rect 14918 14396 14924 14408
rect 14507 14368 14924 14396
rect 14507 14365 14519 14368
rect 14461 14359 14519 14365
rect 14918 14356 14924 14368
rect 14976 14356 14982 14408
rect 16298 14396 16304 14408
rect 16259 14368 16304 14396
rect 16298 14356 16304 14368
rect 16356 14356 16362 14408
rect 16390 14356 16396 14408
rect 16448 14356 16454 14408
rect 17954 14356 17960 14408
rect 18012 14396 18018 14408
rect 18141 14399 18199 14405
rect 18141 14396 18153 14399
rect 18012 14368 18153 14396
rect 18012 14356 18018 14368
rect 18141 14365 18153 14368
rect 18187 14365 18199 14399
rect 18141 14359 18199 14365
rect 19334 14356 19340 14408
rect 19392 14396 19398 14408
rect 19613 14399 19671 14405
rect 19613 14396 19625 14399
rect 19392 14368 19625 14396
rect 19392 14356 19398 14368
rect 19613 14365 19625 14368
rect 19659 14365 19671 14399
rect 19613 14359 19671 14365
rect 9861 14331 9919 14337
rect 9861 14297 9873 14331
rect 9907 14328 9919 14331
rect 13078 14328 13084 14340
rect 9907 14300 13084 14328
rect 9907 14297 9919 14300
rect 9861 14291 9919 14297
rect 13078 14288 13084 14300
rect 13136 14288 13142 14340
rect 13170 14288 13176 14340
rect 13228 14328 13234 14340
rect 13722 14328 13728 14340
rect 13228 14300 13273 14328
rect 13683 14300 13728 14328
rect 13228 14288 13234 14300
rect 13722 14288 13728 14300
rect 13780 14288 13786 14340
rect 14734 14288 14740 14340
rect 14792 14328 14798 14340
rect 15105 14331 15163 14337
rect 15105 14328 15117 14331
rect 14792 14300 15117 14328
rect 14792 14288 14798 14300
rect 15105 14297 15117 14300
rect 15151 14297 15163 14331
rect 15105 14291 15163 14297
rect 15657 14331 15715 14337
rect 15657 14297 15669 14331
rect 15703 14297 15715 14331
rect 15657 14291 15715 14297
rect 15749 14331 15807 14337
rect 15749 14297 15761 14331
rect 15795 14328 15807 14331
rect 16408 14328 16436 14356
rect 17494 14328 17500 14340
rect 15795 14300 16436 14328
rect 17455 14300 17500 14328
rect 15795 14297 15807 14300
rect 15749 14291 15807 14297
rect 1670 14260 1676 14272
rect 1631 14232 1676 14260
rect 1670 14220 1676 14232
rect 1728 14220 1734 14272
rect 11882 14260 11888 14272
rect 11843 14232 11888 14260
rect 11882 14220 11888 14232
rect 11940 14220 11946 14272
rect 14182 14220 14188 14272
rect 14240 14260 14246 14272
rect 15672 14260 15700 14291
rect 17494 14288 17500 14300
rect 17552 14288 17558 14340
rect 18693 14331 18751 14337
rect 18693 14297 18705 14331
rect 18739 14297 18751 14331
rect 18693 14291 18751 14297
rect 14240 14232 15700 14260
rect 16393 14263 16451 14269
rect 14240 14220 14246 14232
rect 16393 14229 16405 14263
rect 16439 14260 16451 14263
rect 18708 14260 18736 14291
rect 18966 14288 18972 14340
rect 19024 14328 19030 14340
rect 20441 14331 20499 14337
rect 19024 14300 20392 14328
rect 19024 14288 19030 14300
rect 16439 14232 18736 14260
rect 19705 14263 19763 14269
rect 16439 14229 16451 14232
rect 16393 14223 16451 14229
rect 19705 14229 19717 14263
rect 19751 14260 19763 14263
rect 20162 14260 20168 14272
rect 19751 14232 20168 14260
rect 19751 14229 19763 14232
rect 19705 14223 19763 14229
rect 20162 14220 20168 14232
rect 20220 14220 20226 14272
rect 20364 14260 20392 14300
rect 20441 14297 20453 14331
rect 20487 14328 20499 14331
rect 20806 14328 20812 14340
rect 20487 14300 20812 14328
rect 20487 14297 20499 14300
rect 20441 14291 20499 14297
rect 20806 14288 20812 14300
rect 20864 14288 20870 14340
rect 20990 14288 20996 14340
rect 21048 14328 21054 14340
rect 21453 14331 21511 14337
rect 21453 14328 21465 14331
rect 21048 14300 21465 14328
rect 21048 14288 21054 14300
rect 21453 14297 21465 14300
rect 21499 14297 21511 14331
rect 21453 14291 21511 14297
rect 21358 14260 21364 14272
rect 20364 14232 21364 14260
rect 21358 14220 21364 14232
rect 21416 14220 21422 14272
rect 21560 14260 21588 14436
rect 22465 14433 22477 14467
rect 22511 14433 22523 14467
rect 22465 14427 22523 14433
rect 23106 14424 23112 14476
rect 23164 14464 23170 14476
rect 23164 14436 23209 14464
rect 23164 14424 23170 14436
rect 23382 14424 23388 14476
rect 23440 14464 23446 14476
rect 24857 14467 24915 14473
rect 24857 14464 24869 14467
rect 23440 14436 24869 14464
rect 23440 14424 23446 14436
rect 24857 14433 24869 14436
rect 24903 14433 24915 14467
rect 24857 14427 24915 14433
rect 25130 14424 25136 14476
rect 25188 14464 25194 14476
rect 27341 14467 27399 14473
rect 27341 14464 27353 14467
rect 25188 14436 27353 14464
rect 25188 14424 25194 14436
rect 27341 14433 27353 14436
rect 27387 14433 27399 14467
rect 27341 14427 27399 14433
rect 26970 14396 26976 14408
rect 26896 14368 26976 14396
rect 22370 14328 22376 14340
rect 22331 14300 22376 14328
rect 22370 14288 22376 14300
rect 22428 14288 22434 14340
rect 22922 14288 22928 14340
rect 22980 14328 22986 14340
rect 23201 14331 23259 14337
rect 23201 14328 23213 14331
rect 22980 14300 23213 14328
rect 22980 14288 22986 14300
rect 23201 14297 23213 14300
rect 23247 14297 23259 14331
rect 23201 14291 23259 14297
rect 25409 14331 25467 14337
rect 25409 14297 25421 14331
rect 25455 14297 25467 14331
rect 25409 14291 25467 14297
rect 24026 14260 24032 14272
rect 21560 14232 24032 14260
rect 24026 14220 24032 14232
rect 24084 14220 24090 14272
rect 25424 14260 25452 14291
rect 25498 14288 25504 14340
rect 25556 14328 25562 14340
rect 25556 14300 25601 14328
rect 25556 14288 25562 14300
rect 25958 14288 25964 14340
rect 26016 14328 26022 14340
rect 26053 14331 26111 14337
rect 26053 14328 26065 14331
rect 26016 14300 26065 14328
rect 26016 14288 26022 14300
rect 26053 14297 26065 14300
rect 26099 14297 26111 14331
rect 26602 14328 26608 14340
rect 26563 14300 26608 14328
rect 26053 14291 26111 14297
rect 26602 14288 26608 14300
rect 26660 14288 26666 14340
rect 26697 14331 26755 14337
rect 26697 14297 26709 14331
rect 26743 14328 26755 14331
rect 26896 14328 26924 14368
rect 26970 14356 26976 14368
rect 27028 14356 27034 14408
rect 27448 14405 27476 14504
rect 29733 14501 29745 14504
rect 29779 14501 29791 14535
rect 29733 14495 29791 14501
rect 28994 14464 29000 14476
rect 28092 14436 29000 14464
rect 27433 14399 27491 14405
rect 27433 14365 27445 14399
rect 27479 14365 27491 14399
rect 27433 14359 27491 14365
rect 27522 14356 27528 14408
rect 27580 14396 27586 14408
rect 28092 14405 28120 14436
rect 28994 14424 29000 14436
rect 29052 14424 29058 14476
rect 28077 14399 28135 14405
rect 28077 14396 28089 14399
rect 27580 14368 28089 14396
rect 27580 14356 27586 14368
rect 28077 14365 28089 14368
rect 28123 14365 28135 14399
rect 28534 14396 28540 14408
rect 28495 14368 28540 14396
rect 28077 14359 28135 14365
rect 28534 14356 28540 14368
rect 28592 14356 28598 14408
rect 28629 14331 28687 14337
rect 28629 14328 28641 14331
rect 26743 14300 26924 14328
rect 26988 14300 28641 14328
rect 26743 14297 26755 14300
rect 26697 14291 26755 14297
rect 26988 14260 27016 14300
rect 28629 14297 28641 14300
rect 28675 14297 28687 14331
rect 28629 14291 28687 14297
rect 25424 14232 27016 14260
rect 27062 14220 27068 14272
rect 27120 14260 27126 14272
rect 27522 14260 27528 14272
rect 27120 14232 27528 14260
rect 27120 14220 27126 14232
rect 27522 14220 27528 14232
rect 27580 14220 27586 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 9217 14059 9275 14065
rect 9217 14025 9229 14059
rect 9263 14056 9275 14059
rect 11606 14056 11612 14068
rect 9263 14028 11612 14056
rect 9263 14025 9275 14028
rect 9217 14019 9275 14025
rect 11606 14016 11612 14028
rect 11664 14016 11670 14068
rect 11882 14016 11888 14068
rect 11940 14056 11946 14068
rect 12434 14056 12440 14068
rect 11940 14028 12440 14056
rect 11940 14016 11946 14028
rect 12434 14016 12440 14028
rect 12492 14016 12498 14068
rect 18414 14056 18420 14068
rect 12912 14028 18420 14056
rect 8021 13991 8079 13997
rect 8021 13957 8033 13991
rect 8067 13988 8079 13991
rect 9766 13988 9772 14000
rect 8067 13960 9772 13988
rect 8067 13957 8079 13960
rect 8021 13951 8079 13957
rect 9766 13948 9772 13960
rect 9824 13988 9830 14000
rect 9824 13960 9904 13988
rect 9824 13948 9830 13960
rect 9876 13929 9904 13960
rect 10318 13948 10324 14000
rect 10376 13988 10382 14000
rect 10413 13991 10471 13997
rect 10413 13988 10425 13991
rect 10376 13960 10425 13988
rect 10376 13948 10382 13960
rect 10413 13957 10425 13960
rect 10459 13957 10471 13991
rect 11238 13988 11244 14000
rect 10413 13951 10471 13957
rect 10520 13960 11244 13988
rect 10520 13929 10548 13960
rect 11238 13948 11244 13960
rect 11296 13948 11302 14000
rect 12912 13997 12940 14028
rect 18414 14016 18420 14028
rect 18472 14016 18478 14068
rect 18601 14059 18659 14065
rect 18601 14025 18613 14059
rect 18647 14056 18659 14059
rect 18647 14028 20392 14056
rect 18647 14025 18659 14028
rect 18601 14019 18659 14025
rect 12805 13991 12863 13997
rect 12805 13988 12817 13991
rect 11348 13960 12817 13988
rect 8573 13923 8631 13929
rect 8573 13889 8585 13923
rect 8619 13920 8631 13923
rect 9861 13923 9919 13929
rect 8619 13892 9812 13920
rect 8619 13889 8631 13892
rect 8573 13883 8631 13889
rect 7834 13812 7840 13864
rect 7892 13852 7898 13864
rect 9784 13852 9812 13892
rect 9861 13889 9873 13923
rect 9907 13889 9919 13923
rect 9861 13883 9919 13889
rect 10505 13923 10563 13929
rect 10505 13889 10517 13923
rect 10551 13889 10563 13923
rect 10505 13883 10563 13889
rect 10965 13923 11023 13929
rect 10965 13889 10977 13923
rect 11011 13889 11023 13923
rect 10965 13883 11023 13889
rect 10870 13852 10876 13864
rect 7892 13824 9720 13852
rect 9784 13824 10876 13852
rect 7892 13812 7898 13824
rect 9692 13793 9720 13824
rect 10870 13812 10876 13824
rect 10928 13852 10934 13864
rect 10980 13852 11008 13883
rect 11146 13880 11152 13932
rect 11204 13920 11210 13932
rect 11348 13920 11376 13960
rect 12805 13957 12817 13960
rect 12851 13957 12863 13991
rect 12805 13951 12863 13957
rect 12897 13991 12955 13997
rect 12897 13957 12909 13991
rect 12943 13957 12955 13991
rect 12897 13951 12955 13957
rect 13633 13991 13691 13997
rect 13633 13957 13645 13991
rect 13679 13988 13691 13991
rect 13906 13988 13912 14000
rect 13679 13960 13912 13988
rect 13679 13957 13691 13960
rect 13633 13951 13691 13957
rect 13906 13948 13912 13960
rect 13964 13948 13970 14000
rect 15565 13991 15623 13997
rect 15565 13988 15577 13991
rect 14384 13960 15577 13988
rect 11204 13892 11376 13920
rect 11204 13880 11210 13892
rect 11422 13880 11428 13932
rect 11480 13920 11486 13932
rect 11701 13923 11759 13929
rect 11701 13920 11713 13923
rect 11480 13892 11713 13920
rect 11480 13880 11486 13892
rect 11701 13889 11713 13892
rect 11747 13889 11759 13923
rect 11701 13883 11759 13889
rect 10928 13824 11008 13852
rect 11057 13855 11115 13861
rect 10928 13812 10934 13824
rect 11057 13821 11069 13855
rect 11103 13852 11115 13855
rect 11103 13824 13308 13852
rect 11103 13821 11115 13824
rect 11057 13815 11115 13821
rect 9677 13787 9735 13793
rect 9677 13753 9689 13787
rect 9723 13753 9735 13787
rect 9677 13747 9735 13753
rect 11238 13744 11244 13796
rect 11296 13784 11302 13796
rect 12342 13784 12348 13796
rect 11296 13756 11836 13784
rect 12303 13756 12348 13784
rect 11296 13744 11302 13756
rect 7926 13676 7932 13728
rect 7984 13716 7990 13728
rect 11698 13716 11704 13728
rect 7984 13688 11704 13716
rect 7984 13676 7990 13688
rect 11698 13676 11704 13688
rect 11756 13676 11762 13728
rect 11808 13716 11836 13756
rect 12342 13744 12348 13756
rect 12400 13744 12406 13796
rect 12434 13744 12440 13796
rect 12492 13784 12498 13796
rect 12802 13784 12808 13796
rect 12492 13756 12808 13784
rect 12492 13744 12498 13756
rect 12802 13744 12808 13756
rect 12860 13744 12866 13796
rect 12526 13716 12532 13728
rect 11808 13688 12532 13716
rect 12526 13676 12532 13688
rect 12584 13676 12590 13728
rect 13280 13716 13308 13824
rect 13354 13812 13360 13864
rect 13412 13852 13418 13864
rect 13541 13855 13599 13861
rect 13541 13852 13553 13855
rect 13412 13824 13553 13852
rect 13412 13812 13418 13824
rect 13541 13821 13553 13824
rect 13587 13852 13599 13855
rect 13630 13852 13636 13864
rect 13587 13824 13636 13852
rect 13587 13821 13599 13824
rect 13541 13815 13599 13821
rect 13630 13812 13636 13824
rect 13688 13812 13694 13864
rect 13814 13812 13820 13864
rect 13872 13852 13878 13864
rect 14384 13852 14412 13960
rect 15565 13957 15577 13960
rect 15611 13957 15623 13991
rect 15565 13951 15623 13957
rect 15657 13991 15715 13997
rect 15657 13957 15669 13991
rect 15703 13988 15715 13991
rect 16666 13988 16672 14000
rect 15703 13960 16672 13988
rect 15703 13957 15715 13960
rect 15657 13951 15715 13957
rect 16666 13948 16672 13960
rect 16724 13948 16730 14000
rect 17034 13988 17040 14000
rect 16995 13960 17040 13988
rect 17034 13948 17040 13960
rect 17092 13948 17098 14000
rect 19058 13948 19064 14000
rect 19116 13988 19122 14000
rect 19153 13991 19211 13997
rect 19153 13988 19165 13991
rect 19116 13960 19165 13988
rect 19116 13948 19122 13960
rect 19153 13957 19165 13960
rect 19199 13957 19211 13991
rect 19153 13951 19211 13957
rect 19705 13991 19763 13997
rect 19705 13957 19717 13991
rect 19751 13988 19763 13991
rect 20254 13988 20260 14000
rect 19751 13960 20260 13988
rect 19751 13957 19763 13960
rect 19705 13951 19763 13957
rect 20254 13948 20260 13960
rect 20312 13948 20318 14000
rect 16209 13923 16267 13929
rect 16209 13889 16221 13923
rect 16255 13920 16267 13923
rect 16298 13920 16304 13932
rect 16255 13892 16304 13920
rect 16255 13889 16267 13892
rect 16209 13883 16267 13889
rect 13872 13824 14412 13852
rect 13872 13812 13878 13824
rect 14458 13812 14464 13864
rect 14516 13852 14522 13864
rect 14516 13824 14561 13852
rect 14516 13812 14522 13824
rect 14642 13812 14648 13864
rect 14700 13852 14706 13864
rect 14918 13852 14924 13864
rect 14700 13824 14924 13852
rect 14700 13812 14706 13824
rect 14918 13812 14924 13824
rect 14976 13852 14982 13864
rect 16224 13852 16252 13883
rect 16298 13880 16304 13892
rect 16356 13880 16362 13932
rect 18690 13920 18696 13932
rect 18651 13892 18696 13920
rect 18690 13880 18696 13892
rect 18748 13880 18754 13932
rect 16942 13852 16948 13864
rect 14976 13824 16252 13852
rect 16903 13824 16948 13852
rect 14976 13812 14982 13824
rect 16942 13812 16948 13824
rect 17000 13812 17006 13864
rect 17589 13855 17647 13861
rect 17589 13821 17601 13855
rect 17635 13852 17647 13855
rect 19150 13852 19156 13864
rect 17635 13824 19156 13852
rect 17635 13821 17647 13824
rect 17589 13815 17647 13821
rect 19150 13812 19156 13824
rect 19208 13812 19214 13864
rect 19426 13812 19432 13864
rect 19484 13852 19490 13864
rect 19797 13855 19855 13861
rect 19797 13852 19809 13855
rect 19484 13824 19809 13852
rect 19484 13812 19490 13824
rect 19797 13821 19809 13824
rect 19843 13821 19855 13855
rect 20364 13852 20392 14028
rect 20438 14016 20444 14068
rect 20496 14056 20502 14068
rect 22005 14059 22063 14065
rect 22005 14056 22017 14059
rect 20496 14028 22017 14056
rect 20496 14016 20502 14028
rect 22005 14025 22017 14028
rect 22051 14025 22063 14059
rect 22005 14019 22063 14025
rect 28258 14016 28264 14068
rect 28316 14056 28322 14068
rect 29181 14059 29239 14065
rect 29181 14056 29193 14059
rect 28316 14028 29193 14056
rect 28316 14016 28322 14028
rect 29181 14025 29193 14028
rect 29227 14025 29239 14059
rect 29181 14019 29239 14025
rect 20625 13991 20683 13997
rect 20625 13957 20637 13991
rect 20671 13988 20683 13991
rect 20671 13960 22094 13988
rect 20671 13957 20683 13960
rect 20625 13951 20683 13957
rect 20533 13923 20591 13929
rect 20533 13889 20545 13923
rect 20579 13920 20591 13923
rect 20806 13920 20812 13932
rect 20579 13892 20812 13920
rect 20579 13889 20591 13892
rect 20533 13883 20591 13889
rect 20806 13880 20812 13892
rect 20864 13880 20870 13932
rect 21174 13880 21180 13932
rect 21232 13920 21238 13932
rect 21361 13923 21419 13929
rect 21361 13920 21373 13923
rect 21232 13892 21373 13920
rect 21232 13880 21238 13892
rect 21361 13889 21373 13892
rect 21407 13889 21419 13923
rect 22066 13920 22094 13960
rect 23106 13948 23112 14000
rect 23164 13988 23170 14000
rect 23293 13991 23351 13997
rect 23293 13988 23305 13991
rect 23164 13960 23305 13988
rect 23164 13948 23170 13960
rect 23293 13957 23305 13960
rect 23339 13957 23351 13991
rect 23293 13951 23351 13957
rect 23382 13948 23388 14000
rect 23440 13988 23446 14000
rect 23934 13988 23940 14000
rect 23440 13960 23485 13988
rect 23847 13960 23940 13988
rect 23440 13948 23446 13960
rect 23934 13948 23940 13960
rect 23992 13988 23998 14000
rect 25314 13988 25320 14000
rect 23992 13960 25320 13988
rect 23992 13948 23998 13960
rect 25314 13948 25320 13960
rect 25372 13948 25378 14000
rect 25406 13948 25412 14000
rect 25464 13988 25470 14000
rect 25501 13991 25559 13997
rect 25501 13988 25513 13991
rect 25464 13960 25513 13988
rect 25464 13948 25470 13960
rect 25501 13957 25513 13960
rect 25547 13988 25559 13991
rect 25958 13988 25964 14000
rect 25547 13960 25964 13988
rect 25547 13957 25559 13960
rect 25501 13951 25559 13957
rect 25958 13948 25964 13960
rect 26016 13948 26022 14000
rect 26053 13991 26111 13997
rect 26053 13957 26065 13991
rect 26099 13988 26111 13991
rect 28537 13991 28595 13997
rect 28537 13988 28549 13991
rect 26099 13960 28549 13988
rect 26099 13957 26111 13960
rect 26053 13951 26111 13957
rect 28537 13957 28549 13960
rect 28583 13957 28595 13991
rect 28537 13951 28595 13957
rect 22465 13923 22523 13929
rect 22465 13920 22477 13923
rect 22066 13892 22477 13920
rect 21361 13883 21419 13889
rect 22465 13889 22477 13892
rect 22511 13889 22523 13923
rect 22465 13883 22523 13889
rect 24026 13880 24032 13932
rect 24084 13920 24090 13932
rect 24397 13923 24455 13929
rect 24397 13920 24409 13923
rect 24084 13892 24409 13920
rect 24084 13880 24090 13892
rect 24397 13889 24409 13892
rect 24443 13920 24455 13923
rect 24443 13892 25452 13920
rect 24443 13889 24455 13892
rect 24397 13883 24455 13889
rect 21266 13852 21272 13864
rect 20364 13824 21128 13852
rect 21227 13824 21272 13852
rect 19797 13815 19855 13821
rect 13906 13744 13912 13796
rect 13964 13784 13970 13796
rect 14734 13784 14740 13796
rect 13964 13756 14740 13784
rect 13964 13744 13970 13756
rect 14734 13744 14740 13756
rect 14792 13744 14798 13796
rect 18138 13784 18144 13796
rect 15304 13756 18144 13784
rect 14550 13716 14556 13728
rect 13280 13688 14556 13716
rect 14550 13676 14556 13688
rect 14608 13676 14614 13728
rect 14642 13676 14648 13728
rect 14700 13716 14706 13728
rect 15304 13716 15332 13756
rect 18138 13744 18144 13756
rect 18196 13744 18202 13796
rect 18230 13744 18236 13796
rect 18288 13784 18294 13796
rect 21100 13784 21128 13824
rect 21266 13812 21272 13824
rect 21324 13812 21330 13864
rect 21818 13852 21824 13864
rect 21376 13824 21824 13852
rect 21376 13784 21404 13824
rect 21818 13812 21824 13824
rect 21876 13812 21882 13864
rect 22649 13855 22707 13861
rect 22649 13821 22661 13855
rect 22695 13852 22707 13855
rect 23382 13852 23388 13864
rect 22695 13824 23388 13852
rect 22695 13821 22707 13824
rect 22649 13815 22707 13821
rect 23382 13812 23388 13824
rect 23440 13812 23446 13864
rect 24489 13855 24547 13861
rect 24489 13821 24501 13855
rect 24535 13852 24547 13855
rect 25038 13852 25044 13864
rect 24535 13824 25044 13852
rect 24535 13821 24547 13824
rect 24489 13815 24547 13821
rect 25038 13812 25044 13824
rect 25096 13812 25102 13864
rect 18288 13756 20760 13784
rect 21100 13756 21404 13784
rect 18288 13744 18294 13756
rect 14700 13688 15332 13716
rect 14700 13676 14706 13688
rect 16206 13676 16212 13728
rect 16264 13716 16270 13728
rect 20622 13716 20628 13728
rect 16264 13688 20628 13716
rect 16264 13676 16270 13688
rect 20622 13676 20628 13688
rect 20680 13676 20686 13728
rect 20732 13716 20760 13756
rect 21726 13744 21732 13796
rect 21784 13784 21790 13796
rect 21784 13756 23428 13784
rect 21784 13744 21790 13756
rect 22002 13716 22008 13728
rect 20732 13688 22008 13716
rect 22002 13676 22008 13688
rect 22060 13676 22066 13728
rect 23400 13716 23428 13756
rect 24026 13744 24032 13796
rect 24084 13784 24090 13796
rect 25424 13784 25452 13892
rect 26878 13880 26884 13932
rect 26936 13920 26942 13932
rect 27338 13920 27344 13932
rect 26936 13892 27344 13920
rect 26936 13880 26942 13892
rect 27338 13880 27344 13892
rect 27396 13880 27402 13932
rect 27522 13880 27528 13932
rect 27580 13920 27586 13932
rect 27985 13923 28043 13929
rect 27985 13920 27997 13923
rect 27580 13892 27997 13920
rect 27580 13880 27586 13892
rect 27985 13889 27997 13892
rect 28031 13889 28043 13923
rect 27985 13883 28043 13889
rect 25774 13812 25780 13864
rect 25832 13852 25838 13864
rect 26145 13855 26203 13861
rect 26145 13852 26157 13855
rect 25832 13824 26157 13852
rect 25832 13812 25838 13824
rect 26145 13821 26157 13824
rect 26191 13821 26203 13855
rect 27246 13852 27252 13864
rect 26145 13815 26203 13821
rect 26252 13824 27252 13852
rect 26252 13784 26280 13824
rect 27246 13812 27252 13824
rect 27304 13812 27310 13864
rect 27890 13852 27896 13864
rect 27851 13824 27896 13852
rect 27890 13812 27896 13824
rect 27948 13812 27954 13864
rect 28000 13852 28028 13883
rect 28074 13880 28080 13932
rect 28132 13920 28138 13932
rect 28629 13923 28687 13929
rect 28629 13920 28641 13923
rect 28132 13892 28641 13920
rect 28132 13880 28138 13892
rect 28629 13889 28641 13892
rect 28675 13920 28687 13923
rect 28718 13920 28724 13932
rect 28675 13892 28724 13920
rect 28675 13889 28687 13892
rect 28629 13883 28687 13889
rect 28718 13880 28724 13892
rect 28776 13880 28782 13932
rect 29270 13920 29276 13932
rect 29231 13892 29276 13920
rect 29270 13880 29276 13892
rect 29328 13920 29334 13932
rect 29454 13920 29460 13932
rect 29328 13892 29460 13920
rect 29328 13880 29334 13892
rect 29454 13880 29460 13892
rect 29512 13920 29518 13932
rect 30285 13923 30343 13929
rect 30285 13920 30297 13923
rect 29512 13892 30297 13920
rect 29512 13880 29518 13892
rect 30285 13889 30297 13892
rect 30331 13889 30343 13923
rect 30285 13883 30343 13889
rect 37553 13923 37611 13929
rect 37553 13889 37565 13923
rect 37599 13920 37611 13923
rect 38194 13920 38200 13932
rect 37599 13892 38200 13920
rect 37599 13889 37611 13892
rect 37553 13883 37611 13889
rect 38194 13880 38200 13892
rect 38252 13880 38258 13932
rect 29733 13855 29791 13861
rect 29733 13852 29745 13855
rect 28000 13824 29745 13852
rect 29733 13821 29745 13824
rect 29779 13821 29791 13855
rect 29733 13815 29791 13821
rect 29822 13812 29828 13864
rect 29880 13852 29886 13864
rect 38013 13855 38071 13861
rect 38013 13852 38025 13855
rect 29880 13824 38025 13852
rect 29880 13812 29886 13824
rect 38013 13821 38025 13824
rect 38059 13821 38071 13855
rect 38013 13815 38071 13821
rect 27614 13784 27620 13796
rect 24084 13756 25360 13784
rect 25424 13756 26280 13784
rect 27080 13756 27620 13784
rect 24084 13744 24090 13756
rect 24670 13716 24676 13728
rect 23400 13688 24676 13716
rect 24670 13676 24676 13688
rect 24728 13676 24734 13728
rect 25332 13716 25360 13756
rect 27080 13716 27108 13756
rect 27614 13744 27620 13756
rect 27672 13744 27678 13796
rect 27246 13716 27252 13728
rect 25332 13688 27108 13716
rect 27207 13688 27252 13716
rect 27246 13676 27252 13688
rect 27304 13676 27310 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 9401 13515 9459 13521
rect 9401 13481 9413 13515
rect 9447 13512 9459 13515
rect 10962 13512 10968 13524
rect 9447 13484 10968 13512
rect 9447 13481 9459 13484
rect 9401 13475 9459 13481
rect 10962 13472 10968 13484
rect 11020 13472 11026 13524
rect 13538 13512 13544 13524
rect 11072 13484 13544 13512
rect 9122 13404 9128 13456
rect 9180 13444 9186 13456
rect 11072 13444 11100 13484
rect 13538 13472 13544 13484
rect 13596 13472 13602 13524
rect 13722 13512 13728 13524
rect 13648 13484 13728 13512
rect 9180 13416 11100 13444
rect 9180 13404 9186 13416
rect 11698 13404 11704 13456
rect 11756 13444 11762 13456
rect 12158 13444 12164 13456
rect 11756 13416 12164 13444
rect 11756 13404 11762 13416
rect 12158 13404 12164 13416
rect 12216 13404 12222 13456
rect 12529 13447 12587 13453
rect 12529 13413 12541 13447
rect 12575 13444 12587 13447
rect 13354 13444 13360 13456
rect 12575 13416 13360 13444
rect 12575 13413 12587 13416
rect 12529 13407 12587 13413
rect 13354 13404 13360 13416
rect 13412 13404 13418 13456
rect 13648 13453 13676 13484
rect 13722 13472 13728 13484
rect 13780 13512 13786 13524
rect 16206 13512 16212 13524
rect 13780 13484 16212 13512
rect 13780 13472 13786 13484
rect 13633 13447 13691 13453
rect 13633 13413 13645 13447
rect 13679 13413 13691 13447
rect 13633 13407 13691 13413
rect 14458 13404 14464 13456
rect 14516 13444 14522 13456
rect 16040 13453 16068 13484
rect 16206 13472 16212 13484
rect 16264 13472 16270 13524
rect 16298 13472 16304 13524
rect 16356 13512 16362 13524
rect 18230 13512 18236 13524
rect 16356 13484 18236 13512
rect 16356 13472 16362 13484
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 18598 13472 18604 13524
rect 18656 13512 18662 13524
rect 21726 13512 21732 13524
rect 18656 13484 21732 13512
rect 18656 13472 18662 13484
rect 21726 13472 21732 13484
rect 21784 13472 21790 13524
rect 22002 13472 22008 13524
rect 22060 13512 22066 13524
rect 27062 13512 27068 13524
rect 22060 13484 25912 13512
rect 27023 13484 27068 13512
rect 22060 13472 22066 13484
rect 16025 13447 16083 13453
rect 14516 13416 15608 13444
rect 14516 13404 14522 13416
rect 8573 13379 8631 13385
rect 8573 13345 8585 13379
rect 8619 13376 8631 13379
rect 11054 13376 11060 13388
rect 8619 13348 11060 13376
rect 8619 13345 8631 13348
rect 8573 13339 8631 13345
rect 11054 13336 11060 13348
rect 11112 13336 11118 13388
rect 15473 13379 15531 13385
rect 15473 13376 15485 13379
rect 11164 13348 15485 13376
rect 6917 13311 6975 13317
rect 6917 13277 6929 13311
rect 6963 13308 6975 13311
rect 8846 13308 8852 13320
rect 6963 13280 8852 13308
rect 6963 13277 6975 13280
rect 6917 13271 6975 13277
rect 8846 13268 8852 13280
rect 8904 13308 8910 13320
rect 9309 13311 9367 13317
rect 9309 13308 9321 13311
rect 8904 13280 9321 13308
rect 8904 13268 8910 13280
rect 9309 13277 9321 13280
rect 9355 13277 9367 13311
rect 9953 13311 10011 13317
rect 9953 13308 9965 13311
rect 9309 13271 9367 13277
rect 9876 13280 9965 13308
rect 9876 13252 9904 13280
rect 9953 13277 9965 13280
rect 9999 13277 10011 13311
rect 9953 13271 10011 13277
rect 10781 13311 10839 13317
rect 10781 13277 10793 13311
rect 10827 13308 10839 13311
rect 11164 13308 11192 13348
rect 15473 13345 15485 13348
rect 15519 13345 15531 13379
rect 15580 13376 15608 13416
rect 16025 13413 16037 13447
rect 16071 13413 16083 13447
rect 16025 13407 16083 13413
rect 16224 13416 23336 13444
rect 16224 13376 16252 13416
rect 18506 13376 18512 13388
rect 15580 13348 16252 13376
rect 18467 13348 18512 13376
rect 15473 13339 15531 13345
rect 18506 13336 18512 13348
rect 18564 13336 18570 13388
rect 18785 13379 18843 13385
rect 18785 13345 18797 13379
rect 18831 13376 18843 13379
rect 19058 13376 19064 13388
rect 18831 13348 19064 13376
rect 18831 13345 18843 13348
rect 18785 13339 18843 13345
rect 19058 13336 19064 13348
rect 19116 13336 19122 13388
rect 19518 13376 19524 13388
rect 19431 13348 19524 13376
rect 19518 13336 19524 13348
rect 19576 13376 19582 13388
rect 19886 13376 19892 13388
rect 19576 13348 19892 13376
rect 19576 13336 19582 13348
rect 19886 13336 19892 13348
rect 19944 13336 19950 13388
rect 21729 13379 21787 13385
rect 21729 13345 21741 13379
rect 21775 13376 21787 13379
rect 21910 13376 21916 13388
rect 21775 13348 21916 13376
rect 21775 13345 21787 13348
rect 21729 13339 21787 13345
rect 21910 13336 21916 13348
rect 21968 13336 21974 13388
rect 23014 13376 23020 13388
rect 22975 13348 23020 13376
rect 23014 13336 23020 13348
rect 23072 13336 23078 13388
rect 23308 13376 23336 13416
rect 23382 13404 23388 13456
rect 23440 13444 23446 13456
rect 25774 13444 25780 13456
rect 23440 13416 25780 13444
rect 23440 13404 23446 13416
rect 23934 13376 23940 13388
rect 23308 13348 23940 13376
rect 23934 13336 23940 13348
rect 23992 13336 23998 13388
rect 24029 13379 24087 13385
rect 24029 13345 24041 13379
rect 24075 13376 24087 13379
rect 24118 13376 24124 13388
rect 24075 13348 24124 13376
rect 24075 13345 24087 13348
rect 24029 13339 24087 13345
rect 24118 13336 24124 13348
rect 24176 13336 24182 13388
rect 24946 13376 24952 13388
rect 24907 13348 24952 13376
rect 24946 13336 24952 13348
rect 25004 13336 25010 13388
rect 25240 13385 25268 13416
rect 25774 13404 25780 13416
rect 25832 13404 25838 13456
rect 25884 13385 25912 13484
rect 27062 13472 27068 13484
rect 27120 13472 27126 13524
rect 27338 13472 27344 13524
rect 27396 13512 27402 13524
rect 28905 13515 28963 13521
rect 28905 13512 28917 13515
rect 27396 13484 28917 13512
rect 27396 13472 27402 13484
rect 28905 13481 28917 13484
rect 28951 13481 28963 13515
rect 28905 13475 28963 13481
rect 25958 13404 25964 13456
rect 26016 13444 26022 13456
rect 28626 13444 28632 13456
rect 26016 13416 28632 13444
rect 26016 13404 26022 13416
rect 28626 13404 28632 13416
rect 28684 13404 28690 13456
rect 25225 13379 25283 13385
rect 25225 13345 25237 13379
rect 25271 13345 25283 13379
rect 25225 13339 25283 13345
rect 25869 13379 25927 13385
rect 25869 13345 25881 13379
rect 25915 13345 25927 13379
rect 25869 13339 25927 13345
rect 26050 13336 26056 13388
rect 26108 13376 26114 13388
rect 28534 13376 28540 13388
rect 26108 13348 28540 13376
rect 26108 13336 26114 13348
rect 28534 13336 28540 13348
rect 28592 13336 28598 13388
rect 28718 13336 28724 13388
rect 28776 13376 28782 13388
rect 29733 13379 29791 13385
rect 29733 13376 29745 13379
rect 28776 13348 29745 13376
rect 28776 13336 28782 13348
rect 29733 13345 29745 13348
rect 29779 13345 29791 13379
rect 29733 13339 29791 13345
rect 10827 13280 11192 13308
rect 10827 13277 10839 13280
rect 10781 13271 10839 13277
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 11296 13280 11341 13308
rect 11296 13268 11302 13280
rect 11790 13268 11796 13320
rect 11848 13308 11854 13320
rect 11885 13311 11943 13317
rect 11885 13308 11897 13311
rect 11848 13280 11897 13308
rect 11848 13268 11854 13280
rect 11885 13277 11897 13280
rect 11931 13277 11943 13311
rect 12066 13308 12072 13320
rect 12027 13280 12072 13308
rect 11885 13271 11943 13277
rect 12066 13268 12072 13280
rect 12124 13268 12130 13320
rect 12158 13268 12164 13320
rect 12216 13308 12222 13320
rect 14458 13308 14464 13320
rect 12216 13280 12480 13308
rect 14419 13280 14464 13308
rect 12216 13268 12222 13280
rect 7469 13243 7527 13249
rect 7469 13209 7481 13243
rect 7515 13240 7527 13243
rect 9858 13240 9864 13252
rect 7515 13212 9864 13240
rect 7515 13209 7527 13212
rect 7469 13203 7527 13209
rect 9858 13200 9864 13212
rect 9916 13200 9922 13252
rect 10045 13243 10103 13249
rect 10045 13209 10057 13243
rect 10091 13240 10103 13243
rect 12342 13240 12348 13252
rect 10091 13212 12348 13240
rect 10091 13209 10103 13212
rect 10045 13203 10103 13209
rect 12342 13200 12348 13212
rect 12400 13200 12406 13252
rect 12452 13240 12480 13280
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 20254 13268 20260 13320
rect 20312 13308 20318 13320
rect 20898 13308 20904 13320
rect 20312 13280 20904 13308
rect 20312 13268 20318 13280
rect 20898 13268 20904 13280
rect 20956 13268 20962 13320
rect 13078 13240 13084 13252
rect 12452 13212 13084 13240
rect 13078 13200 13084 13212
rect 13136 13200 13142 13252
rect 13173 13243 13231 13249
rect 13173 13209 13185 13243
rect 13219 13209 13231 13243
rect 13173 13203 13231 13209
rect 8021 13175 8079 13181
rect 8021 13141 8033 13175
rect 8067 13172 8079 13175
rect 10594 13172 10600 13184
rect 8067 13144 10600 13172
rect 8067 13141 8079 13144
rect 8021 13135 8079 13141
rect 10594 13132 10600 13144
rect 10652 13172 10658 13184
rect 10962 13172 10968 13184
rect 10652 13144 10968 13172
rect 10652 13132 10658 13144
rect 10962 13132 10968 13144
rect 11020 13132 11026 13184
rect 11333 13175 11391 13181
rect 11333 13141 11345 13175
rect 11379 13172 11391 13175
rect 11790 13172 11796 13184
rect 11379 13144 11796 13172
rect 11379 13141 11391 13144
rect 11333 13135 11391 13141
rect 11790 13132 11796 13144
rect 11848 13132 11854 13184
rect 12250 13132 12256 13184
rect 12308 13172 12314 13184
rect 13188 13172 13216 13203
rect 13354 13200 13360 13252
rect 13412 13240 13418 13252
rect 13412 13212 14504 13240
rect 13412 13200 13418 13212
rect 12308 13144 13216 13172
rect 12308 13132 12314 13144
rect 13814 13132 13820 13184
rect 13872 13172 13878 13184
rect 14369 13175 14427 13181
rect 14369 13172 14381 13175
rect 13872 13144 14381 13172
rect 13872 13132 13878 13144
rect 14369 13141 14381 13144
rect 14415 13141 14427 13175
rect 14476 13172 14504 13212
rect 14550 13200 14556 13252
rect 14608 13240 14614 13252
rect 15565 13243 15623 13249
rect 15565 13240 15577 13243
rect 14608 13212 15577 13240
rect 14608 13200 14614 13212
rect 15565 13209 15577 13212
rect 15611 13209 15623 13243
rect 15565 13203 15623 13209
rect 16669 13243 16727 13249
rect 16669 13209 16681 13243
rect 16715 13209 16727 13243
rect 16669 13203 16727 13209
rect 15470 13172 15476 13184
rect 14476 13144 15476 13172
rect 14369 13135 14427 13141
rect 15470 13132 15476 13144
rect 15528 13172 15534 13184
rect 16684 13172 16712 13203
rect 16758 13200 16764 13252
rect 16816 13240 16822 13252
rect 17313 13243 17371 13249
rect 16816 13212 16861 13240
rect 16816 13200 16822 13212
rect 17313 13209 17325 13243
rect 17359 13240 17371 13243
rect 18230 13240 18236 13252
rect 17359 13212 18236 13240
rect 17359 13209 17371 13212
rect 17313 13203 17371 13209
rect 18230 13200 18236 13212
rect 18288 13200 18294 13252
rect 18693 13243 18751 13249
rect 18693 13209 18705 13243
rect 18739 13209 18751 13243
rect 19610 13240 19616 13252
rect 19571 13212 19616 13240
rect 18693 13203 18751 13209
rect 15528 13144 16712 13172
rect 18708 13172 18736 13203
rect 19610 13200 19616 13212
rect 19668 13200 19674 13252
rect 20165 13243 20223 13249
rect 20165 13209 20177 13243
rect 20211 13240 20223 13243
rect 20346 13240 20352 13252
rect 20211 13212 20352 13240
rect 20211 13209 20223 13212
rect 20165 13203 20223 13209
rect 20346 13200 20352 13212
rect 20404 13200 20410 13252
rect 21082 13200 21088 13252
rect 21140 13240 21146 13252
rect 21913 13243 21971 13249
rect 21913 13240 21925 13243
rect 21140 13212 21925 13240
rect 21140 13200 21146 13212
rect 21913 13209 21925 13212
rect 21959 13209 21971 13243
rect 21913 13203 21971 13209
rect 22005 13243 22063 13249
rect 22005 13209 22017 13243
rect 22051 13209 22063 13243
rect 22005 13203 22063 13209
rect 23109 13243 23167 13249
rect 23109 13209 23121 13243
rect 23155 13240 23167 13243
rect 24026 13240 24032 13252
rect 23155 13212 24032 13240
rect 23155 13209 23167 13212
rect 23109 13203 23167 13209
rect 20530 13172 20536 13184
rect 18708 13144 20536 13172
rect 15528 13132 15534 13144
rect 20530 13132 20536 13144
rect 20588 13132 20594 13184
rect 22020 13172 22048 13203
rect 24026 13200 24032 13212
rect 24084 13200 24090 13252
rect 24136 13240 24164 13336
rect 26513 13311 26571 13317
rect 26513 13277 26525 13311
rect 26559 13308 26571 13311
rect 26786 13308 26792 13320
rect 26559 13280 26792 13308
rect 26559 13277 26571 13280
rect 26513 13271 26571 13277
rect 26786 13268 26792 13280
rect 26844 13268 26850 13320
rect 26970 13308 26976 13320
rect 26931 13280 26976 13308
rect 26970 13268 26976 13280
rect 27028 13268 27034 13320
rect 24946 13240 24952 13252
rect 24136 13212 24952 13240
rect 24946 13200 24952 13212
rect 25004 13200 25010 13252
rect 25130 13240 25136 13252
rect 25091 13212 25136 13240
rect 25130 13200 25136 13212
rect 25188 13200 25194 13252
rect 25222 13200 25228 13252
rect 25280 13240 25286 13252
rect 25682 13240 25688 13252
rect 25280 13212 25688 13240
rect 25280 13200 25286 13212
rect 25682 13200 25688 13212
rect 25740 13200 25746 13252
rect 25961 13243 26019 13249
rect 25961 13209 25973 13243
rect 26007 13240 26019 13243
rect 27522 13240 27528 13252
rect 26007 13212 27528 13240
rect 26007 13209 26019 13212
rect 25961 13203 26019 13209
rect 27522 13200 27528 13212
rect 27580 13200 27586 13252
rect 27617 13243 27675 13249
rect 27617 13209 27629 13243
rect 27663 13240 27675 13243
rect 27798 13240 27804 13252
rect 27663 13212 27804 13240
rect 27663 13209 27675 13212
rect 27617 13203 27675 13209
rect 27798 13200 27804 13212
rect 27856 13200 27862 13252
rect 28166 13240 28172 13252
rect 28127 13212 28172 13240
rect 28166 13200 28172 13212
rect 28224 13200 28230 13252
rect 28258 13200 28264 13252
rect 28316 13240 28322 13252
rect 28316 13212 28409 13240
rect 28316 13200 28322 13212
rect 23474 13172 23480 13184
rect 22020 13144 23480 13172
rect 23474 13132 23480 13144
rect 23532 13132 23538 13184
rect 24118 13132 24124 13184
rect 24176 13172 24182 13184
rect 26694 13172 26700 13184
rect 24176 13144 26700 13172
rect 24176 13132 24182 13144
rect 26694 13132 26700 13144
rect 26752 13132 26758 13184
rect 27062 13132 27068 13184
rect 27120 13172 27126 13184
rect 28276 13172 28304 13200
rect 27120 13144 28304 13172
rect 27120 13132 27126 13144
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 7837 12971 7895 12977
rect 7837 12937 7849 12971
rect 7883 12968 7895 12971
rect 7926 12968 7932 12980
rect 7883 12940 7932 12968
rect 7883 12937 7895 12940
rect 7837 12931 7895 12937
rect 7926 12928 7932 12940
rect 7984 12928 7990 12980
rect 9122 12968 9128 12980
rect 9083 12940 9128 12968
rect 9122 12928 9128 12940
rect 9180 12928 9186 12980
rect 11974 12928 11980 12980
rect 12032 12968 12038 12980
rect 13446 12968 13452 12980
rect 12032 12940 13452 12968
rect 12032 12928 12038 12940
rect 13446 12928 13452 12940
rect 13504 12928 13510 12980
rect 18230 12928 18236 12980
rect 18288 12968 18294 12980
rect 18690 12968 18696 12980
rect 18288 12940 18696 12968
rect 18288 12928 18294 12940
rect 18690 12928 18696 12940
rect 18748 12928 18754 12980
rect 19426 12928 19432 12980
rect 19484 12968 19490 12980
rect 19613 12971 19671 12977
rect 19613 12968 19625 12971
rect 19484 12940 19625 12968
rect 19484 12928 19490 12940
rect 19613 12937 19625 12940
rect 19659 12937 19671 12971
rect 19613 12931 19671 12937
rect 19720 12940 20576 12968
rect 6733 12903 6791 12909
rect 6733 12869 6745 12903
rect 6779 12900 6791 12903
rect 9674 12900 9680 12912
rect 6779 12872 9680 12900
rect 6779 12869 6791 12872
rect 6733 12863 6791 12869
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12832 1915 12835
rect 5534 12832 5540 12844
rect 1903 12804 5540 12832
rect 1903 12801 1915 12804
rect 1857 12795 1915 12801
rect 5534 12792 5540 12804
rect 5592 12792 5598 12844
rect 7742 12832 7748 12844
rect 7703 12804 7748 12832
rect 7742 12792 7748 12804
rect 7800 12792 7806 12844
rect 8404 12841 8432 12872
rect 9674 12860 9680 12872
rect 9732 12860 9738 12912
rect 10428 12872 11100 12900
rect 8389 12835 8447 12841
rect 8389 12801 8401 12835
rect 8435 12801 8447 12835
rect 9030 12832 9036 12844
rect 8389 12795 8447 12801
rect 8588 12804 9036 12832
rect 7285 12767 7343 12773
rect 7285 12733 7297 12767
rect 7331 12764 7343 12767
rect 8588 12764 8616 12804
rect 9030 12792 9036 12804
rect 9088 12792 9094 12844
rect 9858 12832 9864 12844
rect 9819 12804 9864 12832
rect 9858 12792 9864 12804
rect 9916 12792 9922 12844
rect 7331 12736 8616 12764
rect 9769 12767 9827 12773
rect 7331 12733 7343 12736
rect 7285 12727 7343 12733
rect 9769 12733 9781 12767
rect 9815 12764 9827 12767
rect 10428 12764 10456 12872
rect 10505 12835 10563 12841
rect 10505 12801 10517 12835
rect 10551 12832 10563 12835
rect 10686 12832 10692 12844
rect 10551 12804 10692 12832
rect 10551 12801 10563 12804
rect 10505 12795 10563 12801
rect 10686 12792 10692 12804
rect 10744 12792 10750 12844
rect 10962 12832 10968 12844
rect 10923 12804 10968 12832
rect 10962 12792 10968 12804
rect 11020 12792 11026 12844
rect 11072 12832 11100 12872
rect 11146 12860 11152 12912
rect 11204 12900 11210 12912
rect 11514 12900 11520 12912
rect 11204 12872 11520 12900
rect 11204 12860 11210 12872
rect 11514 12860 11520 12872
rect 11572 12860 11578 12912
rect 11606 12860 11612 12912
rect 11664 12900 11670 12912
rect 11793 12903 11851 12909
rect 11793 12900 11805 12903
rect 11664 12872 11805 12900
rect 11664 12860 11670 12872
rect 11793 12869 11805 12872
rect 11839 12869 11851 12903
rect 11793 12863 11851 12869
rect 11885 12903 11943 12909
rect 11885 12869 11897 12903
rect 11931 12900 11943 12903
rect 12066 12900 12072 12912
rect 11931 12872 12072 12900
rect 11931 12869 11943 12872
rect 11885 12863 11943 12869
rect 12066 12860 12072 12872
rect 12124 12860 12130 12912
rect 13357 12903 13415 12909
rect 13357 12900 13369 12903
rect 12912 12872 13369 12900
rect 11072 12804 11284 12832
rect 9815 12736 10456 12764
rect 11256 12764 11284 12804
rect 12912 12764 12940 12872
rect 13357 12869 13369 12872
rect 13403 12869 13415 12903
rect 13357 12863 13415 12869
rect 14921 12903 14979 12909
rect 14921 12869 14933 12903
rect 14967 12900 14979 12903
rect 15378 12900 15384 12912
rect 14967 12872 15384 12900
rect 14967 12869 14979 12872
rect 14921 12863 14979 12869
rect 15378 12860 15384 12872
rect 15436 12860 15442 12912
rect 15749 12903 15807 12909
rect 15749 12869 15761 12903
rect 15795 12900 15807 12903
rect 17218 12900 17224 12912
rect 15795 12872 17224 12900
rect 15795 12869 15807 12872
rect 15749 12863 15807 12869
rect 17218 12860 17224 12872
rect 17276 12860 17282 12912
rect 18049 12903 18107 12909
rect 18049 12900 18061 12903
rect 17328 12872 18061 12900
rect 16301 12835 16359 12841
rect 16301 12801 16313 12835
rect 16347 12832 16359 12835
rect 16390 12832 16396 12844
rect 16347 12804 16396 12832
rect 16347 12801 16359 12804
rect 16301 12795 16359 12801
rect 16390 12792 16396 12804
rect 16448 12792 16454 12844
rect 11256 12752 11560 12764
rect 11900 12752 12940 12764
rect 11256 12736 12940 12752
rect 9815 12733 9827 12736
rect 9769 12727 9827 12733
rect 11532 12724 11928 12736
rect 13078 12724 13084 12776
rect 13136 12764 13142 12776
rect 13265 12767 13323 12773
rect 13265 12764 13277 12767
rect 13136 12736 13277 12764
rect 13136 12724 13142 12736
rect 13265 12733 13277 12736
rect 13311 12733 13323 12767
rect 13265 12727 13323 12733
rect 14182 12724 14188 12776
rect 14240 12764 14246 12776
rect 14734 12764 14740 12776
rect 14240 12736 14740 12764
rect 14240 12724 14246 12736
rect 14734 12724 14740 12736
rect 14792 12724 14798 12776
rect 15010 12764 15016 12776
rect 14971 12736 15016 12764
rect 15010 12724 15016 12736
rect 15068 12724 15074 12776
rect 15470 12724 15476 12776
rect 15528 12764 15534 12776
rect 15657 12767 15715 12773
rect 15657 12764 15669 12767
rect 15528 12736 15669 12764
rect 15528 12724 15534 12736
rect 15657 12733 15669 12736
rect 15703 12733 15715 12767
rect 17328 12764 17356 12872
rect 18049 12869 18061 12872
rect 18095 12869 18107 12903
rect 18049 12863 18107 12869
rect 18322 12860 18328 12912
rect 18380 12900 18386 12912
rect 19720 12900 19748 12940
rect 20438 12900 20444 12912
rect 18380 12872 19748 12900
rect 20399 12872 20444 12900
rect 18380 12860 18386 12872
rect 20438 12860 20444 12872
rect 20496 12860 20502 12912
rect 20548 12909 20576 12940
rect 20806 12928 20812 12980
rect 20864 12968 20870 12980
rect 22738 12968 22744 12980
rect 20864 12940 22744 12968
rect 20864 12928 20870 12940
rect 22738 12928 22744 12940
rect 22796 12968 22802 12980
rect 22796 12940 24348 12968
rect 22796 12928 22802 12940
rect 20533 12903 20591 12909
rect 20533 12869 20545 12903
rect 20579 12869 20591 12903
rect 20533 12863 20591 12869
rect 21358 12860 21364 12912
rect 21416 12900 21422 12912
rect 21453 12903 21511 12909
rect 21453 12900 21465 12903
rect 21416 12872 21465 12900
rect 21416 12860 21422 12872
rect 21453 12869 21465 12872
rect 21499 12900 21511 12903
rect 21726 12900 21732 12912
rect 21499 12872 21732 12900
rect 21499 12869 21511 12872
rect 21453 12863 21511 12869
rect 21726 12860 21732 12872
rect 21784 12860 21790 12912
rect 22833 12903 22891 12909
rect 22833 12869 22845 12903
rect 22879 12900 22891 12903
rect 22922 12900 22928 12912
rect 22879 12872 22928 12900
rect 22879 12869 22891 12872
rect 22833 12863 22891 12869
rect 22922 12860 22928 12872
rect 22980 12860 22986 12912
rect 23474 12900 23480 12912
rect 23435 12872 23480 12900
rect 23474 12860 23480 12872
rect 23532 12860 23538 12912
rect 24029 12903 24087 12909
rect 24029 12869 24041 12903
rect 24075 12900 24087 12903
rect 24118 12900 24124 12912
rect 24075 12872 24124 12900
rect 24075 12869 24087 12872
rect 24029 12863 24087 12869
rect 24118 12860 24124 12872
rect 24176 12860 24182 12912
rect 17402 12792 17408 12844
rect 17460 12832 17466 12844
rect 17770 12832 17776 12844
rect 17460 12804 17776 12832
rect 17460 12792 17466 12804
rect 17770 12792 17776 12804
rect 17828 12792 17834 12844
rect 18800 12804 20116 12832
rect 15657 12727 15715 12733
rect 15764 12736 17356 12764
rect 17957 12767 18015 12773
rect 8481 12699 8539 12705
rect 8481 12665 8493 12699
rect 8527 12696 8539 12699
rect 12066 12696 12072 12708
rect 8527 12668 12072 12696
rect 8527 12665 8539 12668
rect 8481 12659 8539 12665
rect 12066 12656 12072 12668
rect 12124 12656 12130 12708
rect 12342 12696 12348 12708
rect 12303 12668 12348 12696
rect 12342 12656 12348 12668
rect 12400 12656 12406 12708
rect 13817 12699 13875 12705
rect 13817 12665 13829 12699
rect 13863 12696 13875 12699
rect 14918 12696 14924 12708
rect 13863 12668 14924 12696
rect 13863 12665 13875 12668
rect 13817 12659 13875 12665
rect 14918 12656 14924 12668
rect 14976 12656 14982 12708
rect 1670 12628 1676 12640
rect 1631 12600 1676 12628
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 10413 12631 10471 12637
rect 10413 12597 10425 12631
rect 10459 12628 10471 12631
rect 10778 12628 10784 12640
rect 10459 12600 10784 12628
rect 10459 12597 10471 12600
rect 10413 12591 10471 12597
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 11057 12631 11115 12637
rect 11057 12597 11069 12631
rect 11103 12628 11115 12631
rect 15764 12628 15792 12736
rect 17957 12733 17969 12767
rect 18003 12764 18015 12767
rect 18230 12764 18236 12776
rect 18003 12736 18236 12764
rect 18003 12733 18015 12736
rect 17957 12727 18015 12733
rect 18230 12724 18236 12736
rect 18288 12724 18294 12776
rect 18506 12764 18512 12776
rect 18419 12736 18512 12764
rect 18506 12724 18512 12736
rect 18564 12764 18570 12776
rect 18800 12764 18828 12804
rect 18564 12736 18828 12764
rect 18564 12724 18570 12736
rect 19334 12724 19340 12776
rect 19392 12764 19398 12776
rect 19518 12764 19524 12776
rect 19392 12736 19524 12764
rect 19392 12724 19398 12736
rect 19518 12724 19524 12736
rect 19576 12724 19582 12776
rect 20088 12764 20116 12804
rect 23382 12792 23388 12844
rect 23440 12832 23446 12844
rect 23440 12804 23520 12832
rect 23440 12792 23446 12804
rect 20990 12764 20996 12776
rect 20088 12736 20996 12764
rect 20990 12724 20996 12736
rect 21048 12724 21054 12776
rect 22278 12764 22284 12776
rect 22239 12736 22284 12764
rect 22278 12724 22284 12736
rect 22336 12724 22342 12776
rect 22925 12767 22983 12773
rect 22925 12733 22937 12767
rect 22971 12733 22983 12767
rect 23492 12764 23520 12804
rect 24121 12767 24179 12773
rect 24121 12764 24133 12767
rect 23492 12736 24133 12764
rect 22925 12727 22983 12733
rect 24121 12733 24133 12736
rect 24167 12733 24179 12767
rect 24320 12764 24348 12940
rect 25866 12928 25872 12980
rect 25924 12968 25930 12980
rect 25961 12971 26019 12977
rect 25961 12968 25973 12971
rect 25924 12940 25973 12968
rect 25924 12928 25930 12940
rect 25961 12937 25973 12940
rect 26007 12937 26019 12971
rect 25961 12931 26019 12937
rect 27522 12928 27528 12980
rect 27580 12968 27586 12980
rect 28537 12971 28595 12977
rect 28537 12968 28549 12971
rect 27580 12940 28549 12968
rect 27580 12928 27586 12940
rect 28537 12937 28549 12940
rect 28583 12937 28595 12971
rect 35894 12968 35900 12980
rect 28537 12931 28595 12937
rect 29656 12940 35900 12968
rect 24670 12900 24676 12912
rect 24631 12872 24676 12900
rect 24670 12860 24676 12872
rect 24728 12860 24734 12912
rect 25038 12860 25044 12912
rect 25096 12900 25102 12912
rect 25248 12903 25306 12909
rect 25248 12900 25260 12903
rect 25096 12872 25260 12900
rect 25096 12860 25102 12872
rect 25248 12869 25260 12872
rect 25294 12869 25306 12903
rect 25248 12863 25306 12869
rect 25774 12860 25780 12912
rect 25832 12900 25838 12912
rect 29656 12909 29684 12940
rect 35894 12928 35900 12940
rect 35952 12928 35958 12980
rect 27249 12903 27307 12909
rect 27249 12900 27261 12903
rect 25832 12872 27261 12900
rect 25832 12860 25838 12872
rect 27249 12869 27261 12872
rect 27295 12869 27307 12903
rect 29641 12903 29699 12909
rect 29641 12900 29653 12903
rect 27249 12863 27307 12869
rect 27356 12872 29653 12900
rect 25682 12832 25688 12844
rect 25516 12804 25688 12832
rect 25317 12767 25375 12773
rect 24320 12736 24900 12764
rect 24121 12727 24179 12733
rect 17313 12699 17371 12705
rect 17313 12665 17325 12699
rect 17359 12696 17371 12699
rect 22940 12696 22968 12727
rect 23382 12696 23388 12708
rect 17359 12668 23388 12696
rect 17359 12665 17371 12668
rect 17313 12659 17371 12665
rect 23382 12656 23388 12668
rect 23440 12656 23446 12708
rect 24872 12696 24900 12736
rect 25317 12733 25329 12767
rect 25363 12764 25375 12767
rect 25516 12764 25544 12804
rect 25682 12792 25688 12804
rect 25740 12792 25746 12844
rect 26050 12832 26056 12844
rect 26011 12804 26056 12832
rect 26050 12792 26056 12804
rect 26108 12792 26114 12844
rect 27356 12841 27384 12872
rect 29641 12869 29653 12872
rect 29687 12869 29699 12903
rect 29641 12863 29699 12869
rect 27341 12835 27399 12841
rect 27341 12832 27353 12835
rect 26620 12804 27353 12832
rect 25363 12736 25544 12764
rect 25363 12733 25375 12736
rect 25317 12727 25375 12733
rect 26513 12699 26571 12705
rect 26513 12696 26525 12699
rect 24872 12668 26525 12696
rect 26513 12665 26525 12668
rect 26559 12665 26571 12699
rect 26513 12659 26571 12665
rect 11103 12600 15792 12628
rect 11103 12597 11115 12600
rect 11057 12591 11115 12597
rect 15930 12588 15936 12640
rect 15988 12628 15994 12640
rect 18506 12628 18512 12640
rect 15988 12600 18512 12628
rect 15988 12588 15994 12600
rect 18506 12588 18512 12600
rect 18564 12588 18570 12640
rect 18690 12588 18696 12640
rect 18748 12628 18754 12640
rect 21542 12628 21548 12640
rect 18748 12600 21548 12628
rect 18748 12588 18754 12600
rect 21542 12588 21548 12600
rect 21600 12628 21606 12640
rect 22922 12628 22928 12640
rect 21600 12600 22928 12628
rect 21600 12588 21606 12600
rect 22922 12588 22928 12600
rect 22980 12588 22986 12640
rect 23934 12588 23940 12640
rect 23992 12628 23998 12640
rect 26620 12628 26648 12804
rect 27341 12801 27353 12804
rect 27387 12801 27399 12835
rect 27341 12795 27399 12801
rect 27985 12835 28043 12841
rect 27985 12801 27997 12835
rect 28031 12801 28043 12835
rect 28626 12832 28632 12844
rect 28587 12804 28632 12832
rect 27985 12795 28043 12801
rect 28000 12764 28028 12795
rect 28626 12792 28632 12804
rect 28684 12832 28690 12844
rect 30745 12835 30803 12841
rect 30745 12832 30757 12835
rect 28684 12804 30757 12832
rect 28684 12792 28690 12804
rect 30745 12801 30757 12804
rect 30791 12801 30803 12835
rect 30745 12795 30803 12801
rect 28718 12764 28724 12776
rect 28000 12736 28724 12764
rect 28718 12724 28724 12736
rect 28776 12764 28782 12776
rect 30193 12767 30251 12773
rect 30193 12764 30205 12767
rect 28776 12736 30205 12764
rect 28776 12724 28782 12736
rect 30193 12733 30205 12736
rect 30239 12733 30251 12767
rect 30193 12727 30251 12733
rect 27706 12656 27712 12708
rect 27764 12696 27770 12708
rect 27893 12699 27951 12705
rect 27893 12696 27905 12699
rect 27764 12668 27905 12696
rect 27764 12656 27770 12668
rect 27893 12665 27905 12668
rect 27939 12665 27951 12699
rect 27893 12659 27951 12665
rect 23992 12600 26648 12628
rect 23992 12588 23998 12600
rect 27522 12588 27528 12640
rect 27580 12628 27586 12640
rect 29089 12631 29147 12637
rect 29089 12628 29101 12631
rect 27580 12600 29101 12628
rect 27580 12588 27586 12600
rect 29089 12597 29101 12600
rect 29135 12597 29147 12631
rect 29089 12591 29147 12597
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 7837 12427 7895 12433
rect 7837 12424 7849 12427
rect 5592 12396 7849 12424
rect 5592 12384 5598 12396
rect 7837 12393 7849 12396
rect 7883 12393 7895 12427
rect 7837 12387 7895 12393
rect 9309 12427 9367 12433
rect 9309 12393 9321 12427
rect 9355 12424 9367 12427
rect 10134 12424 10140 12436
rect 9355 12396 10140 12424
rect 9355 12393 9367 12396
rect 9309 12387 9367 12393
rect 10134 12384 10140 12396
rect 10192 12384 10198 12436
rect 10597 12427 10655 12433
rect 10597 12393 10609 12427
rect 10643 12424 10655 12427
rect 10778 12424 10784 12436
rect 10643 12396 10784 12424
rect 10643 12393 10655 12396
rect 10597 12387 10655 12393
rect 10778 12384 10784 12396
rect 10836 12384 10842 12436
rect 11238 12424 11244 12436
rect 11199 12396 11244 12424
rect 11238 12384 11244 12396
rect 11296 12384 11302 12436
rect 19702 12424 19708 12436
rect 12360 12396 19708 12424
rect 7285 12359 7343 12365
rect 7285 12325 7297 12359
rect 7331 12356 7343 12359
rect 9766 12356 9772 12368
rect 7331 12328 9772 12356
rect 7331 12325 7343 12328
rect 7285 12319 7343 12325
rect 9766 12316 9772 12328
rect 9824 12316 9830 12368
rect 11146 12316 11152 12368
rect 11204 12356 11210 12368
rect 12360 12356 12388 12396
rect 19702 12384 19708 12396
rect 19760 12384 19766 12436
rect 20346 12424 20352 12436
rect 19812 12396 20352 12424
rect 11204 12328 12388 12356
rect 12437 12359 12495 12365
rect 11204 12316 11210 12328
rect 12437 12325 12449 12359
rect 12483 12356 12495 12359
rect 13170 12356 13176 12368
rect 12483 12328 13176 12356
rect 12483 12325 12495 12328
rect 12437 12319 12495 12325
rect 13170 12316 13176 12328
rect 13228 12316 13234 12368
rect 13446 12316 13452 12368
rect 13504 12356 13510 12368
rect 14550 12356 14556 12368
rect 13504 12328 14556 12356
rect 13504 12316 13510 12328
rect 14550 12316 14556 12328
rect 14608 12356 14614 12368
rect 16390 12356 16396 12368
rect 14608 12328 16396 12356
rect 14608 12316 14614 12328
rect 16390 12316 16396 12328
rect 16448 12356 16454 12368
rect 17034 12356 17040 12368
rect 16448 12328 17040 12356
rect 16448 12316 16454 12328
rect 17034 12316 17040 12328
rect 17092 12356 17098 12368
rect 18785 12359 18843 12365
rect 17092 12328 17540 12356
rect 17092 12316 17098 12328
rect 12894 12288 12900 12300
rect 7944 12260 12900 12288
rect 7944 12229 7972 12260
rect 12894 12248 12900 12260
rect 12952 12248 12958 12300
rect 13081 12291 13139 12297
rect 13081 12257 13093 12291
rect 13127 12288 13139 12291
rect 13354 12288 13360 12300
rect 13127 12260 13360 12288
rect 13127 12257 13139 12260
rect 13081 12251 13139 12257
rect 13354 12248 13360 12260
rect 13412 12248 13418 12300
rect 13722 12288 13728 12300
rect 13683 12260 13728 12288
rect 13722 12248 13728 12260
rect 13780 12248 13786 12300
rect 13998 12248 14004 12300
rect 14056 12288 14062 12300
rect 14918 12288 14924 12300
rect 14056 12260 14924 12288
rect 14056 12248 14062 12260
rect 14918 12248 14924 12260
rect 14976 12288 14982 12300
rect 15749 12291 15807 12297
rect 15749 12288 15761 12291
rect 14976 12260 15761 12288
rect 14976 12248 14982 12260
rect 15749 12257 15761 12260
rect 15795 12257 15807 12291
rect 15749 12251 15807 12257
rect 7929 12223 7987 12229
rect 7929 12189 7941 12223
rect 7975 12189 7987 12223
rect 7929 12183 7987 12189
rect 8573 12223 8631 12229
rect 8573 12189 8585 12223
rect 8619 12189 8631 12223
rect 8573 12183 8631 12189
rect 7742 12152 7748 12164
rect 6656 12124 7748 12152
rect 1854 12044 1860 12096
rect 1912 12084 1918 12096
rect 2590 12084 2596 12096
rect 1912 12056 2596 12084
rect 1912 12044 1918 12056
rect 2590 12044 2596 12056
rect 2648 12084 2654 12096
rect 6656 12093 6684 12124
rect 7742 12112 7748 12124
rect 7800 12112 7806 12164
rect 8588 12152 8616 12183
rect 9030 12180 9036 12232
rect 9088 12220 9094 12232
rect 9217 12223 9275 12229
rect 9217 12220 9229 12223
rect 9088 12192 9229 12220
rect 9088 12180 9094 12192
rect 9217 12189 9229 12192
rect 9263 12189 9275 12223
rect 9217 12183 9275 12189
rect 9490 12180 9496 12232
rect 9548 12220 9554 12232
rect 9861 12223 9919 12229
rect 9861 12220 9873 12223
rect 9548 12192 9873 12220
rect 9548 12180 9554 12192
rect 9861 12189 9873 12192
rect 9907 12189 9919 12223
rect 10686 12220 10692 12232
rect 10647 12192 10692 12220
rect 9861 12183 9919 12189
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 11333 12223 11391 12229
rect 11333 12189 11345 12223
rect 11379 12220 11391 12223
rect 11698 12220 11704 12232
rect 11379 12192 11704 12220
rect 11379 12189 11391 12192
rect 11333 12183 11391 12189
rect 11698 12180 11704 12192
rect 11756 12180 11762 12232
rect 17512 12229 17540 12328
rect 18785 12325 18797 12359
rect 18831 12356 18843 12359
rect 18874 12356 18880 12368
rect 18831 12328 18880 12356
rect 18831 12325 18843 12328
rect 18785 12319 18843 12325
rect 18874 12316 18880 12328
rect 18932 12356 18938 12368
rect 19812 12356 19840 12396
rect 20346 12384 20352 12396
rect 20404 12384 20410 12436
rect 20438 12384 20444 12436
rect 20496 12424 20502 12436
rect 21637 12427 21695 12433
rect 21637 12424 21649 12427
rect 20496 12396 21649 12424
rect 20496 12384 20502 12396
rect 21637 12393 21649 12396
rect 21683 12393 21695 12427
rect 25774 12424 25780 12436
rect 21637 12387 21695 12393
rect 21744 12396 25780 12424
rect 18932 12328 19840 12356
rect 18932 12316 18938 12328
rect 20714 12316 20720 12368
rect 20772 12356 20778 12368
rect 21744 12356 21772 12396
rect 25774 12384 25780 12396
rect 25832 12384 25838 12436
rect 27614 12384 27620 12436
rect 27672 12424 27678 12436
rect 27709 12427 27767 12433
rect 27709 12424 27721 12427
rect 27672 12396 27721 12424
rect 27672 12384 27678 12396
rect 27709 12393 27721 12396
rect 27755 12393 27767 12427
rect 29822 12424 29828 12436
rect 29783 12396 29828 12424
rect 27709 12387 27767 12393
rect 29822 12384 29828 12396
rect 29880 12384 29886 12436
rect 30282 12384 30288 12436
rect 30340 12424 30346 12436
rect 38010 12424 38016 12436
rect 30340 12396 38016 12424
rect 30340 12384 30346 12396
rect 38010 12384 38016 12396
rect 38068 12384 38074 12436
rect 20772 12328 21772 12356
rect 22833 12359 22891 12365
rect 20772 12316 20778 12328
rect 22833 12325 22845 12359
rect 22879 12356 22891 12359
rect 23290 12356 23296 12368
rect 22879 12328 23296 12356
rect 22879 12325 22891 12328
rect 22833 12319 22891 12325
rect 23290 12316 23296 12328
rect 23348 12316 23354 12368
rect 23658 12316 23664 12368
rect 23716 12356 23722 12368
rect 24673 12359 24731 12365
rect 24673 12356 24685 12359
rect 23716 12328 24685 12356
rect 23716 12316 23722 12328
rect 24673 12325 24685 12328
rect 24719 12325 24731 12359
rect 27065 12359 27123 12365
rect 27065 12356 27077 12359
rect 24673 12319 24731 12325
rect 24780 12328 27077 12356
rect 18233 12291 18291 12297
rect 18233 12257 18245 12291
rect 18279 12288 18291 12291
rect 18966 12288 18972 12300
rect 18279 12260 18972 12288
rect 18279 12257 18291 12260
rect 18233 12251 18291 12257
rect 18966 12248 18972 12260
rect 19024 12248 19030 12300
rect 19242 12248 19248 12300
rect 19300 12288 19306 12300
rect 20165 12291 20223 12297
rect 20165 12288 20177 12291
rect 19300 12260 20177 12288
rect 19300 12248 19306 12260
rect 20165 12257 20177 12260
rect 20211 12288 20223 12291
rect 20254 12288 20260 12300
rect 20211 12260 20260 12288
rect 20211 12257 20223 12260
rect 20165 12251 20223 12257
rect 20254 12248 20260 12260
rect 20312 12248 20318 12300
rect 20346 12248 20352 12300
rect 20404 12288 20410 12300
rect 23382 12288 23388 12300
rect 20404 12260 22876 12288
rect 23343 12260 23388 12288
rect 20404 12248 20410 12260
rect 17497 12223 17555 12229
rect 17497 12189 17509 12223
rect 17543 12189 17555 12223
rect 19426 12220 19432 12232
rect 19387 12192 19432 12220
rect 17497 12183 17555 12189
rect 19426 12180 19432 12192
rect 19484 12180 19490 12232
rect 21358 12180 21364 12232
rect 21416 12220 21422 12232
rect 22097 12223 22155 12229
rect 22097 12220 22109 12223
rect 21416 12192 22109 12220
rect 21416 12180 21422 12192
rect 22097 12189 22109 12192
rect 22143 12189 22155 12223
rect 22278 12220 22284 12232
rect 22239 12192 22284 12220
rect 22097 12183 22155 12189
rect 22278 12180 22284 12192
rect 22336 12180 22342 12232
rect 8754 12152 8760 12164
rect 8588 12124 8760 12152
rect 8754 12112 8760 12124
rect 8812 12152 8818 12164
rect 9582 12152 9588 12164
rect 8812 12124 9588 12152
rect 8812 12112 8818 12124
rect 9582 12112 9588 12124
rect 9640 12112 9646 12164
rect 9953 12155 10011 12161
rect 9953 12121 9965 12155
rect 9999 12152 10011 12155
rect 9999 12124 11376 12152
rect 9999 12121 10011 12124
rect 9953 12115 10011 12121
rect 6641 12087 6699 12093
rect 6641 12084 6653 12087
rect 2648 12056 6653 12084
rect 2648 12044 2654 12056
rect 6641 12053 6653 12056
rect 6687 12053 6699 12087
rect 6641 12047 6699 12053
rect 8481 12087 8539 12093
rect 8481 12053 8493 12087
rect 8527 12084 8539 12087
rect 10410 12084 10416 12096
rect 8527 12056 10416 12084
rect 8527 12053 8539 12056
rect 8481 12047 8539 12053
rect 10410 12044 10416 12056
rect 10468 12044 10474 12096
rect 11348 12084 11376 12124
rect 11422 12112 11428 12164
rect 11480 12152 11486 12164
rect 11885 12155 11943 12161
rect 11885 12152 11897 12155
rect 11480 12124 11897 12152
rect 11480 12112 11486 12124
rect 11885 12121 11897 12124
rect 11931 12121 11943 12155
rect 11885 12115 11943 12121
rect 11974 12112 11980 12164
rect 12032 12152 12038 12164
rect 12032 12124 12077 12152
rect 12032 12112 12038 12124
rect 12526 12112 12532 12164
rect 12584 12152 12590 12164
rect 12710 12152 12716 12164
rect 12584 12124 12716 12152
rect 12584 12112 12590 12124
rect 12710 12112 12716 12124
rect 12768 12112 12774 12164
rect 13173 12155 13231 12161
rect 13173 12121 13185 12155
rect 13219 12121 13231 12155
rect 13173 12115 13231 12121
rect 13188 12084 13216 12115
rect 13722 12112 13728 12164
rect 13780 12152 13786 12164
rect 14553 12155 14611 12161
rect 14553 12152 14565 12155
rect 13780 12124 14565 12152
rect 13780 12112 13786 12124
rect 14553 12121 14565 12124
rect 14599 12121 14611 12155
rect 14553 12115 14611 12121
rect 15105 12155 15163 12161
rect 15105 12121 15117 12155
rect 15151 12121 15163 12155
rect 15105 12115 15163 12121
rect 15197 12155 15255 12161
rect 15197 12121 15209 12155
rect 15243 12152 15255 12155
rect 15562 12152 15568 12164
rect 15243 12124 15568 12152
rect 15243 12121 15255 12124
rect 15197 12115 15255 12121
rect 11348 12056 13216 12084
rect 13446 12044 13452 12096
rect 13504 12084 13510 12096
rect 15120 12084 15148 12115
rect 15562 12112 15568 12124
rect 15620 12112 15626 12164
rect 16666 12152 16672 12164
rect 16627 12124 16672 12152
rect 16666 12112 16672 12124
rect 16724 12112 16730 12164
rect 16761 12155 16819 12161
rect 16761 12121 16773 12155
rect 16807 12152 16819 12155
rect 17310 12152 17316 12164
rect 16807 12124 17316 12152
rect 16807 12121 16819 12124
rect 16761 12115 16819 12121
rect 17310 12112 17316 12124
rect 17368 12112 17374 12164
rect 18325 12155 18383 12161
rect 18325 12121 18337 12155
rect 18371 12152 18383 12155
rect 19334 12152 19340 12164
rect 18371 12124 19340 12152
rect 18371 12121 18383 12124
rect 18325 12115 18383 12121
rect 19334 12112 19340 12124
rect 19392 12112 19398 12164
rect 19702 12112 19708 12164
rect 19760 12152 19766 12164
rect 20257 12155 20315 12161
rect 20257 12152 20269 12155
rect 19760 12124 20269 12152
rect 19760 12112 19766 12124
rect 20257 12121 20269 12124
rect 20303 12121 20315 12155
rect 20257 12115 20315 12121
rect 21177 12155 21235 12161
rect 21177 12121 21189 12155
rect 21223 12152 21235 12155
rect 21726 12152 21732 12164
rect 21223 12124 21732 12152
rect 21223 12121 21235 12124
rect 21177 12115 21235 12121
rect 21726 12112 21732 12124
rect 21784 12112 21790 12164
rect 13504 12056 15148 12084
rect 17589 12087 17647 12093
rect 13504 12044 13510 12056
rect 17589 12053 17601 12087
rect 17635 12084 17647 12087
rect 19058 12084 19064 12096
rect 17635 12056 19064 12084
rect 17635 12053 17647 12056
rect 17589 12047 17647 12053
rect 19058 12044 19064 12056
rect 19116 12044 19122 12096
rect 19521 12087 19579 12093
rect 19521 12053 19533 12087
rect 19567 12084 19579 12087
rect 20806 12084 20812 12096
rect 19567 12056 20812 12084
rect 19567 12053 19579 12056
rect 19521 12047 19579 12053
rect 20806 12044 20812 12056
rect 20864 12044 20870 12096
rect 22848 12084 22876 12260
rect 23382 12248 23388 12260
rect 23440 12248 23446 12300
rect 23566 12248 23572 12300
rect 23624 12288 23630 12300
rect 24780 12288 24808 12328
rect 27065 12325 27077 12328
rect 27111 12325 27123 12359
rect 27065 12319 27123 12325
rect 27430 12316 27436 12368
rect 27488 12356 27494 12368
rect 29840 12356 29868 12384
rect 27488 12328 29868 12356
rect 27488 12316 27494 12328
rect 23624 12260 24808 12288
rect 23624 12248 23630 12260
rect 25130 12248 25136 12300
rect 25188 12288 25194 12300
rect 27890 12288 27896 12300
rect 25188 12260 27896 12288
rect 25188 12248 25194 12260
rect 27890 12248 27896 12260
rect 27948 12248 27954 12300
rect 26513 12223 26571 12229
rect 26513 12189 26525 12223
rect 26559 12220 26571 12223
rect 26602 12220 26608 12232
rect 26559 12192 26608 12220
rect 26559 12189 26571 12192
rect 26513 12183 26571 12189
rect 26602 12180 26608 12192
rect 26660 12180 26666 12232
rect 27157 12223 27215 12229
rect 27157 12189 27169 12223
rect 27203 12220 27215 12223
rect 27430 12220 27436 12232
rect 27203 12192 27436 12220
rect 27203 12189 27215 12192
rect 27157 12183 27215 12189
rect 27430 12180 27436 12192
rect 27488 12180 27494 12232
rect 27614 12180 27620 12232
rect 27672 12220 27678 12232
rect 27672 12192 27717 12220
rect 27672 12180 27678 12192
rect 27982 12180 27988 12232
rect 28040 12220 28046 12232
rect 28445 12223 28503 12229
rect 28445 12220 28457 12223
rect 28040 12192 28457 12220
rect 28040 12180 28046 12192
rect 28445 12189 28457 12192
rect 28491 12189 28503 12223
rect 28445 12183 28503 12189
rect 28902 12180 28908 12232
rect 28960 12220 28966 12232
rect 29089 12223 29147 12229
rect 29089 12220 29101 12223
rect 28960 12192 29101 12220
rect 28960 12180 28966 12192
rect 29089 12189 29101 12192
rect 29135 12220 29147 12223
rect 30285 12223 30343 12229
rect 30285 12220 30297 12223
rect 29135 12192 30297 12220
rect 29135 12189 29147 12192
rect 29089 12183 29147 12189
rect 30285 12189 30297 12192
rect 30331 12189 30343 12223
rect 30285 12183 30343 12189
rect 22922 12112 22928 12164
rect 22980 12152 22986 12164
rect 23198 12152 23204 12164
rect 22980 12124 23204 12152
rect 22980 12112 22986 12124
rect 23198 12112 23204 12124
rect 23256 12112 23262 12164
rect 23474 12152 23480 12164
rect 23435 12124 23480 12152
rect 23474 12112 23480 12124
rect 23532 12112 23538 12164
rect 23658 12112 23664 12164
rect 23716 12152 23722 12164
rect 24029 12155 24087 12161
rect 24029 12152 24041 12155
rect 23716 12124 24041 12152
rect 23716 12112 23722 12124
rect 24029 12121 24041 12124
rect 24075 12152 24087 12155
rect 24854 12152 24860 12164
rect 24075 12124 24860 12152
rect 24075 12121 24087 12124
rect 24029 12115 24087 12121
rect 24854 12112 24860 12124
rect 24912 12112 24918 12164
rect 25130 12152 25136 12164
rect 25091 12124 25136 12152
rect 25130 12112 25136 12124
rect 25188 12112 25194 12164
rect 25222 12112 25228 12164
rect 25280 12152 25286 12164
rect 25498 12152 25504 12164
rect 25280 12124 25504 12152
rect 25280 12112 25286 12124
rect 25498 12112 25504 12124
rect 25556 12112 25562 12164
rect 25869 12155 25927 12161
rect 25869 12121 25881 12155
rect 25915 12121 25927 12155
rect 25869 12115 25927 12121
rect 25961 12155 26019 12161
rect 25961 12121 25973 12155
rect 26007 12152 26019 12155
rect 28997 12155 29055 12161
rect 28997 12152 29009 12155
rect 26007 12124 29009 12152
rect 26007 12121 26019 12124
rect 25961 12115 26019 12121
rect 28997 12121 29009 12124
rect 29043 12121 29055 12155
rect 28997 12115 29055 12121
rect 25884 12084 25912 12115
rect 28350 12084 28356 12096
rect 22848 12056 25912 12084
rect 28311 12056 28356 12084
rect 28350 12044 28356 12056
rect 28408 12044 28414 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 7929 11883 7987 11889
rect 7929 11849 7941 11883
rect 7975 11880 7987 11883
rect 9030 11880 9036 11892
rect 7975 11852 9036 11880
rect 7975 11849 7987 11852
rect 7929 11843 7987 11849
rect 9030 11840 9036 11852
rect 9088 11840 9094 11892
rect 10318 11840 10324 11892
rect 10376 11880 10382 11892
rect 10413 11883 10471 11889
rect 10413 11880 10425 11883
rect 10376 11852 10425 11880
rect 10376 11840 10382 11852
rect 10413 11849 10425 11852
rect 10459 11849 10471 11883
rect 10413 11843 10471 11849
rect 11057 11883 11115 11889
rect 11057 11849 11069 11883
rect 11103 11880 11115 11883
rect 11146 11880 11152 11892
rect 11103 11852 11152 11880
rect 11103 11849 11115 11852
rect 11057 11843 11115 11849
rect 11146 11840 11152 11852
rect 11204 11840 11210 11892
rect 12161 11883 12219 11889
rect 12161 11849 12173 11883
rect 12207 11880 12219 11883
rect 12207 11852 15700 11880
rect 12207 11849 12219 11852
rect 12161 11843 12219 11849
rect 9861 11815 9919 11821
rect 9861 11781 9873 11815
rect 9907 11812 9919 11815
rect 12250 11812 12256 11824
rect 9907 11784 12256 11812
rect 9907 11781 9919 11784
rect 9861 11775 9919 11781
rect 12250 11772 12256 11784
rect 12308 11772 12314 11824
rect 12526 11772 12532 11824
rect 12584 11812 12590 11824
rect 12805 11815 12863 11821
rect 12805 11812 12817 11815
rect 12584 11784 12817 11812
rect 12584 11772 12590 11784
rect 12805 11781 12817 11784
rect 12851 11781 12863 11815
rect 12805 11775 12863 11781
rect 12894 11772 12900 11824
rect 12952 11812 12958 11824
rect 13357 11815 13415 11821
rect 13357 11812 13369 11815
rect 12952 11784 13369 11812
rect 12952 11772 12958 11784
rect 13357 11781 13369 11784
rect 13403 11812 13415 11815
rect 13722 11812 13728 11824
rect 13403 11784 13728 11812
rect 13403 11781 13415 11784
rect 13357 11775 13415 11781
rect 13722 11772 13728 11784
rect 13780 11772 13786 11824
rect 13906 11772 13912 11824
rect 13964 11812 13970 11824
rect 14001 11815 14059 11821
rect 14001 11812 14013 11815
rect 13964 11784 14013 11812
rect 13964 11772 13970 11784
rect 14001 11781 14013 11784
rect 14047 11781 14059 11815
rect 14918 11812 14924 11824
rect 14879 11784 14924 11812
rect 14001 11775 14059 11781
rect 14918 11772 14924 11784
rect 14976 11772 14982 11824
rect 15672 11821 15700 11852
rect 17310 11840 17316 11892
rect 17368 11880 17374 11892
rect 23658 11880 23664 11892
rect 17368 11852 23664 11880
rect 17368 11840 17374 11852
rect 23658 11840 23664 11852
rect 23716 11840 23722 11892
rect 28537 11883 28595 11889
rect 28537 11880 28549 11883
rect 23860 11852 28549 11880
rect 15657 11815 15715 11821
rect 15657 11781 15669 11815
rect 15703 11781 15715 11815
rect 15657 11775 15715 11781
rect 15749 11815 15807 11821
rect 15749 11781 15761 11815
rect 15795 11812 15807 11815
rect 18230 11812 18236 11824
rect 15795 11784 17724 11812
rect 18191 11784 18236 11812
rect 15795 11781 15807 11784
rect 15749 11775 15807 11781
rect 8110 11704 8116 11756
rect 8168 11744 8174 11756
rect 8389 11747 8447 11753
rect 8389 11744 8401 11747
rect 8168 11716 8401 11744
rect 8168 11704 8174 11716
rect 8389 11713 8401 11716
rect 8435 11713 8447 11747
rect 8389 11707 8447 11713
rect 9033 11747 9091 11753
rect 9033 11713 9045 11747
rect 9079 11713 9091 11747
rect 10502 11744 10508 11756
rect 10463 11716 10508 11744
rect 9033 11707 9091 11713
rect 9048 11676 9076 11707
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 10962 11744 10968 11756
rect 10704 11716 10968 11744
rect 10704 11676 10732 11716
rect 10962 11704 10968 11716
rect 11020 11704 11026 11756
rect 11146 11744 11152 11756
rect 11107 11716 11152 11744
rect 11146 11704 11152 11716
rect 11204 11704 11210 11756
rect 16298 11704 16304 11756
rect 16356 11744 16362 11756
rect 17034 11744 17040 11756
rect 16356 11716 16401 11744
rect 16995 11716 17040 11744
rect 16356 11704 16362 11716
rect 17034 11704 17040 11716
rect 17092 11704 17098 11756
rect 12713 11679 12771 11685
rect 7300 11648 10732 11676
rect 10796 11648 12664 11676
rect 7300 11552 7328 11648
rect 8481 11611 8539 11617
rect 8481 11577 8493 11611
rect 8527 11608 8539 11611
rect 10796 11608 10824 11648
rect 8527 11580 10824 11608
rect 8527 11577 8539 11580
rect 8481 11571 8539 11577
rect 11054 11568 11060 11620
rect 11112 11608 11118 11620
rect 11238 11608 11244 11620
rect 11112 11580 11244 11608
rect 11112 11568 11118 11580
rect 11238 11568 11244 11580
rect 11296 11568 11302 11620
rect 11330 11568 11336 11620
rect 11388 11608 11394 11620
rect 12434 11608 12440 11620
rect 11388 11580 12440 11608
rect 11388 11568 11394 11580
rect 12434 11568 12440 11580
rect 12492 11568 12498 11620
rect 12636 11608 12664 11648
rect 12713 11645 12725 11679
rect 12759 11676 12771 11679
rect 13170 11676 13176 11688
rect 12759 11648 13176 11676
rect 12759 11645 12771 11648
rect 12713 11639 12771 11645
rect 13170 11636 13176 11648
rect 13228 11636 13234 11688
rect 13909 11679 13967 11685
rect 13909 11645 13921 11679
rect 13955 11676 13967 11679
rect 13998 11676 14004 11688
rect 13955 11648 14004 11676
rect 13955 11645 13967 11648
rect 13909 11639 13967 11645
rect 13998 11636 14004 11648
rect 14056 11676 14062 11688
rect 17586 11676 17592 11688
rect 14056 11648 17592 11676
rect 14056 11636 14062 11648
rect 17586 11636 17592 11648
rect 17644 11636 17650 11688
rect 15470 11608 15476 11620
rect 12636 11580 15476 11608
rect 15470 11568 15476 11580
rect 15528 11568 15534 11620
rect 17696 11608 17724 11784
rect 18230 11772 18236 11784
rect 18288 11772 18294 11824
rect 19058 11812 19064 11824
rect 19019 11784 19064 11812
rect 19058 11772 19064 11784
rect 19116 11772 19122 11824
rect 20162 11772 20168 11824
rect 20220 11812 20226 11824
rect 20257 11815 20315 11821
rect 20257 11812 20269 11815
rect 20220 11784 20269 11812
rect 20220 11772 20226 11784
rect 20257 11781 20269 11784
rect 20303 11781 20315 11815
rect 20257 11775 20315 11781
rect 20806 11772 20812 11824
rect 20864 11812 20870 11824
rect 22189 11815 22247 11821
rect 22189 11812 22201 11815
rect 20864 11784 22201 11812
rect 20864 11772 20870 11784
rect 22189 11781 22201 11784
rect 22235 11781 22247 11815
rect 22189 11775 22247 11781
rect 22370 11772 22376 11824
rect 22428 11812 22434 11824
rect 22428 11784 22784 11812
rect 22428 11772 22434 11784
rect 21358 11744 21364 11756
rect 21319 11716 21364 11744
rect 21358 11704 21364 11716
rect 21416 11704 21422 11756
rect 21453 11747 21511 11753
rect 21453 11713 21465 11747
rect 21499 11744 21511 11747
rect 21542 11744 21548 11756
rect 21499 11716 21548 11744
rect 21499 11713 21511 11716
rect 21453 11707 21511 11713
rect 21542 11704 21548 11716
rect 21600 11744 21606 11756
rect 21818 11744 21824 11756
rect 21600 11716 21824 11744
rect 21600 11704 21606 11716
rect 21818 11704 21824 11716
rect 21876 11704 21882 11756
rect 22756 11753 22784 11784
rect 23014 11772 23020 11824
rect 23072 11812 23078 11824
rect 23860 11821 23888 11852
rect 28537 11849 28549 11852
rect 28583 11849 28595 11883
rect 28537 11843 28595 11849
rect 23293 11815 23351 11821
rect 23293 11812 23305 11815
rect 23072 11784 23305 11812
rect 23072 11772 23078 11784
rect 23293 11781 23305 11784
rect 23339 11781 23351 11815
rect 23293 11775 23351 11781
rect 23845 11815 23903 11821
rect 23845 11781 23857 11815
rect 23891 11781 23903 11815
rect 23845 11775 23903 11781
rect 23934 11772 23940 11824
rect 23992 11812 23998 11824
rect 24578 11812 24584 11824
rect 23992 11784 24584 11812
rect 23992 11772 23998 11784
rect 24578 11772 24584 11784
rect 24636 11772 24642 11824
rect 24854 11812 24860 11824
rect 24815 11784 24860 11812
rect 24854 11772 24860 11784
rect 24912 11772 24918 11824
rect 25409 11815 25467 11821
rect 25409 11781 25421 11815
rect 25455 11812 25467 11815
rect 26145 11815 26203 11821
rect 26145 11812 26157 11815
rect 25455 11784 26157 11812
rect 25455 11781 25467 11784
rect 25409 11775 25467 11781
rect 26145 11781 26157 11784
rect 26191 11781 26203 11815
rect 26145 11775 26203 11781
rect 26326 11772 26332 11824
rect 26384 11812 26390 11824
rect 27890 11812 27896 11824
rect 26384 11784 27896 11812
rect 26384 11772 26390 11784
rect 27890 11772 27896 11784
rect 27948 11772 27954 11824
rect 22741 11747 22799 11753
rect 22741 11713 22753 11747
rect 22787 11744 22799 11747
rect 23198 11744 23204 11756
rect 22787 11716 23204 11744
rect 22787 11713 22799 11716
rect 22741 11707 22799 11713
rect 23198 11704 23204 11716
rect 23256 11704 23262 11756
rect 26237 11747 26295 11753
rect 26237 11713 26249 11747
rect 26283 11713 26295 11747
rect 27338 11744 27344 11756
rect 27299 11716 27344 11744
rect 26237 11707 26295 11713
rect 17862 11676 17868 11688
rect 17823 11648 17868 11676
rect 17862 11636 17868 11648
rect 17920 11636 17926 11688
rect 18325 11679 18383 11685
rect 18325 11645 18337 11679
rect 18371 11676 18383 11679
rect 18690 11676 18696 11688
rect 18371 11648 18696 11676
rect 18371 11645 18383 11648
rect 18325 11639 18383 11645
rect 18690 11636 18696 11648
rect 18748 11636 18754 11688
rect 18966 11676 18972 11688
rect 18927 11648 18972 11676
rect 18966 11636 18972 11648
rect 19024 11636 19030 11688
rect 19978 11636 19984 11688
rect 20036 11676 20042 11688
rect 20165 11679 20223 11685
rect 20165 11676 20177 11679
rect 20036 11648 20177 11676
rect 20036 11636 20042 11648
rect 20165 11645 20177 11648
rect 20211 11645 20223 11679
rect 20165 11639 20223 11645
rect 20441 11679 20499 11685
rect 20441 11645 20453 11679
rect 20487 11645 20499 11679
rect 20441 11639 20499 11645
rect 19150 11608 19156 11620
rect 17696 11580 19156 11608
rect 19150 11568 19156 11580
rect 19208 11568 19214 11620
rect 19521 11611 19579 11617
rect 19521 11577 19533 11611
rect 19567 11608 19579 11611
rect 20456 11608 20484 11639
rect 22094 11636 22100 11688
rect 22152 11676 22158 11688
rect 23566 11676 23572 11688
rect 22152 11648 23572 11676
rect 22152 11636 22158 11648
rect 23566 11636 23572 11648
rect 23624 11636 23630 11688
rect 23937 11679 23995 11685
rect 23937 11645 23949 11679
rect 23983 11676 23995 11679
rect 25222 11676 25228 11688
rect 23983 11648 25228 11676
rect 23983 11645 23995 11648
rect 23937 11639 23995 11645
rect 25222 11636 25228 11648
rect 25280 11636 25286 11688
rect 25498 11676 25504 11688
rect 25459 11648 25504 11676
rect 25498 11636 25504 11648
rect 25556 11636 25562 11688
rect 26252 11676 26280 11707
rect 27338 11704 27344 11716
rect 27396 11704 27402 11756
rect 27430 11704 27436 11756
rect 27488 11744 27494 11756
rect 27801 11747 27859 11753
rect 27801 11744 27813 11747
rect 27488 11716 27813 11744
rect 27488 11704 27494 11716
rect 27801 11713 27813 11716
rect 27847 11713 27859 11747
rect 28442 11744 28448 11756
rect 28403 11716 28448 11744
rect 27801 11707 27859 11713
rect 28442 11704 28448 11716
rect 28500 11704 28506 11756
rect 37553 11747 37611 11753
rect 37553 11713 37565 11747
rect 37599 11744 37611 11747
rect 38194 11744 38200 11756
rect 37599 11716 38200 11744
rect 37599 11713 37611 11716
rect 37553 11707 37611 11713
rect 38194 11704 38200 11716
rect 38252 11704 38258 11756
rect 29089 11679 29147 11685
rect 29089 11676 29101 11679
rect 25608 11648 29101 11676
rect 22554 11608 22560 11620
rect 19567 11580 22560 11608
rect 19567 11577 19579 11580
rect 19521 11571 19579 11577
rect 22554 11568 22560 11580
rect 22612 11568 22618 11620
rect 23382 11568 23388 11620
rect 23440 11608 23446 11620
rect 25608 11608 25636 11648
rect 29089 11645 29101 11648
rect 29135 11645 29147 11679
rect 29089 11639 29147 11645
rect 27893 11611 27951 11617
rect 27893 11608 27905 11611
rect 23440 11580 25636 11608
rect 25700 11580 27905 11608
rect 23440 11568 23446 11580
rect 7282 11540 7288 11552
rect 7243 11512 7288 11540
rect 7282 11500 7288 11512
rect 7340 11500 7346 11552
rect 9122 11540 9128 11552
rect 9083 11512 9128 11540
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 10410 11500 10416 11552
rect 10468 11540 10474 11552
rect 13354 11540 13360 11552
rect 10468 11512 13360 11540
rect 10468 11500 10474 11512
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 17129 11543 17187 11549
rect 17129 11509 17141 11543
rect 17175 11540 17187 11543
rect 20714 11540 20720 11552
rect 17175 11512 20720 11540
rect 17175 11509 17187 11512
rect 17129 11503 17187 11509
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 23474 11500 23480 11552
rect 23532 11540 23538 11552
rect 25700 11540 25728 11580
rect 27893 11577 27905 11580
rect 27939 11577 27951 11611
rect 27893 11571 27951 11577
rect 30742 11568 30748 11620
rect 30800 11608 30806 11620
rect 38013 11611 38071 11617
rect 38013 11608 38025 11611
rect 30800 11580 38025 11608
rect 30800 11568 30806 11580
rect 38013 11577 38025 11580
rect 38059 11577 38071 11611
rect 38013 11571 38071 11577
rect 23532 11512 25728 11540
rect 23532 11500 23538 11512
rect 25866 11500 25872 11552
rect 25924 11540 25930 11552
rect 27062 11540 27068 11552
rect 25924 11512 27068 11540
rect 25924 11500 25930 11512
rect 27062 11500 27068 11512
rect 27120 11500 27126 11552
rect 27246 11540 27252 11552
rect 27207 11512 27252 11540
rect 27246 11500 27252 11512
rect 27304 11500 27310 11552
rect 27522 11500 27528 11552
rect 27580 11540 27586 11552
rect 29641 11543 29699 11549
rect 29641 11540 29653 11543
rect 27580 11512 29653 11540
rect 27580 11500 27586 11512
rect 29641 11509 29653 11512
rect 29687 11509 29699 11543
rect 29641 11503 29699 11509
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 11241 11339 11299 11345
rect 11241 11305 11253 11339
rect 11287 11336 11299 11339
rect 13446 11336 13452 11348
rect 11287 11308 13452 11336
rect 11287 11305 11299 11308
rect 11241 11299 11299 11305
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 13630 11296 13636 11348
rect 13688 11336 13694 11348
rect 14277 11339 14335 11345
rect 14277 11336 14289 11339
rect 13688 11308 14289 11336
rect 13688 11296 13694 11308
rect 14277 11305 14289 11308
rect 14323 11305 14335 11339
rect 14277 11299 14335 11305
rect 15562 11296 15568 11348
rect 15620 11336 15626 11348
rect 15620 11308 19840 11336
rect 15620 11296 15626 11308
rect 11606 11268 11612 11280
rect 9140 11240 11612 11268
rect 9140 11141 9168 11240
rect 11606 11228 11612 11240
rect 11664 11228 11670 11280
rect 15010 11268 15016 11280
rect 12176 11240 15016 11268
rect 12176 11209 12204 11240
rect 15010 11228 15016 11240
rect 15068 11228 15074 11280
rect 16206 11268 16212 11280
rect 15120 11240 16212 11268
rect 10413 11203 10471 11209
rect 10413 11169 10425 11203
rect 10459 11200 10471 11203
rect 12161 11203 12219 11209
rect 12161 11200 12173 11203
rect 10459 11172 12173 11200
rect 10459 11169 10471 11172
rect 10413 11163 10471 11169
rect 12161 11169 12173 11172
rect 12207 11169 12219 11203
rect 12161 11163 12219 11169
rect 12250 11160 12256 11212
rect 12308 11200 12314 11212
rect 13081 11203 13139 11209
rect 13081 11200 13093 11203
rect 12308 11172 13093 11200
rect 12308 11160 12314 11172
rect 13081 11169 13093 11172
rect 13127 11169 13139 11203
rect 13081 11163 13139 11169
rect 13538 11160 13544 11212
rect 13596 11200 13602 11212
rect 14737 11203 14795 11209
rect 14737 11200 14749 11203
rect 13596 11172 14749 11200
rect 13596 11160 13602 11172
rect 14737 11169 14749 11172
rect 14783 11169 14795 11203
rect 14737 11163 14795 11169
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11132 8079 11135
rect 9125 11135 9183 11141
rect 9125 11132 9137 11135
rect 8067 11104 9137 11132
rect 8067 11101 8079 11104
rect 8021 11095 8079 11101
rect 9125 11101 9137 11104
rect 9171 11101 9183 11135
rect 11330 11132 11336 11144
rect 11291 11104 11336 11132
rect 9125 11095 9183 11101
rect 11330 11092 11336 11104
rect 11388 11092 11394 11144
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11132 13783 11135
rect 13998 11132 14004 11144
rect 13771 11104 14004 11132
rect 13771 11101 13783 11104
rect 13725 11095 13783 11101
rect 13998 11092 14004 11104
rect 14056 11092 14062 11144
rect 14918 11132 14924 11144
rect 14879 11104 14924 11132
rect 14918 11092 14924 11104
rect 14976 11092 14982 11144
rect 2866 11024 2872 11076
rect 2924 11064 2930 11076
rect 7834 11064 7840 11076
rect 2924 11036 7840 11064
rect 2924 11024 2930 11036
rect 7834 11024 7840 11036
rect 7892 11024 7898 11076
rect 8570 11064 8576 11076
rect 8531 11036 8576 11064
rect 8570 11024 8576 11036
rect 8628 11064 8634 11076
rect 9490 11064 9496 11076
rect 8628 11036 9496 11064
rect 8628 11024 8634 11036
rect 9490 11024 9496 11036
rect 9548 11024 9554 11076
rect 9766 11064 9772 11076
rect 9727 11036 9772 11064
rect 9766 11024 9772 11036
rect 9824 11024 9830 11076
rect 10318 11064 10324 11076
rect 10279 11036 10324 11064
rect 10318 11024 10324 11036
rect 10376 11024 10382 11076
rect 10410 11024 10416 11076
rect 10468 11064 10474 11076
rect 11422 11064 11428 11076
rect 10468 11036 11428 11064
rect 10468 11024 10474 11036
rect 11422 11024 11428 11036
rect 11480 11024 11486 11076
rect 11514 11024 11520 11076
rect 11572 11064 11578 11076
rect 11885 11067 11943 11073
rect 11885 11064 11897 11067
rect 11572 11036 11897 11064
rect 11572 11024 11578 11036
rect 11885 11033 11897 11036
rect 11931 11033 11943 11067
rect 11885 11027 11943 11033
rect 11977 11067 12035 11073
rect 11977 11033 11989 11067
rect 12023 11033 12035 11067
rect 11977 11027 12035 11033
rect 9214 10996 9220 11008
rect 9175 10968 9220 10996
rect 9214 10956 9220 10968
rect 9272 10956 9278 11008
rect 9858 10956 9864 11008
rect 9916 10996 9922 11008
rect 11992 10996 12020 11027
rect 13170 11024 13176 11076
rect 13228 11064 13234 11076
rect 13228 11036 13273 11064
rect 13228 11024 13234 11036
rect 13446 11024 13452 11076
rect 13504 11064 13510 11076
rect 15120 11064 15148 11240
rect 16206 11228 16212 11240
rect 16264 11268 16270 11280
rect 16669 11271 16727 11277
rect 16669 11268 16681 11271
rect 16264 11240 16681 11268
rect 16264 11228 16270 11240
rect 16669 11237 16681 11240
rect 16715 11237 16727 11271
rect 16669 11231 16727 11237
rect 19150 11228 19156 11280
rect 19208 11268 19214 11280
rect 19426 11268 19432 11280
rect 19208 11240 19432 11268
rect 19208 11228 19214 11240
rect 19426 11228 19432 11240
rect 19484 11228 19490 11280
rect 19812 11268 19840 11308
rect 19886 11296 19892 11348
rect 19944 11336 19950 11348
rect 21266 11336 21272 11348
rect 19944 11308 21272 11336
rect 19944 11296 19950 11308
rect 21266 11296 21272 11308
rect 21324 11296 21330 11348
rect 21358 11296 21364 11348
rect 21416 11336 21422 11348
rect 27246 11336 27252 11348
rect 21416 11308 27252 11336
rect 21416 11296 21422 11308
rect 27246 11296 27252 11308
rect 27304 11296 27310 11348
rect 20622 11268 20628 11280
rect 19812 11240 20628 11268
rect 20622 11228 20628 11240
rect 20680 11228 20686 11280
rect 21177 11271 21235 11277
rect 21177 11237 21189 11271
rect 21223 11268 21235 11271
rect 22370 11268 22376 11280
rect 21223 11240 22376 11268
rect 21223 11237 21235 11240
rect 21177 11231 21235 11237
rect 22370 11228 22376 11240
rect 22428 11228 22434 11280
rect 22554 11228 22560 11280
rect 22612 11268 22618 11280
rect 24670 11268 24676 11280
rect 22612 11240 24676 11268
rect 22612 11228 22618 11240
rect 24670 11228 24676 11240
rect 24728 11228 24734 11280
rect 28350 11268 28356 11280
rect 25700 11240 28356 11268
rect 15470 11200 15476 11212
rect 15431 11172 15476 11200
rect 15470 11160 15476 11172
rect 15528 11160 15534 11212
rect 16117 11203 16175 11209
rect 16117 11169 16129 11203
rect 16163 11200 16175 11203
rect 19242 11200 19248 11212
rect 16163 11172 19248 11200
rect 16163 11169 16175 11172
rect 16117 11163 16175 11169
rect 19242 11160 19248 11172
rect 19300 11160 19306 11212
rect 19886 11200 19892 11212
rect 19847 11172 19892 11200
rect 19886 11160 19892 11172
rect 19944 11160 19950 11212
rect 20073 11203 20131 11209
rect 20073 11169 20085 11203
rect 20119 11200 20131 11203
rect 21821 11203 21879 11209
rect 21821 11200 21833 11203
rect 20119 11172 21833 11200
rect 20119 11169 20131 11172
rect 20073 11163 20131 11169
rect 21821 11169 21833 11172
rect 21867 11200 21879 11203
rect 22094 11200 22100 11212
rect 21867 11172 22100 11200
rect 21867 11169 21879 11172
rect 21821 11163 21879 11169
rect 22094 11160 22100 11172
rect 22152 11160 22158 11212
rect 22278 11160 22284 11212
rect 22336 11200 22342 11212
rect 23569 11203 23627 11209
rect 23569 11200 23581 11203
rect 22336 11172 23581 11200
rect 22336 11160 22342 11172
rect 23569 11169 23581 11172
rect 23615 11200 23627 11203
rect 24578 11200 24584 11212
rect 23615 11172 24584 11200
rect 23615 11169 23627 11172
rect 23569 11163 23627 11169
rect 24578 11160 24584 11172
rect 24636 11200 24642 11212
rect 25225 11203 25283 11209
rect 25225 11200 25237 11203
rect 24636 11172 25237 11200
rect 24636 11160 24642 11172
rect 25225 11169 25237 11172
rect 25271 11169 25283 11203
rect 25225 11163 25283 11169
rect 18417 11135 18475 11141
rect 18417 11101 18429 11135
rect 18463 11132 18475 11135
rect 18506 11132 18512 11144
rect 18463 11104 18512 11132
rect 18463 11101 18475 11104
rect 18417 11095 18475 11101
rect 18506 11092 18512 11104
rect 18564 11092 18570 11144
rect 19429 11135 19487 11141
rect 19429 11101 19441 11135
rect 19475 11132 19487 11135
rect 20438 11132 20444 11144
rect 19475 11104 20444 11132
rect 19475 11101 19487 11104
rect 19429 11095 19487 11101
rect 20438 11092 20444 11104
rect 20496 11092 20502 11144
rect 15562 11064 15568 11076
rect 13504 11036 15148 11064
rect 15523 11036 15568 11064
rect 13504 11024 13510 11036
rect 15562 11024 15568 11036
rect 15620 11024 15626 11076
rect 18138 11064 18144 11076
rect 17710 11036 18000 11064
rect 18051 11036 18144 11064
rect 9916 10968 12020 10996
rect 9916 10956 9922 10968
rect 12710 10956 12716 11008
rect 12768 10996 12774 11008
rect 13814 10996 13820 11008
rect 12768 10968 13820 10996
rect 12768 10956 12774 10968
rect 13814 10956 13820 10968
rect 13872 10956 13878 11008
rect 17972 10996 18000 11036
rect 18138 11024 18144 11036
rect 18196 11024 18202 11076
rect 18690 11024 18696 11076
rect 18748 11064 18754 11076
rect 20625 11067 20683 11073
rect 20625 11064 20637 11067
rect 18748 11036 20637 11064
rect 18748 11024 18754 11036
rect 20625 11033 20637 11036
rect 20671 11033 20683 11067
rect 20625 11027 20683 11033
rect 18046 10996 18052 11008
rect 17972 10968 18052 10996
rect 18046 10956 18052 10968
rect 18104 10956 18110 11008
rect 18156 10996 18184 11024
rect 19058 10996 19064 11008
rect 18156 10968 19064 10996
rect 19058 10956 19064 10968
rect 19116 10956 19122 11008
rect 19518 10956 19524 11008
rect 19576 10996 19582 11008
rect 20070 10996 20076 11008
rect 19576 10968 20076 10996
rect 19576 10956 19582 10968
rect 20070 10956 20076 10968
rect 20128 10956 20134 11008
rect 20640 10996 20668 11027
rect 20714 11024 20720 11076
rect 20772 11064 20778 11076
rect 20772 11036 20817 11064
rect 20772 11024 20778 11036
rect 21266 11024 21272 11076
rect 21324 11064 21330 11076
rect 21324 11036 21496 11064
rect 21324 11024 21330 11036
rect 20898 10996 20904 11008
rect 20640 10968 20904 10996
rect 20898 10956 20904 10968
rect 20956 10996 20962 11008
rect 21358 10996 21364 11008
rect 20956 10968 21364 10996
rect 20956 10956 20962 10968
rect 21358 10956 21364 10968
rect 21416 10956 21422 11008
rect 21468 10996 21496 11036
rect 21910 11024 21916 11076
rect 21968 11064 21974 11076
rect 21968 11036 22013 11064
rect 21968 11024 21974 11036
rect 22278 11024 22284 11076
rect 22336 11064 22342 11076
rect 22465 11067 22523 11073
rect 22465 11064 22477 11067
rect 22336 11036 22477 11064
rect 22336 11024 22342 11036
rect 22465 11033 22477 11036
rect 22511 11064 22523 11067
rect 22925 11067 22983 11073
rect 22925 11064 22937 11067
rect 22511 11036 22937 11064
rect 22511 11033 22523 11036
rect 22465 11027 22523 11033
rect 22925 11033 22937 11036
rect 22971 11033 22983 11067
rect 23474 11064 23480 11076
rect 23435 11036 23480 11064
rect 22925 11027 22983 11033
rect 23474 11024 23480 11036
rect 23532 11024 23538 11076
rect 25133 11067 25191 11073
rect 25133 11033 25145 11067
rect 25179 11033 25191 11067
rect 25700 11064 25728 11240
rect 28350 11228 28356 11240
rect 28408 11228 28414 11280
rect 25774 11160 25780 11212
rect 25832 11200 25838 11212
rect 26418 11200 26424 11212
rect 25832 11172 25877 11200
rect 26379 11172 26424 11200
rect 25832 11160 25838 11172
rect 26418 11160 26424 11172
rect 26476 11160 26482 11212
rect 26602 11160 26608 11212
rect 26660 11200 26666 11212
rect 27341 11203 27399 11209
rect 27341 11200 27353 11203
rect 26660 11172 27353 11200
rect 26660 11160 26666 11172
rect 27341 11169 27353 11172
rect 27387 11169 27399 11203
rect 27341 11163 27399 11169
rect 27982 11092 27988 11144
rect 28040 11132 28046 11144
rect 28353 11135 28411 11141
rect 28353 11132 28365 11135
rect 28040 11104 28365 11132
rect 28040 11092 28046 11104
rect 28353 11101 28365 11104
rect 28399 11132 28411 11135
rect 28813 11135 28871 11141
rect 28813 11132 28825 11135
rect 28399 11104 28825 11132
rect 28399 11101 28411 11104
rect 28353 11095 28411 11101
rect 28813 11101 28825 11104
rect 28859 11132 28871 11135
rect 29733 11135 29791 11141
rect 29733 11132 29745 11135
rect 28859 11104 29745 11132
rect 28859 11101 28871 11104
rect 28813 11095 28871 11101
rect 29733 11101 29745 11104
rect 29779 11101 29791 11135
rect 29733 11095 29791 11101
rect 25133 11027 25191 11033
rect 25332 11036 25728 11064
rect 23382 10996 23388 11008
rect 21468 10968 23388 10996
rect 23382 10956 23388 10968
rect 23440 10956 23446 11008
rect 25148 10996 25176 11027
rect 25332 10996 25360 11036
rect 26142 11024 26148 11076
rect 26200 11024 26206 11076
rect 26326 11064 26332 11076
rect 26287 11036 26332 11064
rect 26326 11024 26332 11036
rect 26384 11024 26390 11076
rect 27065 11067 27123 11073
rect 27065 11064 27077 11067
rect 26528 11036 27077 11064
rect 25148 10968 25360 10996
rect 26160 10996 26188 11024
rect 26528 10996 26556 11036
rect 27065 11033 27077 11036
rect 27111 11033 27123 11067
rect 27065 11027 27123 11033
rect 27157 11067 27215 11073
rect 27157 11033 27169 11067
rect 27203 11064 27215 11067
rect 27203 11036 27660 11064
rect 27203 11033 27215 11036
rect 27157 11027 27215 11033
rect 27632 11008 27660 11036
rect 26160 10968 26556 10996
rect 27614 10956 27620 11008
rect 27672 10956 27678 11008
rect 28258 10996 28264 11008
rect 28219 10968 28264 10996
rect 28258 10956 28264 10968
rect 28316 10956 28322 11008
rect 30190 10956 30196 11008
rect 30248 10996 30254 11008
rect 34790 10996 34796 11008
rect 30248 10968 34796 10996
rect 30248 10956 30254 10968
rect 34790 10956 34796 10968
rect 34848 10956 34854 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 8754 10792 8760 10804
rect 8715 10764 8760 10792
rect 8754 10752 8760 10764
rect 8812 10752 8818 10804
rect 9214 10752 9220 10804
rect 9272 10792 9278 10804
rect 9272 10764 14596 10792
rect 9272 10752 9278 10764
rect 10413 10727 10471 10733
rect 10413 10693 10425 10727
rect 10459 10724 10471 10727
rect 12250 10724 12256 10736
rect 10459 10696 12256 10724
rect 10459 10693 10471 10696
rect 10413 10687 10471 10693
rect 12250 10684 12256 10696
rect 12308 10684 12314 10736
rect 12529 10727 12587 10733
rect 12529 10693 12541 10727
rect 12575 10724 12587 10727
rect 13078 10724 13084 10736
rect 12575 10696 13084 10724
rect 12575 10693 12587 10696
rect 12529 10687 12587 10693
rect 13078 10684 13084 10696
rect 13136 10684 13142 10736
rect 13262 10684 13268 10736
rect 13320 10724 13326 10736
rect 13357 10727 13415 10733
rect 13357 10724 13369 10727
rect 13320 10696 13369 10724
rect 13320 10684 13326 10696
rect 13357 10693 13369 10696
rect 13403 10693 13415 10727
rect 13357 10687 13415 10693
rect 13909 10727 13967 10733
rect 13909 10693 13921 10727
rect 13955 10724 13967 10727
rect 13998 10724 14004 10736
rect 13955 10696 14004 10724
rect 13955 10693 13967 10696
rect 13909 10687 13967 10693
rect 13998 10684 14004 10696
rect 14056 10684 14062 10736
rect 14568 10733 14596 10764
rect 14734 10752 14740 10804
rect 14792 10792 14798 10804
rect 18506 10792 18512 10804
rect 14792 10764 16988 10792
rect 14792 10752 14798 10764
rect 14553 10727 14611 10733
rect 14553 10693 14565 10727
rect 14599 10693 14611 10727
rect 14553 10687 14611 10693
rect 14642 10684 14648 10736
rect 14700 10724 14706 10736
rect 15749 10727 15807 10733
rect 15749 10724 15761 10727
rect 14700 10696 15761 10724
rect 14700 10684 14706 10696
rect 15749 10693 15761 10696
rect 15795 10693 15807 10727
rect 15749 10687 15807 10693
rect 16301 10727 16359 10733
rect 16301 10693 16313 10727
rect 16347 10724 16359 10727
rect 16574 10724 16580 10736
rect 16347 10696 16580 10724
rect 16347 10693 16359 10696
rect 16301 10687 16359 10693
rect 16574 10684 16580 10696
rect 16632 10684 16638 10736
rect 1578 10616 1584 10668
rect 1636 10656 1642 10668
rect 1673 10659 1731 10665
rect 1673 10656 1685 10659
rect 1636 10628 1685 10656
rect 1636 10616 1642 10628
rect 1673 10625 1685 10628
rect 1719 10625 1731 10659
rect 1673 10619 1731 10625
rect 8846 10616 8852 10668
rect 8904 10656 8910 10668
rect 9677 10659 9735 10665
rect 9677 10656 9689 10659
rect 8904 10628 9689 10656
rect 8904 10616 8910 10628
rect 9677 10625 9689 10628
rect 9723 10625 9735 10659
rect 9677 10619 9735 10625
rect 10505 10659 10563 10665
rect 10505 10625 10517 10659
rect 10551 10625 10563 10659
rect 10505 10619 10563 10625
rect 11149 10659 11207 10665
rect 11149 10625 11161 10659
rect 11195 10656 11207 10659
rect 11238 10656 11244 10668
rect 11195 10628 11244 10656
rect 11195 10625 11207 10628
rect 11149 10619 11207 10625
rect 10520 10588 10548 10619
rect 11238 10616 11244 10628
rect 11296 10616 11302 10668
rect 11330 10616 11336 10668
rect 11388 10656 11394 10668
rect 11977 10659 12035 10665
rect 11977 10656 11989 10659
rect 11388 10628 11989 10656
rect 11388 10616 11394 10628
rect 11977 10625 11989 10628
rect 12023 10625 12035 10659
rect 11977 10619 12035 10625
rect 10520 10560 11100 10588
rect 1857 10523 1915 10529
rect 1857 10489 1869 10523
rect 1903 10520 1915 10523
rect 8846 10520 8852 10532
rect 1903 10492 8852 10520
rect 1903 10489 1915 10492
rect 1857 10483 1915 10489
rect 8846 10480 8852 10492
rect 8904 10480 8910 10532
rect 9769 10523 9827 10529
rect 9769 10489 9781 10523
rect 9815 10520 9827 10523
rect 10962 10520 10968 10532
rect 9815 10492 10968 10520
rect 9815 10489 9827 10492
rect 9769 10483 9827 10489
rect 10962 10480 10968 10492
rect 11020 10480 11026 10532
rect 11072 10520 11100 10560
rect 12250 10548 12256 10600
rect 12308 10588 12314 10600
rect 12526 10588 12532 10600
rect 12308 10560 12532 10588
rect 12308 10548 12314 10560
rect 12526 10548 12532 10560
rect 12584 10548 12590 10600
rect 12621 10591 12679 10597
rect 12621 10557 12633 10591
rect 12667 10588 12679 10591
rect 13262 10588 13268 10600
rect 12667 10560 13125 10588
rect 13223 10560 13268 10588
rect 12667 10557 12679 10560
rect 12621 10551 12679 10557
rect 11606 10520 11612 10532
rect 11072 10492 11612 10520
rect 11606 10480 11612 10492
rect 11664 10480 11670 10532
rect 13097 10520 13125 10560
rect 13262 10548 13268 10560
rect 13320 10548 13326 10600
rect 13998 10548 14004 10600
rect 14056 10588 14062 10600
rect 14461 10591 14519 10597
rect 14461 10588 14473 10591
rect 14056 10560 14473 10588
rect 14056 10548 14062 10560
rect 14461 10557 14473 10560
rect 14507 10557 14519 10591
rect 14461 10551 14519 10557
rect 14918 10548 14924 10600
rect 14976 10588 14982 10600
rect 15657 10591 15715 10597
rect 15657 10588 15669 10591
rect 14976 10560 15669 10588
rect 14976 10548 14982 10560
rect 15657 10557 15669 10560
rect 15703 10557 15715 10591
rect 16960 10588 16988 10764
rect 17236 10764 18512 10792
rect 17034 10616 17040 10668
rect 17092 10656 17098 10668
rect 17236 10665 17264 10764
rect 18506 10752 18512 10764
rect 18564 10792 18570 10804
rect 18564 10764 18828 10792
rect 18564 10752 18570 10764
rect 18800 10724 18828 10764
rect 19150 10752 19156 10804
rect 19208 10792 19214 10804
rect 21266 10792 21272 10804
rect 19208 10764 21272 10792
rect 19208 10752 19214 10764
rect 21266 10752 21272 10764
rect 21324 10752 21330 10804
rect 21361 10795 21419 10801
rect 21361 10761 21373 10795
rect 21407 10792 21419 10795
rect 21634 10792 21640 10804
rect 21407 10764 21640 10792
rect 21407 10761 21419 10764
rect 21361 10755 21419 10761
rect 21634 10752 21640 10764
rect 21692 10752 21698 10804
rect 22066 10764 24348 10792
rect 20162 10724 20168 10736
rect 18800 10696 20168 10724
rect 17221 10659 17279 10665
rect 17221 10656 17233 10659
rect 17092 10628 17233 10656
rect 17092 10616 17098 10628
rect 17221 10625 17233 10628
rect 17267 10625 17279 10659
rect 19518 10656 19524 10668
rect 18630 10628 19524 10656
rect 17221 10619 17279 10625
rect 19518 10616 19524 10628
rect 19576 10616 19582 10668
rect 19628 10665 19656 10696
rect 20162 10684 20168 10696
rect 20220 10684 20226 10736
rect 22066 10724 22094 10764
rect 24320 10733 24348 10764
rect 21376 10696 22094 10724
rect 24305 10727 24363 10733
rect 19613 10659 19671 10665
rect 19613 10625 19625 10659
rect 19659 10625 19671 10659
rect 19613 10619 19671 10625
rect 20990 10616 20996 10668
rect 21048 10616 21054 10668
rect 17497 10591 17555 10597
rect 17497 10588 17509 10591
rect 16960 10560 17509 10588
rect 15657 10551 15715 10557
rect 17497 10557 17509 10560
rect 17543 10588 17555 10591
rect 18874 10588 18880 10600
rect 17543 10560 18880 10588
rect 17543 10557 17555 10560
rect 17497 10551 17555 10557
rect 18874 10548 18880 10560
rect 18932 10548 18938 10600
rect 18969 10591 19027 10597
rect 18969 10557 18981 10591
rect 19015 10588 19027 10591
rect 19058 10588 19064 10600
rect 19015 10560 19064 10588
rect 19015 10557 19027 10560
rect 18969 10551 19027 10557
rect 19058 10548 19064 10560
rect 19116 10548 19122 10600
rect 19889 10591 19947 10597
rect 19889 10557 19901 10591
rect 19935 10588 19947 10591
rect 21266 10588 21272 10600
rect 19935 10560 21272 10588
rect 19935 10557 19947 10560
rect 19889 10551 19947 10557
rect 21266 10548 21272 10560
rect 21324 10548 21330 10600
rect 14826 10520 14832 10532
rect 13097 10492 14832 10520
rect 14826 10480 14832 10492
rect 14884 10480 14890 10532
rect 15010 10520 15016 10532
rect 14923 10492 15016 10520
rect 15010 10480 15016 10492
rect 15068 10480 15074 10532
rect 8110 10452 8116 10464
rect 8071 10424 8116 10452
rect 8110 10412 8116 10424
rect 8168 10412 8174 10464
rect 11054 10452 11060 10464
rect 11015 10424 11060 10452
rect 11054 10412 11060 10424
rect 11112 10412 11118 10464
rect 12526 10412 12532 10464
rect 12584 10452 12590 10464
rect 12802 10452 12808 10464
rect 12584 10424 12808 10452
rect 12584 10412 12590 10424
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 15028 10452 15056 10480
rect 21376 10452 21404 10696
rect 24305 10693 24317 10727
rect 24351 10693 24363 10727
rect 24854 10724 24860 10736
rect 24815 10696 24860 10724
rect 24305 10687 24363 10693
rect 24854 10684 24860 10696
rect 24912 10684 24918 10736
rect 25685 10727 25743 10733
rect 25685 10693 25697 10727
rect 25731 10724 25743 10727
rect 25774 10724 25780 10736
rect 25731 10696 25780 10724
rect 25731 10693 25743 10696
rect 25685 10687 25743 10693
rect 25774 10684 25780 10696
rect 25832 10684 25838 10736
rect 27341 10727 27399 10733
rect 27341 10693 27353 10727
rect 27387 10724 27399 10727
rect 28258 10724 28264 10736
rect 27387 10696 28264 10724
rect 27387 10693 27399 10696
rect 27341 10687 27399 10693
rect 28258 10684 28264 10696
rect 28316 10684 28322 10736
rect 28905 10659 28963 10665
rect 23414 10628 24348 10656
rect 21634 10548 21640 10600
rect 21692 10588 21698 10600
rect 22005 10591 22063 10597
rect 22005 10588 22017 10591
rect 21692 10560 22017 10588
rect 21692 10548 21698 10560
rect 22005 10557 22017 10560
rect 22051 10557 22063 10591
rect 22005 10551 22063 10557
rect 22281 10591 22339 10597
rect 22281 10557 22293 10591
rect 22327 10588 22339 10591
rect 23750 10588 23756 10600
rect 22327 10560 23756 10588
rect 22327 10557 22339 10560
rect 22281 10551 22339 10557
rect 23750 10548 23756 10560
rect 23808 10548 23814 10600
rect 24320 10520 24348 10628
rect 28905 10625 28917 10659
rect 28951 10656 28963 10659
rect 28994 10656 29000 10668
rect 28951 10628 29000 10656
rect 28951 10625 28963 10628
rect 28905 10619 28963 10625
rect 28994 10616 29000 10628
rect 29052 10616 29058 10668
rect 37553 10659 37611 10665
rect 37553 10625 37565 10659
rect 37599 10656 37611 10659
rect 38194 10656 38200 10668
rect 37599 10628 38200 10656
rect 37599 10625 37611 10628
rect 37553 10619 37611 10625
rect 38194 10616 38200 10628
rect 38252 10616 38258 10668
rect 24949 10591 25007 10597
rect 24949 10557 24961 10591
rect 24995 10588 25007 10591
rect 25130 10588 25136 10600
rect 24995 10560 25136 10588
rect 24995 10557 25007 10560
rect 24949 10551 25007 10557
rect 25130 10548 25136 10560
rect 25188 10548 25194 10600
rect 25590 10588 25596 10600
rect 25551 10560 25596 10588
rect 25590 10548 25596 10560
rect 25648 10548 25654 10600
rect 25682 10548 25688 10600
rect 25740 10588 25746 10600
rect 25869 10591 25927 10597
rect 25869 10588 25881 10591
rect 25740 10560 25881 10588
rect 25740 10548 25746 10560
rect 25869 10557 25881 10560
rect 25915 10557 25927 10591
rect 25869 10551 25927 10557
rect 27062 10548 27068 10600
rect 27120 10588 27126 10600
rect 27249 10591 27307 10597
rect 27249 10588 27261 10591
rect 27120 10560 27261 10588
rect 27120 10548 27126 10560
rect 27249 10557 27261 10560
rect 27295 10557 27307 10591
rect 27890 10588 27896 10600
rect 27851 10560 27896 10588
rect 27249 10551 27307 10557
rect 27890 10548 27896 10560
rect 27948 10548 27954 10600
rect 28721 10591 28779 10597
rect 28721 10557 28733 10591
rect 28767 10588 28779 10591
rect 28810 10588 28816 10600
rect 28767 10560 28816 10588
rect 28767 10557 28779 10560
rect 28721 10551 28779 10557
rect 28810 10548 28816 10560
rect 28868 10548 28874 10600
rect 27706 10520 27712 10532
rect 24320 10492 27712 10520
rect 27706 10480 27712 10492
rect 27764 10480 27770 10532
rect 28350 10480 28356 10532
rect 28408 10520 28414 10532
rect 29917 10523 29975 10529
rect 29917 10520 29929 10523
rect 28408 10492 29929 10520
rect 28408 10480 28414 10492
rect 29917 10489 29929 10492
rect 29963 10489 29975 10523
rect 29917 10483 29975 10489
rect 36998 10480 37004 10532
rect 37056 10520 37062 10532
rect 38013 10523 38071 10529
rect 38013 10520 38025 10523
rect 37056 10492 38025 10520
rect 37056 10480 37062 10492
rect 38013 10489 38025 10492
rect 38059 10489 38071 10523
rect 38013 10483 38071 10489
rect 15028 10424 21404 10452
rect 22830 10412 22836 10464
rect 22888 10452 22894 10464
rect 23753 10455 23811 10461
rect 23753 10452 23765 10455
rect 22888 10424 23765 10452
rect 22888 10412 22894 10424
rect 23753 10421 23765 10424
rect 23799 10421 23811 10455
rect 23753 10415 23811 10421
rect 25130 10412 25136 10464
rect 25188 10452 25194 10464
rect 28902 10452 28908 10464
rect 25188 10424 28908 10452
rect 25188 10412 25194 10424
rect 28902 10412 28908 10424
rect 28960 10412 28966 10464
rect 29362 10452 29368 10464
rect 29323 10424 29368 10452
rect 29362 10412 29368 10424
rect 29420 10412 29426 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 1578 10248 1584 10260
rect 1539 10220 1584 10248
rect 1578 10208 1584 10220
rect 1636 10208 1642 10260
rect 8573 10251 8631 10257
rect 8573 10217 8585 10251
rect 8619 10248 8631 10251
rect 8754 10248 8760 10260
rect 8619 10220 8760 10248
rect 8619 10217 8631 10220
rect 8573 10211 8631 10217
rect 8754 10208 8760 10220
rect 8812 10208 8818 10260
rect 9674 10208 9680 10260
rect 9732 10248 9738 10260
rect 10962 10248 10968 10260
rect 9732 10220 10968 10248
rect 9732 10208 9738 10220
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 11054 10208 11060 10260
rect 11112 10248 11118 10260
rect 16666 10248 16672 10260
rect 11112 10220 16672 10248
rect 11112 10208 11118 10220
rect 16666 10208 16672 10220
rect 16724 10208 16730 10260
rect 17494 10248 17500 10260
rect 16776 10220 17500 10248
rect 9030 10140 9036 10192
rect 9088 10180 9094 10192
rect 10502 10180 10508 10192
rect 9088 10152 10508 10180
rect 9088 10140 9094 10152
rect 10502 10140 10508 10152
rect 10560 10140 10566 10192
rect 10594 10140 10600 10192
rect 10652 10180 10658 10192
rect 11149 10183 11207 10189
rect 10652 10152 10732 10180
rect 10652 10140 10658 10152
rect 9858 10112 9864 10124
rect 9819 10084 9864 10112
rect 9858 10072 9864 10084
rect 9916 10072 9922 10124
rect 10605 10057 10663 10063
rect 8754 10004 8760 10056
rect 8812 10044 8818 10056
rect 9769 10047 9827 10053
rect 9769 10044 9781 10047
rect 8812 10016 9781 10044
rect 8812 10004 8818 10016
rect 9769 10013 9781 10016
rect 9815 10013 9827 10047
rect 10605 10023 10617 10057
rect 10651 10054 10663 10057
rect 10704 10054 10732 10152
rect 11149 10149 11161 10183
rect 11195 10180 11207 10183
rect 12158 10180 12164 10192
rect 11195 10152 12164 10180
rect 11195 10149 11207 10152
rect 11149 10143 11207 10149
rect 12158 10140 12164 10152
rect 12216 10140 12222 10192
rect 12986 10180 12992 10192
rect 12360 10152 12992 10180
rect 12360 10121 12388 10152
rect 12986 10140 12992 10152
rect 13044 10180 13050 10192
rect 13541 10183 13599 10189
rect 13541 10180 13553 10183
rect 13044 10152 13553 10180
rect 13044 10140 13050 10152
rect 13541 10149 13553 10152
rect 13587 10149 13599 10183
rect 13541 10143 13599 10149
rect 16301 10183 16359 10189
rect 16301 10149 16313 10183
rect 16347 10180 16359 10183
rect 16390 10180 16396 10192
rect 16347 10152 16396 10180
rect 16347 10149 16359 10152
rect 16301 10143 16359 10149
rect 16390 10140 16396 10152
rect 16448 10140 16454 10192
rect 12345 10115 12403 10121
rect 12345 10081 12357 10115
rect 12391 10081 12403 10115
rect 14918 10112 14924 10124
rect 12345 10075 12403 10081
rect 12820 10084 14924 10112
rect 10651 10026 10732 10054
rect 10651 10023 10663 10026
rect 10605 10017 10663 10023
rect 9769 10007 9827 10013
rect 10962 10004 10968 10056
rect 11020 10044 11026 10056
rect 11057 10047 11115 10053
rect 11057 10044 11069 10047
rect 11020 10016 11069 10044
rect 11020 10004 11026 10016
rect 11057 10013 11069 10016
rect 11103 10013 11115 10047
rect 11057 10007 11115 10013
rect 11330 10004 11336 10056
rect 11388 10044 11394 10056
rect 11701 10047 11759 10053
rect 11701 10044 11713 10047
rect 11388 10016 11713 10044
rect 11388 10004 11394 10016
rect 11701 10013 11713 10016
rect 11747 10013 11759 10047
rect 11701 10007 11759 10013
rect 12820 9988 12848 10084
rect 14918 10072 14924 10084
rect 14976 10072 14982 10124
rect 15194 10072 15200 10124
rect 15252 10112 15258 10124
rect 16776 10112 16804 10220
rect 17494 10208 17500 10220
rect 17552 10248 17558 10260
rect 19150 10248 19156 10260
rect 17552 10220 19156 10248
rect 17552 10208 17558 10220
rect 19150 10208 19156 10220
rect 19208 10208 19214 10260
rect 21358 10208 21364 10260
rect 21416 10248 21422 10260
rect 21416 10220 22968 10248
rect 21416 10208 21422 10220
rect 18414 10140 18420 10192
rect 18472 10180 18478 10192
rect 19242 10180 19248 10192
rect 18472 10152 19248 10180
rect 18472 10140 18478 10152
rect 19242 10140 19248 10152
rect 19300 10140 19306 10192
rect 19610 10140 19616 10192
rect 19668 10180 19674 10192
rect 22940 10180 22968 10220
rect 23290 10208 23296 10260
rect 23348 10248 23354 10260
rect 23937 10251 23995 10257
rect 23937 10248 23949 10251
rect 23348 10220 23949 10248
rect 23348 10208 23354 10220
rect 23937 10217 23949 10220
rect 23983 10217 23995 10251
rect 23937 10211 23995 10217
rect 25038 10208 25044 10260
rect 25096 10248 25102 10260
rect 25958 10248 25964 10260
rect 25096 10220 25964 10248
rect 25096 10208 25102 10220
rect 25958 10208 25964 10220
rect 26016 10248 26022 10260
rect 29086 10248 29092 10260
rect 26016 10220 29092 10248
rect 26016 10208 26022 10220
rect 29086 10208 29092 10220
rect 29144 10208 29150 10260
rect 25130 10180 25136 10192
rect 19668 10152 21772 10180
rect 22940 10152 25136 10180
rect 19668 10140 19674 10152
rect 17034 10112 17040 10124
rect 15252 10084 16804 10112
rect 16995 10084 17040 10112
rect 15252 10072 15258 10084
rect 17034 10072 17040 10084
rect 17092 10072 17098 10124
rect 17310 10112 17316 10124
rect 17271 10084 17316 10112
rect 17310 10072 17316 10084
rect 17368 10112 17374 10124
rect 17862 10112 17868 10124
rect 17368 10084 17868 10112
rect 17368 10072 17374 10084
rect 17862 10072 17868 10084
rect 17920 10112 17926 10124
rect 20732 10121 20760 10152
rect 20717 10115 20775 10121
rect 17920 10084 19380 10112
rect 17920 10072 17926 10084
rect 14458 10004 14464 10056
rect 14516 10044 14522 10056
rect 14553 10047 14611 10053
rect 14553 10044 14565 10047
rect 14516 10016 14565 10044
rect 14516 10004 14522 10016
rect 14553 10013 14565 10016
rect 14599 10013 14611 10047
rect 19352 10046 19380 10084
rect 20717 10081 20729 10115
rect 20763 10081 20775 10115
rect 20717 10075 20775 10081
rect 20898 10072 20904 10124
rect 20956 10112 20962 10124
rect 20993 10115 21051 10121
rect 20993 10112 21005 10115
rect 20956 10084 21005 10112
rect 20956 10072 20962 10084
rect 20993 10081 21005 10084
rect 21039 10081 21051 10115
rect 21634 10112 21640 10124
rect 21595 10084 21640 10112
rect 20993 10075 21051 10081
rect 21634 10072 21640 10084
rect 21692 10072 21698 10124
rect 21744 10112 21772 10152
rect 25130 10140 25136 10152
rect 25188 10140 25194 10192
rect 25314 10140 25320 10192
rect 25372 10180 25378 10192
rect 26513 10183 26571 10189
rect 26513 10180 26525 10183
rect 25372 10152 26525 10180
rect 25372 10140 25378 10152
rect 26513 10149 26525 10152
rect 26559 10149 26571 10183
rect 26513 10143 26571 10149
rect 26602 10140 26608 10192
rect 26660 10180 26666 10192
rect 28258 10180 28264 10192
rect 26660 10152 28264 10180
rect 26660 10140 26666 10152
rect 28258 10140 28264 10152
rect 28316 10140 28322 10192
rect 22278 10112 22284 10124
rect 21744 10084 22284 10112
rect 22278 10072 22284 10084
rect 22336 10072 22342 10124
rect 29362 10112 29368 10124
rect 27816 10084 29368 10112
rect 19429 10047 19487 10053
rect 19429 10046 19441 10047
rect 19352 10018 19441 10046
rect 14553 10007 14611 10013
rect 19429 10013 19441 10018
rect 19475 10013 19487 10047
rect 19429 10007 19487 10013
rect 19536 10044 19656 10046
rect 20346 10044 20352 10056
rect 19536 10018 20352 10044
rect 10505 9979 10563 9985
rect 10505 9945 10517 9979
rect 10551 9976 10563 9979
rect 12250 9976 12256 9988
rect 10551 9948 11836 9976
rect 12211 9948 12256 9976
rect 10551 9945 10563 9948
rect 10505 9939 10563 9945
rect 9309 9911 9367 9917
rect 9309 9877 9321 9911
rect 9355 9908 9367 9911
rect 9398 9908 9404 9920
rect 9355 9880 9404 9908
rect 9355 9877 9367 9880
rect 9309 9871 9367 9877
rect 9398 9868 9404 9880
rect 9456 9908 9462 9920
rect 11238 9908 11244 9920
rect 9456 9880 11244 9908
rect 9456 9868 9462 9880
rect 11238 9868 11244 9880
rect 11296 9868 11302 9920
rect 11808 9908 11836 9948
rect 12250 9936 12256 9948
rect 12308 9936 12314 9988
rect 12802 9936 12808 9988
rect 12860 9976 12866 9988
rect 12989 9979 13047 9985
rect 12989 9976 13001 9979
rect 12860 9948 13001 9976
rect 12860 9936 12866 9948
rect 12989 9945 13001 9948
rect 13035 9945 13047 9979
rect 12989 9939 13047 9945
rect 13081 9979 13139 9985
rect 13081 9945 13093 9979
rect 13127 9976 13139 9979
rect 13354 9976 13360 9988
rect 13127 9948 13360 9976
rect 13127 9945 13139 9948
rect 13081 9939 13139 9945
rect 13354 9936 13360 9948
rect 13412 9936 13418 9988
rect 14829 9979 14887 9985
rect 14829 9945 14841 9979
rect 14875 9976 14887 9979
rect 14918 9976 14924 9988
rect 14875 9948 14924 9976
rect 14875 9945 14887 9948
rect 14829 9939 14887 9945
rect 14918 9936 14924 9948
rect 14976 9936 14982 9988
rect 16482 9976 16488 9988
rect 16054 9948 16488 9976
rect 16482 9936 16488 9948
rect 16540 9936 16546 9988
rect 16758 9936 16764 9988
rect 16816 9976 16822 9988
rect 17310 9976 17316 9988
rect 16816 9948 17316 9976
rect 16816 9936 16822 9948
rect 17310 9936 17316 9948
rect 17368 9936 17374 9988
rect 18322 9936 18328 9988
rect 18380 9936 18386 9988
rect 19536 9976 19564 10018
rect 19628 10016 20352 10018
rect 20346 10004 20352 10016
rect 20404 10004 20410 10056
rect 24762 10044 24768 10056
rect 23046 10016 24768 10044
rect 24762 10004 24768 10016
rect 24820 10004 24826 10056
rect 27522 10004 27528 10056
rect 27580 10044 27586 10056
rect 27816 10053 27844 10084
rect 29362 10072 29368 10084
rect 29420 10072 29426 10124
rect 27801 10047 27859 10053
rect 27801 10044 27813 10047
rect 27580 10016 27813 10044
rect 27580 10004 27586 10016
rect 27801 10013 27813 10016
rect 27847 10013 27859 10047
rect 28994 10044 29000 10056
rect 28907 10016 29000 10044
rect 27801 10007 27859 10013
rect 28994 10004 29000 10016
rect 29052 10044 29058 10056
rect 30190 10044 30196 10056
rect 29052 10016 30196 10044
rect 29052 10004 29058 10016
rect 30190 10004 30196 10016
rect 30248 10004 30254 10056
rect 19168 9948 19564 9976
rect 19168 9920 19196 9948
rect 19610 9936 19616 9988
rect 19668 9976 19674 9988
rect 20898 9976 20904 9988
rect 19668 9948 20668 9976
rect 20859 9948 20904 9976
rect 19668 9936 19674 9948
rect 20640 9920 20668 9948
rect 20898 9936 20904 9948
rect 20956 9936 20962 9988
rect 21450 9936 21456 9988
rect 21508 9976 21514 9988
rect 21910 9976 21916 9988
rect 21508 9948 21916 9976
rect 21508 9936 21514 9948
rect 21910 9936 21916 9948
rect 21968 9936 21974 9988
rect 24670 9936 24676 9988
rect 24728 9976 24734 9988
rect 24949 9979 25007 9985
rect 24949 9976 24961 9979
rect 24728 9948 24961 9976
rect 24728 9936 24734 9948
rect 24949 9945 24961 9948
rect 24995 9945 25007 9979
rect 24949 9939 25007 9945
rect 25038 9936 25044 9988
rect 25096 9976 25102 9988
rect 25958 9976 25964 9988
rect 25096 9948 25141 9976
rect 25919 9948 25964 9976
rect 25096 9936 25102 9948
rect 25958 9936 25964 9948
rect 26016 9936 26022 9988
rect 26142 9936 26148 9988
rect 26200 9976 26206 9988
rect 26973 9979 27031 9985
rect 26973 9976 26985 9979
rect 26200 9948 26985 9976
rect 26200 9936 26206 9948
rect 26973 9945 26985 9948
rect 27019 9945 27031 9979
rect 26973 9939 27031 9945
rect 27062 9936 27068 9988
rect 27120 9976 27126 9988
rect 27120 9948 27165 9976
rect 27120 9936 27126 9948
rect 28626 9936 28632 9988
rect 28684 9976 28690 9988
rect 28721 9979 28779 9985
rect 28721 9976 28733 9979
rect 28684 9948 28733 9976
rect 28684 9936 28690 9948
rect 28721 9945 28733 9948
rect 28767 9945 28779 9979
rect 29914 9976 29920 9988
rect 29875 9948 29920 9976
rect 28721 9939 28779 9945
rect 29914 9936 29920 9948
rect 29972 9936 29978 9988
rect 13170 9908 13176 9920
rect 11808 9880 13176 9908
rect 13170 9868 13176 9880
rect 13228 9868 13234 9920
rect 18782 9868 18788 9920
rect 18840 9908 18846 9920
rect 19150 9908 19156 9920
rect 18840 9880 19156 9908
rect 18840 9868 18846 9880
rect 19150 9868 19156 9880
rect 19208 9868 19214 9920
rect 19521 9911 19579 9917
rect 19521 9877 19533 9911
rect 19567 9908 19579 9911
rect 19702 9908 19708 9920
rect 19567 9880 19708 9908
rect 19567 9877 19579 9880
rect 19521 9871 19579 9877
rect 19702 9868 19708 9880
rect 19760 9868 19766 9920
rect 20622 9868 20628 9920
rect 20680 9908 20686 9920
rect 23290 9908 23296 9920
rect 20680 9880 23296 9908
rect 20680 9868 20686 9880
rect 23290 9868 23296 9880
rect 23348 9868 23354 9920
rect 23382 9868 23388 9920
rect 23440 9908 23446 9920
rect 23440 9880 23485 9908
rect 23440 9868 23446 9880
rect 26234 9868 26240 9920
rect 26292 9908 26298 9920
rect 27709 9911 27767 9917
rect 27709 9908 27721 9911
rect 26292 9880 27721 9908
rect 26292 9868 26298 9880
rect 27709 9877 27721 9880
rect 27755 9877 27767 9911
rect 27709 9871 27767 9877
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 9122 9664 9128 9716
rect 9180 9704 9186 9716
rect 12802 9704 12808 9716
rect 9180 9676 12808 9704
rect 9180 9664 9186 9676
rect 12802 9664 12808 9676
rect 12860 9664 12866 9716
rect 13998 9704 14004 9716
rect 12912 9676 13400 9704
rect 13959 9676 14004 9704
rect 9674 9596 9680 9648
rect 9732 9636 9738 9648
rect 9769 9639 9827 9645
rect 9769 9636 9781 9639
rect 9732 9608 9781 9636
rect 9732 9596 9738 9608
rect 9769 9605 9781 9608
rect 9815 9605 9827 9639
rect 9769 9599 9827 9605
rect 10318 9596 10324 9648
rect 10376 9636 10382 9648
rect 10413 9639 10471 9645
rect 10413 9636 10425 9639
rect 10376 9608 10425 9636
rect 10376 9596 10382 9608
rect 10413 9605 10425 9608
rect 10459 9605 10471 9639
rect 11238 9636 11244 9648
rect 10413 9599 10471 9605
rect 10520 9608 11244 9636
rect 10520 9577 10548 9608
rect 11238 9596 11244 9608
rect 11296 9596 11302 9648
rect 12912 9636 12940 9676
rect 11992 9608 12940 9636
rect 12989 9639 13047 9645
rect 11992 9577 12020 9608
rect 12989 9605 13001 9639
rect 13035 9636 13047 9639
rect 13372 9636 13400 9676
rect 13998 9664 14004 9676
rect 14056 9664 14062 9716
rect 14826 9664 14832 9716
rect 14884 9704 14890 9716
rect 17954 9704 17960 9716
rect 14884 9676 17960 9704
rect 14884 9664 14890 9676
rect 14734 9636 14740 9648
rect 13035 9608 13308 9636
rect 13372 9608 14740 9636
rect 13035 9605 13047 9608
rect 12989 9599 13047 9605
rect 13280 9580 13308 9608
rect 14734 9596 14740 9608
rect 14792 9596 14798 9648
rect 10505 9571 10563 9577
rect 10505 9537 10517 9571
rect 10551 9537 10563 9571
rect 10505 9531 10563 9537
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9537 11207 9571
rect 11149 9531 11207 9537
rect 11977 9571 12035 9577
rect 11977 9537 11989 9571
rect 12023 9537 12035 9571
rect 11977 9531 12035 9537
rect 9309 9503 9367 9509
rect 9309 9469 9321 9503
rect 9355 9500 9367 9503
rect 11164 9500 11192 9531
rect 13262 9528 13268 9580
rect 13320 9528 13326 9580
rect 16224 9568 16252 9676
rect 17954 9664 17960 9676
rect 18012 9664 18018 9716
rect 19058 9664 19064 9716
rect 19116 9704 19122 9716
rect 19116 9676 20944 9704
rect 19116 9664 19122 9676
rect 16482 9596 16488 9648
rect 16540 9636 16546 9648
rect 17497 9639 17555 9645
rect 17497 9636 17509 9639
rect 16540 9608 17509 9636
rect 16540 9596 16546 9608
rect 17497 9605 17509 9608
rect 17543 9605 17555 9639
rect 17497 9599 17555 9605
rect 17589 9639 17647 9645
rect 17589 9605 17601 9639
rect 17635 9636 17647 9639
rect 18138 9636 18144 9648
rect 17635 9608 18144 9636
rect 17635 9605 17647 9608
rect 17589 9599 17647 9605
rect 18138 9596 18144 9608
rect 18196 9596 18202 9648
rect 20916 9636 20944 9676
rect 20990 9664 20996 9716
rect 21048 9704 21054 9716
rect 21048 9676 24716 9704
rect 21048 9664 21054 9676
rect 21361 9639 21419 9645
rect 19458 9608 20852 9636
rect 20916 9608 21312 9636
rect 16945 9571 17003 9577
rect 16945 9568 16957 9571
rect 12342 9500 12348 9512
rect 9355 9472 12348 9500
rect 9355 9469 9367 9472
rect 9309 9463 9367 9469
rect 12342 9460 12348 9472
rect 12400 9460 12406 9512
rect 12618 9460 12624 9512
rect 12676 9500 12682 9512
rect 13081 9503 13139 9509
rect 13081 9500 13093 9503
rect 12676 9472 13093 9500
rect 12676 9460 12682 9472
rect 13081 9469 13093 9472
rect 13127 9469 13139 9503
rect 14458 9500 14464 9512
rect 14419 9472 14464 9500
rect 13081 9463 13139 9469
rect 14458 9460 14464 9472
rect 14516 9460 14522 9512
rect 7190 9392 7196 9444
rect 7248 9432 7254 9444
rect 10965 9435 11023 9441
rect 10965 9432 10977 9435
rect 7248 9404 10977 9432
rect 7248 9392 7254 9404
rect 10965 9401 10977 9404
rect 11011 9401 11023 9435
rect 10965 9395 11023 9401
rect 12529 9435 12587 9441
rect 12529 9401 12541 9435
rect 12575 9432 12587 9435
rect 12894 9432 12900 9444
rect 12575 9404 12900 9432
rect 12575 9401 12587 9404
rect 12529 9395 12587 9401
rect 12894 9392 12900 9404
rect 12952 9392 12958 9444
rect 8754 9364 8760 9376
rect 8715 9336 8760 9364
rect 8754 9324 8760 9336
rect 8812 9324 8818 9376
rect 10410 9324 10416 9376
rect 10468 9364 10474 9376
rect 10778 9364 10784 9376
rect 10468 9336 10784 9364
rect 10468 9324 10474 9336
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 11885 9367 11943 9373
rect 11885 9333 11897 9367
rect 11931 9364 11943 9367
rect 13906 9364 13912 9376
rect 11931 9336 13912 9364
rect 11931 9333 11943 9336
rect 11885 9327 11943 9333
rect 13906 9324 13912 9336
rect 13964 9324 13970 9376
rect 13998 9324 14004 9376
rect 14056 9364 14062 9376
rect 14724 9367 14782 9373
rect 14724 9364 14736 9367
rect 14056 9336 14736 9364
rect 14056 9324 14062 9336
rect 14724 9333 14736 9336
rect 14770 9364 14782 9367
rect 15746 9364 15752 9376
rect 14770 9336 15752 9364
rect 14770 9333 14782 9336
rect 14724 9327 14782 9333
rect 15746 9324 15752 9336
rect 15804 9324 15810 9376
rect 15856 9364 15884 9554
rect 16224 9540 16957 9568
rect 16945 9537 16957 9540
rect 16991 9537 17003 9571
rect 16945 9531 17003 9537
rect 20162 9528 20168 9580
rect 20220 9568 20226 9580
rect 20220 9540 20265 9568
rect 20220 9528 20226 9540
rect 20346 9528 20352 9580
rect 20404 9568 20410 9580
rect 20625 9571 20683 9577
rect 20625 9568 20637 9571
rect 20404 9540 20637 9568
rect 20404 9528 20410 9540
rect 20625 9537 20637 9540
rect 20671 9537 20683 9571
rect 20625 9531 20683 9537
rect 16209 9503 16267 9509
rect 16209 9469 16221 9503
rect 16255 9500 16267 9503
rect 16758 9500 16764 9512
rect 16255 9472 16764 9500
rect 16255 9469 16267 9472
rect 16209 9463 16267 9469
rect 16758 9460 16764 9472
rect 16816 9460 16822 9512
rect 16850 9460 16856 9512
rect 16908 9500 16914 9512
rect 17770 9500 17776 9512
rect 16908 9472 17776 9500
rect 16908 9460 16914 9472
rect 17770 9460 17776 9472
rect 17828 9500 17834 9512
rect 18141 9503 18199 9509
rect 18141 9500 18153 9503
rect 17828 9472 18153 9500
rect 17828 9460 17834 9472
rect 18141 9469 18153 9472
rect 18187 9469 18199 9503
rect 19334 9500 19340 9512
rect 18141 9463 18199 9469
rect 18248 9472 19340 9500
rect 16390 9392 16396 9444
rect 16448 9432 16454 9444
rect 18248 9432 18276 9472
rect 19334 9460 19340 9472
rect 19392 9460 19398 9512
rect 19889 9503 19947 9509
rect 19889 9469 19901 9503
rect 19935 9500 19947 9503
rect 20824 9500 20852 9608
rect 21284 9577 21312 9608
rect 21361 9605 21373 9639
rect 21407 9636 21419 9639
rect 22186 9636 22192 9648
rect 21407 9608 22192 9636
rect 21407 9605 21419 9608
rect 21361 9599 21419 9605
rect 22186 9596 22192 9608
rect 22244 9596 22250 9648
rect 24210 9636 24216 9648
rect 23506 9608 24216 9636
rect 24210 9596 24216 9608
rect 24268 9596 24274 9648
rect 24394 9636 24400 9648
rect 24355 9608 24400 9636
rect 24394 9596 24400 9608
rect 24452 9596 24458 9648
rect 21269 9571 21327 9577
rect 21269 9537 21281 9571
rect 21315 9537 21327 9571
rect 21269 9531 21327 9537
rect 21634 9528 21640 9580
rect 21692 9568 21698 9580
rect 22005 9571 22063 9577
rect 22005 9568 22017 9571
rect 21692 9540 22017 9568
rect 21692 9528 21698 9540
rect 22005 9537 22017 9540
rect 22051 9537 22063 9571
rect 22005 9531 22063 9537
rect 24118 9528 24124 9580
rect 24176 9568 24182 9580
rect 24305 9571 24363 9577
rect 24305 9568 24317 9571
rect 24176 9540 24317 9568
rect 24176 9528 24182 9540
rect 24305 9537 24317 9540
rect 24351 9537 24363 9571
rect 24688 9568 24716 9676
rect 24762 9664 24768 9716
rect 24820 9704 24826 9716
rect 27430 9704 27436 9716
rect 24820 9676 27436 9704
rect 24820 9664 24826 9676
rect 27430 9664 27436 9676
rect 27488 9664 27494 9716
rect 28350 9704 28356 9716
rect 28000 9676 28356 9704
rect 24946 9636 24952 9648
rect 24907 9608 24952 9636
rect 24946 9596 24952 9608
rect 25004 9596 25010 9648
rect 25501 9639 25559 9645
rect 25501 9605 25513 9639
rect 25547 9636 25559 9639
rect 26234 9636 26240 9648
rect 25547 9608 26240 9636
rect 25547 9605 25559 9608
rect 25501 9599 25559 9605
rect 26234 9596 26240 9608
rect 26292 9596 26298 9648
rect 26418 9596 26424 9648
rect 26476 9636 26482 9648
rect 27249 9639 27307 9645
rect 27249 9636 27261 9639
rect 26476 9608 27261 9636
rect 26476 9596 26482 9608
rect 27249 9605 27261 9608
rect 27295 9605 27307 9639
rect 27522 9636 27528 9648
rect 27249 9599 27307 9605
rect 27356 9608 27528 9636
rect 26326 9568 26332 9580
rect 24688 9540 24992 9568
rect 26287 9540 26332 9568
rect 24305 9531 24363 9537
rect 24964 9512 24992 9540
rect 26326 9528 26332 9540
rect 26384 9528 26390 9580
rect 27356 9577 27384 9608
rect 27522 9596 27528 9608
rect 27580 9596 27586 9648
rect 27614 9596 27620 9648
rect 27672 9636 27678 9648
rect 27893 9639 27951 9645
rect 27893 9636 27905 9639
rect 27672 9608 27905 9636
rect 27672 9596 27678 9608
rect 27893 9605 27905 9608
rect 27939 9605 27951 9639
rect 28000 9636 28028 9676
rect 28350 9664 28356 9676
rect 28408 9664 28414 9716
rect 28534 9664 28540 9716
rect 28592 9704 28598 9716
rect 28592 9676 29040 9704
rect 28592 9664 28598 9676
rect 28000 9608 28120 9636
rect 27893 9599 27951 9605
rect 27341 9571 27399 9577
rect 27341 9537 27353 9571
rect 27387 9537 27399 9571
rect 27341 9531 27399 9537
rect 27985 9571 28043 9577
rect 27985 9537 27997 9571
rect 28031 9568 28043 9571
rect 28092 9568 28120 9608
rect 28166 9596 28172 9648
rect 28224 9636 28230 9648
rect 28905 9639 28963 9645
rect 28905 9636 28917 9639
rect 28224 9608 28917 9636
rect 28224 9596 28230 9608
rect 28905 9605 28917 9608
rect 28951 9605 28963 9639
rect 29012 9636 29040 9676
rect 30837 9639 30895 9645
rect 30837 9636 30849 9639
rect 29012 9608 30849 9636
rect 28905 9599 28963 9605
rect 30837 9605 30849 9608
rect 30883 9636 30895 9639
rect 36998 9636 37004 9648
rect 30883 9608 37004 9636
rect 30883 9605 30895 9608
rect 30837 9599 30895 9605
rect 36998 9596 37004 9608
rect 37056 9596 37062 9648
rect 28031 9540 28120 9568
rect 28031 9537 28043 9540
rect 27985 9531 28043 9537
rect 29914 9528 29920 9580
rect 29972 9568 29978 9580
rect 34241 9571 34299 9577
rect 34241 9568 34253 9571
rect 29972 9540 34253 9568
rect 29972 9528 29978 9540
rect 34241 9537 34253 9540
rect 34287 9537 34299 9571
rect 34241 9531 34299 9537
rect 22281 9503 22339 9509
rect 19935 9472 20760 9500
rect 20824 9472 22054 9500
rect 19935 9469 19947 9472
rect 19889 9463 19947 9469
rect 16448 9404 18276 9432
rect 20732 9432 20760 9472
rect 22048 9448 22054 9472
rect 22106 9448 22112 9500
rect 22281 9469 22293 9503
rect 22327 9500 22339 9503
rect 22370 9500 22376 9512
rect 22327 9472 22376 9500
rect 22327 9469 22339 9472
rect 22281 9463 22339 9469
rect 22370 9460 22376 9472
rect 22428 9460 22434 9512
rect 22646 9460 22652 9512
rect 22704 9500 22710 9512
rect 24854 9500 24860 9512
rect 22704 9472 24860 9500
rect 22704 9460 22710 9472
rect 24854 9460 24860 9472
rect 24912 9460 24918 9512
rect 24946 9460 24952 9512
rect 25004 9460 25010 9512
rect 25593 9503 25651 9509
rect 25593 9469 25605 9503
rect 25639 9500 25651 9503
rect 26237 9503 26295 9509
rect 26237 9500 26249 9503
rect 25639 9472 26249 9500
rect 25639 9469 25651 9472
rect 25593 9463 25651 9469
rect 26237 9469 26249 9472
rect 26283 9500 26295 9503
rect 27062 9500 27068 9512
rect 26283 9472 27068 9500
rect 26283 9469 26295 9472
rect 26237 9463 26295 9469
rect 27062 9460 27068 9472
rect 27120 9460 27126 9512
rect 27154 9460 27160 9512
rect 27212 9500 27218 9512
rect 27798 9500 27804 9512
rect 27212 9472 27804 9500
rect 27212 9460 27218 9472
rect 27798 9460 27804 9472
rect 27856 9460 27862 9512
rect 27890 9460 27896 9512
rect 27948 9500 27954 9512
rect 28813 9503 28871 9509
rect 28813 9500 28825 9503
rect 27948 9472 28825 9500
rect 27948 9460 27954 9472
rect 28813 9469 28825 9472
rect 28859 9469 28871 9503
rect 29086 9500 29092 9512
rect 29047 9472 29092 9500
rect 28813 9463 28871 9469
rect 29086 9460 29092 9472
rect 29144 9460 29150 9512
rect 29362 9460 29368 9512
rect 29420 9500 29426 9512
rect 31389 9503 31447 9509
rect 31389 9500 31401 9503
rect 29420 9472 31401 9500
rect 29420 9460 29426 9472
rect 31389 9469 31401 9472
rect 31435 9469 31447 9503
rect 31389 9463 31447 9469
rect 21174 9432 21180 9444
rect 20732 9404 21180 9432
rect 16448 9392 16454 9404
rect 21174 9392 21180 9404
rect 21232 9432 21238 9444
rect 21542 9432 21548 9444
rect 21232 9404 21548 9432
rect 21232 9392 21238 9404
rect 21542 9392 21548 9404
rect 21600 9392 21606 9444
rect 23290 9392 23296 9444
rect 23348 9432 23354 9444
rect 27522 9432 27528 9444
rect 23348 9404 27528 9432
rect 23348 9392 23354 9404
rect 27522 9392 27528 9404
rect 27580 9392 27586 9444
rect 27614 9392 27620 9444
rect 27672 9432 27678 9444
rect 28994 9432 29000 9444
rect 27672 9404 29000 9432
rect 27672 9392 27678 9404
rect 28994 9392 29000 9404
rect 29052 9392 29058 9444
rect 20070 9364 20076 9376
rect 15856 9336 20076 9364
rect 20070 9324 20076 9336
rect 20128 9324 20134 9376
rect 20714 9364 20720 9376
rect 20675 9336 20720 9364
rect 20714 9324 20720 9336
rect 20772 9324 20778 9376
rect 20806 9324 20812 9376
rect 20864 9364 20870 9376
rect 21266 9364 21272 9376
rect 20864 9336 21272 9364
rect 20864 9324 20870 9336
rect 21266 9324 21272 9336
rect 21324 9324 21330 9376
rect 22002 9324 22008 9376
rect 22060 9364 22066 9376
rect 22738 9364 22744 9376
rect 22060 9336 22744 9364
rect 22060 9324 22066 9336
rect 22738 9324 22744 9336
rect 22796 9364 22802 9376
rect 23382 9364 23388 9376
rect 22796 9336 23388 9364
rect 22796 9324 22802 9336
rect 23382 9324 23388 9336
rect 23440 9324 23446 9376
rect 23750 9364 23756 9376
rect 23711 9336 23756 9364
rect 23750 9324 23756 9336
rect 23808 9324 23814 9376
rect 24118 9324 24124 9376
rect 24176 9364 24182 9376
rect 30285 9367 30343 9373
rect 30285 9364 30297 9367
rect 24176 9336 30297 9364
rect 24176 9324 24182 9336
rect 30285 9333 30297 9336
rect 30331 9333 30343 9367
rect 30285 9327 30343 9333
rect 33686 9324 33692 9376
rect 33744 9364 33750 9376
rect 34333 9367 34391 9373
rect 34333 9364 34345 9367
rect 33744 9336 34345 9364
rect 33744 9324 33750 9336
rect 34333 9333 34345 9336
rect 34379 9333 34391 9367
rect 34333 9327 34391 9333
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 9766 9120 9772 9172
rect 9824 9160 9830 9172
rect 11330 9160 11336 9172
rect 9824 9132 11336 9160
rect 9824 9120 9830 9132
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 11514 9160 11520 9172
rect 11475 9132 11520 9160
rect 11514 9120 11520 9132
rect 11572 9120 11578 9172
rect 11790 9120 11796 9172
rect 11848 9160 11854 9172
rect 11848 9132 15700 9160
rect 11848 9120 11854 9132
rect 13814 9052 13820 9104
rect 13872 9092 13878 9104
rect 14366 9092 14372 9104
rect 13872 9064 14372 9092
rect 13872 9052 13878 9064
rect 14366 9052 14372 9064
rect 14424 9052 14430 9104
rect 15672 9092 15700 9132
rect 16684 9132 24532 9160
rect 16482 9092 16488 9104
rect 15672 9064 16488 9092
rect 16482 9052 16488 9064
rect 16540 9052 16546 9104
rect 1857 9027 1915 9033
rect 1857 8993 1869 9027
rect 1903 9024 1915 9027
rect 7282 9024 7288 9036
rect 1903 8996 7288 9024
rect 1903 8993 1915 8996
rect 1857 8987 1915 8993
rect 7282 8984 7288 8996
rect 7340 8984 7346 9036
rect 9769 9027 9827 9033
rect 9769 8993 9781 9027
rect 9815 9024 9827 9027
rect 10042 9024 10048 9036
rect 9815 8996 10048 9024
rect 9815 8993 9827 8996
rect 9769 8987 9827 8993
rect 10042 8984 10048 8996
rect 10100 9024 10106 9036
rect 10778 9024 10784 9036
rect 10100 8996 10784 9024
rect 10100 8984 10106 8996
rect 10778 8984 10784 8996
rect 10836 9024 10842 9036
rect 12618 9024 12624 9036
rect 10836 8996 11468 9024
rect 12579 8996 12624 9024
rect 10836 8984 10842 8996
rect 1578 8956 1584 8968
rect 1539 8928 1584 8956
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 10962 8956 10968 8968
rect 10923 8928 10968 8956
rect 10962 8916 10968 8928
rect 11020 8916 11026 8968
rect 11440 8965 11468 8996
rect 12618 8984 12624 8996
rect 12676 8984 12682 9036
rect 13633 9027 13691 9033
rect 13633 8993 13645 9027
rect 13679 9024 13691 9027
rect 14642 9024 14648 9036
rect 13679 8996 14648 9024
rect 13679 8993 13691 8996
rect 13633 8987 13691 8993
rect 14642 8984 14648 8996
rect 14700 8984 14706 9036
rect 16390 9024 16396 9036
rect 16351 8996 16396 9024
rect 16390 8984 16396 8996
rect 16448 8984 16454 9036
rect 11425 8959 11483 8965
rect 11425 8925 11437 8959
rect 11471 8925 11483 8959
rect 11425 8919 11483 8925
rect 13725 8959 13783 8965
rect 13725 8925 13737 8959
rect 13771 8956 13783 8959
rect 13998 8956 14004 8968
rect 13771 8928 14004 8956
rect 13771 8925 13783 8928
rect 13725 8919 13783 8925
rect 13998 8916 14004 8928
rect 14056 8916 14062 8968
rect 14366 8956 14372 8968
rect 14327 8928 14372 8956
rect 14366 8916 14372 8928
rect 14424 8916 14430 8968
rect 16684 8956 16712 9132
rect 18138 9052 18144 9104
rect 18196 9092 18202 9104
rect 18966 9092 18972 9104
rect 18196 9064 18972 9092
rect 18196 9052 18202 9064
rect 18966 9052 18972 9064
rect 19024 9092 19030 9104
rect 19521 9095 19579 9101
rect 19521 9092 19533 9095
rect 19024 9064 19533 9092
rect 19024 9052 19030 9064
rect 19521 9061 19533 9064
rect 19567 9061 19579 9095
rect 19521 9055 19579 9061
rect 20714 9052 20720 9104
rect 20772 9092 20778 9104
rect 22278 9092 22284 9104
rect 20772 9064 22284 9092
rect 20772 9052 20778 9064
rect 22278 9052 22284 9064
rect 22336 9052 22342 9104
rect 24504 9092 24532 9132
rect 24578 9120 24584 9172
rect 24636 9160 24642 9172
rect 24673 9163 24731 9169
rect 24673 9160 24685 9163
rect 24636 9132 24685 9160
rect 24636 9120 24642 9132
rect 24673 9129 24685 9132
rect 24719 9129 24731 9163
rect 24673 9123 24731 9129
rect 24762 9120 24768 9172
rect 24820 9160 24826 9172
rect 30742 9160 30748 9172
rect 24820 9132 30748 9160
rect 24820 9120 24826 9132
rect 30742 9120 30748 9132
rect 30800 9120 30806 9172
rect 33505 9163 33563 9169
rect 33505 9129 33517 9163
rect 33551 9160 33563 9163
rect 37918 9160 37924 9172
rect 33551 9132 37924 9160
rect 33551 9129 33563 9132
rect 33505 9123 33563 9129
rect 26786 9092 26792 9104
rect 24504 9064 26792 9092
rect 26786 9052 26792 9064
rect 26844 9052 26850 9104
rect 26896 9064 27292 9092
rect 16850 9024 16856 9036
rect 16811 8996 16856 9024
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 17126 8984 17132 9036
rect 17184 9024 17190 9036
rect 18877 9027 18935 9033
rect 18877 9024 18889 9027
rect 17184 8996 18889 9024
rect 17184 8984 17190 8996
rect 18877 8993 18889 8996
rect 18923 9024 18935 9027
rect 20257 9027 20315 9033
rect 18923 8996 19334 9024
rect 18923 8993 18935 8996
rect 18877 8987 18935 8993
rect 15778 8928 16712 8956
rect 10321 8891 10379 8897
rect 10321 8857 10333 8891
rect 10367 8888 10379 8891
rect 11054 8888 11060 8900
rect 10367 8860 11060 8888
rect 10367 8857 10379 8860
rect 10321 8851 10379 8857
rect 11054 8848 11060 8860
rect 11112 8848 11118 8900
rect 12158 8888 12164 8900
rect 12119 8860 12164 8888
rect 12158 8848 12164 8860
rect 12216 8848 12222 8900
rect 12253 8891 12311 8897
rect 12253 8857 12265 8891
rect 12299 8857 12311 8891
rect 12253 8851 12311 8857
rect 10873 8823 10931 8829
rect 10873 8789 10885 8823
rect 10919 8820 10931 8823
rect 12268 8820 12296 8851
rect 14550 8848 14556 8900
rect 14608 8888 14614 8900
rect 14645 8891 14703 8897
rect 14645 8888 14657 8891
rect 14608 8860 14657 8888
rect 14608 8848 14614 8860
rect 14645 8857 14657 8860
rect 14691 8857 14703 8891
rect 14645 8851 14703 8857
rect 17129 8891 17187 8897
rect 17129 8857 17141 8891
rect 17175 8888 17187 8891
rect 17402 8888 17408 8900
rect 17175 8860 17408 8888
rect 17175 8857 17187 8860
rect 17129 8851 17187 8857
rect 17402 8848 17408 8860
rect 17460 8848 17466 8900
rect 18782 8888 18788 8900
rect 18354 8860 18788 8888
rect 18782 8848 18788 8860
rect 18840 8848 18846 8900
rect 10919 8792 12296 8820
rect 10919 8789 10931 8792
rect 10873 8783 10931 8789
rect 12342 8780 12348 8832
rect 12400 8820 12406 8832
rect 18138 8820 18144 8832
rect 12400 8792 18144 8820
rect 12400 8780 12406 8792
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 19306 8820 19334 8996
rect 20257 8993 20269 9027
rect 20303 9024 20315 9027
rect 21082 9024 21088 9036
rect 20303 8996 21088 9024
rect 20303 8993 20315 8996
rect 20257 8987 20315 8993
rect 21082 8984 21088 8996
rect 21140 8984 21146 9036
rect 21634 8984 21640 9036
rect 21692 9024 21698 9036
rect 23569 9027 23627 9033
rect 23569 9024 23581 9027
rect 21692 8996 23581 9024
rect 21692 8984 21698 8996
rect 23569 8993 23581 8996
rect 23615 9024 23627 9027
rect 24302 9024 24308 9036
rect 23615 8996 24308 9024
rect 23615 8993 23627 8996
rect 23569 8987 23627 8993
rect 24302 8984 24308 8996
rect 24360 8984 24366 9036
rect 24394 8984 24400 9036
rect 24452 9024 24458 9036
rect 25777 9027 25835 9033
rect 25777 9024 25789 9027
rect 24452 8996 25789 9024
rect 24452 8984 24458 8996
rect 25777 8993 25789 8996
rect 25823 8993 25835 9027
rect 25777 8987 25835 8993
rect 25866 8984 25872 9036
rect 25924 9024 25930 9036
rect 26053 9027 26111 9033
rect 26053 9024 26065 9027
rect 25924 8996 26065 9024
rect 25924 8984 25930 8996
rect 26053 8993 26065 8996
rect 26099 9024 26111 9027
rect 26896 9024 26924 9064
rect 26099 8996 26924 9024
rect 26973 9027 27031 9033
rect 26099 8993 26111 8996
rect 26053 8987 26111 8993
rect 26973 8993 26985 9027
rect 27019 9024 27031 9027
rect 27154 9024 27160 9036
rect 27019 8996 27160 9024
rect 27019 8993 27031 8996
rect 26973 8987 27031 8993
rect 27154 8984 27160 8996
rect 27212 8984 27218 9036
rect 27264 9033 27292 9064
rect 27706 9052 27712 9104
rect 27764 9092 27770 9104
rect 28813 9095 28871 9101
rect 28813 9092 28825 9095
rect 27764 9064 28825 9092
rect 27764 9052 27770 9064
rect 28813 9061 28825 9064
rect 28859 9061 28871 9095
rect 28813 9055 28871 9061
rect 27249 9027 27307 9033
rect 27249 8993 27261 9027
rect 27295 9024 27307 9027
rect 30558 9024 30564 9036
rect 27295 8996 30564 9024
rect 27295 8993 27307 8996
rect 27249 8987 27307 8993
rect 30558 8984 30564 8996
rect 30616 8984 30622 9036
rect 19610 8956 19616 8968
rect 19571 8928 19616 8956
rect 19610 8916 19616 8928
rect 19668 8916 19674 8968
rect 20162 8956 20168 8968
rect 20123 8928 20168 8956
rect 20162 8916 20168 8928
rect 20220 8916 20226 8968
rect 20809 8959 20867 8965
rect 20809 8925 20821 8959
rect 20855 8956 20867 8959
rect 20990 8956 20996 8968
rect 20855 8928 20996 8956
rect 20855 8925 20867 8928
rect 20809 8919 20867 8925
rect 20990 8916 20996 8928
rect 21048 8956 21054 8968
rect 21545 8959 21603 8965
rect 21545 8956 21557 8959
rect 21048 8928 21557 8956
rect 21048 8916 21054 8928
rect 21545 8925 21557 8928
rect 21591 8925 21603 8959
rect 24762 8956 24768 8968
rect 24723 8928 24768 8956
rect 21545 8919 21603 8925
rect 24762 8916 24768 8928
rect 24820 8916 24826 8968
rect 28077 8959 28135 8965
rect 28077 8956 28089 8959
rect 28000 8928 28089 8956
rect 20530 8848 20536 8900
rect 20588 8888 20594 8900
rect 20714 8888 20720 8900
rect 20588 8860 20720 8888
rect 20588 8848 20594 8860
rect 20714 8848 20720 8860
rect 20772 8848 20778 8900
rect 20898 8888 20904 8900
rect 20859 8860 20904 8888
rect 20898 8848 20904 8860
rect 20956 8848 20962 8900
rect 23198 8888 23204 8900
rect 22862 8860 23204 8888
rect 23198 8848 23204 8860
rect 23256 8848 23262 8900
rect 23293 8891 23351 8897
rect 23293 8857 23305 8891
rect 23339 8857 23351 8891
rect 23293 8851 23351 8857
rect 21726 8820 21732 8832
rect 19306 8792 21732 8820
rect 21726 8780 21732 8792
rect 21784 8780 21790 8832
rect 22278 8780 22284 8832
rect 22336 8820 22342 8832
rect 23308 8820 23336 8851
rect 25130 8848 25136 8900
rect 25188 8888 25194 8900
rect 25869 8891 25927 8897
rect 25869 8888 25881 8891
rect 25188 8860 25881 8888
rect 25188 8848 25194 8860
rect 25869 8857 25881 8860
rect 25915 8857 25927 8891
rect 25869 8851 25927 8857
rect 26510 8848 26516 8900
rect 26568 8888 26574 8900
rect 27065 8891 27123 8897
rect 27065 8888 27077 8891
rect 26568 8860 27077 8888
rect 26568 8848 26574 8860
rect 27065 8857 27077 8860
rect 27111 8857 27123 8891
rect 27065 8851 27123 8857
rect 22336 8792 23336 8820
rect 22336 8780 22342 8792
rect 26602 8780 26608 8832
rect 26660 8820 26666 8832
rect 28000 8820 28028 8928
rect 28077 8925 28089 8928
rect 28123 8925 28135 8959
rect 28077 8919 28135 8925
rect 28166 8916 28172 8968
rect 28224 8956 28230 8968
rect 28905 8959 28963 8965
rect 28224 8928 28269 8956
rect 28224 8916 28230 8928
rect 28905 8925 28917 8959
rect 28951 8956 28963 8959
rect 30190 8956 30196 8968
rect 28951 8928 28985 8956
rect 30103 8928 30196 8956
rect 28951 8925 28963 8928
rect 28905 8919 28963 8925
rect 28810 8848 28816 8900
rect 28868 8888 28874 8900
rect 28920 8888 28948 8919
rect 30190 8916 30196 8928
rect 30248 8956 30254 8968
rect 32493 8959 32551 8965
rect 32493 8956 32505 8959
rect 30248 8928 32505 8956
rect 30248 8916 30254 8928
rect 32493 8925 32505 8928
rect 32539 8925 32551 8959
rect 32493 8919 32551 8925
rect 32861 8959 32919 8965
rect 32861 8925 32873 8959
rect 32907 8956 32919 8959
rect 33042 8956 33048 8968
rect 32907 8928 33048 8956
rect 32907 8925 32919 8928
rect 32861 8919 32919 8925
rect 33042 8916 33048 8928
rect 33100 8956 33106 8968
rect 33520 8956 33548 9123
rect 37918 9120 37924 9132
rect 37976 9120 37982 9172
rect 33100 8928 33548 8956
rect 33100 8916 33106 8928
rect 29917 8891 29975 8897
rect 29917 8888 29929 8891
rect 28868 8860 29929 8888
rect 28868 8848 28874 8860
rect 29917 8857 29929 8860
rect 29963 8857 29975 8891
rect 29917 8851 29975 8857
rect 26660 8792 28028 8820
rect 26660 8780 26666 8792
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 10962 8576 10968 8628
rect 11020 8616 11026 8628
rect 13906 8616 13912 8628
rect 11020 8588 13912 8616
rect 11020 8576 11026 8588
rect 13906 8576 13912 8588
rect 13964 8576 13970 8628
rect 14001 8619 14059 8625
rect 14001 8585 14013 8619
rect 14047 8616 14059 8619
rect 14182 8616 14188 8628
rect 14047 8588 14188 8616
rect 14047 8585 14059 8588
rect 14001 8579 14059 8585
rect 14182 8576 14188 8588
rect 14240 8576 14246 8628
rect 18138 8576 18144 8628
rect 18196 8616 18202 8628
rect 22554 8616 22560 8628
rect 18196 8588 22560 8616
rect 18196 8576 18202 8588
rect 22554 8576 22560 8588
rect 22612 8576 22618 8628
rect 24118 8616 24124 8628
rect 22664 8588 24124 8616
rect 11149 8551 11207 8557
rect 11149 8517 11161 8551
rect 11195 8548 11207 8551
rect 11238 8548 11244 8560
rect 11195 8520 11244 8548
rect 11195 8517 11207 8520
rect 11149 8511 11207 8517
rect 11238 8508 11244 8520
rect 11296 8508 11302 8560
rect 12066 8508 12072 8560
rect 12124 8548 12130 8560
rect 14734 8548 14740 8560
rect 12124 8520 12296 8548
rect 14695 8520 14740 8548
rect 12124 8508 12130 8520
rect 2869 8483 2927 8489
rect 2869 8449 2881 8483
rect 2915 8480 2927 8483
rect 9766 8480 9772 8492
rect 2915 8452 9772 8480
rect 2915 8449 2927 8452
rect 2869 8443 2927 8449
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 12268 8489 12296 8520
rect 14734 8508 14740 8520
rect 14792 8508 14798 8560
rect 18506 8548 18512 8560
rect 15962 8520 18512 8548
rect 18506 8508 18512 8520
rect 18564 8508 18570 8560
rect 22664 8548 22692 8588
rect 24118 8576 24124 8588
rect 24176 8576 24182 8628
rect 24302 8616 24308 8628
rect 24263 8588 24308 8616
rect 24302 8576 24308 8588
rect 24360 8576 24366 8628
rect 24596 8588 26096 8616
rect 24596 8548 24624 8588
rect 19458 8520 22692 8548
rect 23506 8520 24624 8548
rect 24670 8508 24676 8560
rect 24728 8548 24734 8560
rect 25041 8551 25099 8557
rect 25041 8548 25053 8551
rect 24728 8520 25053 8548
rect 24728 8508 24734 8520
rect 25041 8517 25053 8520
rect 25087 8517 25099 8551
rect 25041 8511 25099 8517
rect 25593 8551 25651 8557
rect 25593 8517 25605 8551
rect 25639 8548 25651 8551
rect 25866 8548 25872 8560
rect 25639 8520 25872 8548
rect 25639 8517 25651 8520
rect 25593 8511 25651 8517
rect 25866 8508 25872 8520
rect 25924 8508 25930 8560
rect 26068 8548 26096 8588
rect 27246 8576 27252 8628
rect 27304 8616 27310 8628
rect 27893 8619 27951 8625
rect 27893 8616 27905 8619
rect 27304 8588 27905 8616
rect 27304 8576 27310 8588
rect 27893 8585 27905 8588
rect 27939 8585 27951 8619
rect 27893 8579 27951 8585
rect 27982 8576 27988 8628
rect 28040 8616 28046 8628
rect 28166 8616 28172 8628
rect 28040 8588 28172 8616
rect 28040 8576 28046 8588
rect 28166 8576 28172 8588
rect 28224 8616 28230 8628
rect 28902 8616 28908 8628
rect 28224 8588 28908 8616
rect 28224 8576 28230 8588
rect 28902 8576 28908 8588
rect 28960 8576 28966 8628
rect 29178 8616 29184 8628
rect 29139 8588 29184 8616
rect 29178 8576 29184 8588
rect 29236 8576 29242 8628
rect 29822 8548 29828 8560
rect 26068 8520 29828 8548
rect 29822 8508 29828 8520
rect 29880 8508 29886 8560
rect 38010 8548 38016 8560
rect 37971 8520 38016 8548
rect 38010 8508 38016 8520
rect 38068 8508 38074 8560
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8449 12311 8483
rect 14090 8480 14096 8492
rect 13662 8452 14096 8480
rect 12253 8443 12311 8449
rect 14090 8440 14096 8452
rect 14148 8440 14154 8492
rect 17310 8480 17316 8492
rect 17271 8452 17316 8480
rect 17310 8440 17316 8452
rect 17368 8440 17374 8492
rect 19978 8480 19984 8492
rect 19939 8452 19984 8480
rect 19978 8440 19984 8452
rect 20036 8440 20042 8492
rect 20625 8483 20683 8489
rect 20625 8449 20637 8483
rect 20671 8480 20683 8483
rect 20806 8480 20812 8492
rect 20671 8452 20812 8480
rect 20671 8449 20683 8452
rect 20625 8443 20683 8449
rect 20806 8440 20812 8452
rect 20864 8440 20870 8492
rect 21174 8480 21180 8492
rect 21135 8452 21180 8480
rect 21174 8440 21180 8452
rect 21232 8440 21238 8492
rect 21269 8483 21327 8489
rect 21269 8449 21281 8483
rect 21315 8449 21327 8483
rect 21269 8443 21327 8449
rect 10597 8415 10655 8421
rect 10597 8381 10609 8415
rect 10643 8412 10655 8415
rect 11054 8412 11060 8424
rect 10643 8384 11060 8412
rect 10643 8381 10655 8384
rect 10597 8375 10655 8381
rect 11054 8372 11060 8384
rect 11112 8412 11118 8424
rect 11701 8415 11759 8421
rect 11701 8412 11713 8415
rect 11112 8384 11713 8412
rect 11112 8372 11118 8384
rect 11701 8381 11713 8384
rect 11747 8412 11759 8415
rect 12066 8412 12072 8424
rect 11747 8384 12072 8412
rect 11747 8381 11759 8384
rect 11701 8375 11759 8381
rect 12066 8372 12072 8384
rect 12124 8372 12130 8424
rect 12526 8412 12532 8424
rect 12487 8384 12532 8412
rect 12526 8372 12532 8384
rect 12584 8372 12590 8424
rect 14458 8412 14464 8424
rect 14419 8384 14464 8412
rect 14458 8372 14464 8384
rect 14516 8372 14522 8424
rect 17957 8415 18015 8421
rect 17957 8381 17969 8415
rect 18003 8381 18015 8415
rect 17957 8375 18015 8381
rect 18233 8415 18291 8421
rect 18233 8381 18245 8415
rect 18279 8412 18291 8415
rect 20533 8415 20591 8421
rect 18279 8384 20484 8412
rect 18279 8381 18291 8384
rect 18233 8375 18291 8381
rect 2774 8304 2780 8356
rect 2832 8344 2838 8356
rect 2832 8316 2877 8344
rect 2832 8304 2838 8316
rect 15746 8304 15752 8356
rect 15804 8344 15810 8356
rect 16209 8347 16267 8353
rect 16209 8344 16221 8347
rect 15804 8316 16221 8344
rect 15804 8304 15810 8316
rect 16209 8313 16221 8316
rect 16255 8313 16267 8347
rect 17494 8344 17500 8356
rect 17455 8316 17500 8344
rect 16209 8307 16267 8313
rect 17494 8304 17500 8316
rect 17552 8304 17558 8356
rect 13906 8236 13912 8288
rect 13964 8276 13970 8288
rect 15286 8276 15292 8288
rect 13964 8248 15292 8276
rect 13964 8236 13970 8248
rect 15286 8236 15292 8248
rect 15344 8276 15350 8288
rect 16022 8276 16028 8288
rect 15344 8248 16028 8276
rect 15344 8236 15350 8248
rect 16022 8236 16028 8248
rect 16080 8236 16086 8288
rect 17972 8276 18000 8375
rect 19242 8304 19248 8356
rect 19300 8344 19306 8356
rect 20456 8344 20484 8384
rect 20533 8381 20545 8415
rect 20579 8412 20591 8415
rect 20714 8412 20720 8424
rect 20579 8384 20720 8412
rect 20579 8381 20591 8384
rect 20533 8375 20591 8381
rect 20714 8372 20720 8384
rect 20772 8372 20778 8424
rect 20898 8372 20904 8424
rect 20956 8412 20962 8424
rect 21284 8412 21312 8443
rect 21634 8440 21640 8492
rect 21692 8480 21698 8492
rect 22005 8483 22063 8489
rect 22005 8480 22017 8483
rect 21692 8452 22017 8480
rect 21692 8440 21698 8452
rect 22005 8449 22017 8452
rect 22051 8449 22063 8483
rect 24762 8480 24768 8492
rect 22005 8443 22063 8449
rect 23492 8452 24768 8480
rect 22278 8412 22284 8424
rect 20956 8384 21312 8412
rect 22239 8384 22284 8412
rect 20956 8372 20962 8384
rect 22278 8372 22284 8384
rect 22336 8372 22342 8424
rect 22646 8372 22652 8424
rect 22704 8412 22710 8424
rect 23492 8412 23520 8452
rect 24762 8440 24768 8452
rect 24820 8440 24826 8492
rect 25774 8440 25780 8492
rect 25832 8480 25838 8492
rect 25958 8480 25964 8492
rect 25832 8452 25964 8480
rect 25832 8440 25838 8452
rect 25958 8440 25964 8452
rect 26016 8480 26022 8492
rect 26053 8483 26111 8489
rect 26053 8480 26065 8483
rect 26016 8452 26065 8480
rect 26016 8440 26022 8452
rect 26053 8449 26065 8452
rect 26099 8449 26111 8483
rect 26053 8443 26111 8449
rect 26418 8440 26424 8492
rect 26476 8480 26482 8492
rect 27341 8483 27399 8489
rect 27341 8480 27353 8483
rect 26476 8452 27353 8480
rect 26476 8440 26482 8452
rect 27341 8449 27353 8452
rect 27387 8480 27399 8483
rect 27614 8480 27620 8492
rect 27387 8452 27620 8480
rect 27387 8449 27399 8452
rect 27341 8443 27399 8449
rect 27614 8440 27620 8452
rect 27672 8440 27678 8492
rect 27982 8480 27988 8492
rect 27943 8452 27988 8480
rect 27982 8440 27988 8452
rect 28040 8440 28046 8492
rect 28626 8480 28632 8492
rect 28587 8452 28632 8480
rect 28626 8440 28632 8452
rect 28684 8440 28690 8492
rect 28902 8440 28908 8492
rect 28960 8480 28966 8492
rect 29089 8483 29147 8489
rect 29089 8480 29101 8483
rect 28960 8452 29101 8480
rect 28960 8440 28966 8452
rect 29089 8449 29101 8452
rect 29135 8449 29147 8483
rect 29089 8443 29147 8449
rect 29917 8483 29975 8489
rect 29917 8449 29929 8483
rect 29963 8480 29975 8483
rect 30006 8480 30012 8492
rect 29963 8452 30012 8480
rect 29963 8449 29975 8452
rect 29917 8443 29975 8449
rect 30006 8440 30012 8452
rect 30064 8480 30070 8492
rect 30561 8483 30619 8489
rect 30561 8480 30573 8483
rect 30064 8452 30573 8480
rect 30064 8440 30070 8452
rect 30561 8449 30573 8452
rect 30607 8449 30619 8483
rect 30561 8443 30619 8449
rect 37553 8483 37611 8489
rect 37553 8449 37565 8483
rect 37599 8480 37611 8483
rect 38194 8480 38200 8492
rect 37599 8452 38200 8480
rect 37599 8449 37611 8452
rect 37553 8443 37611 8449
rect 38194 8440 38200 8452
rect 38252 8440 38258 8492
rect 22704 8384 23520 8412
rect 22704 8372 22710 8384
rect 23658 8372 23664 8424
rect 23716 8412 23722 8424
rect 23753 8415 23811 8421
rect 23753 8412 23765 8415
rect 23716 8384 23765 8412
rect 23716 8372 23722 8384
rect 23753 8381 23765 8384
rect 23799 8412 23811 8415
rect 23934 8412 23940 8424
rect 23799 8384 23940 8412
rect 23799 8381 23811 8384
rect 23753 8375 23811 8381
rect 23934 8372 23940 8384
rect 23992 8372 23998 8424
rect 24486 8372 24492 8424
rect 24544 8412 24550 8424
rect 24949 8415 25007 8421
rect 24949 8412 24961 8415
rect 24544 8384 24961 8412
rect 24544 8372 24550 8384
rect 24949 8381 24961 8384
rect 24995 8381 25007 8415
rect 28537 8415 28595 8421
rect 28537 8412 28549 8415
rect 24949 8375 25007 8381
rect 25056 8384 28549 8412
rect 22002 8344 22008 8356
rect 19300 8316 19472 8344
rect 20456 8316 22008 8344
rect 19300 8304 19306 8316
rect 19334 8276 19340 8288
rect 17972 8248 19340 8276
rect 19334 8236 19340 8248
rect 19392 8236 19398 8288
rect 19444 8276 19472 8316
rect 22002 8304 22008 8316
rect 22060 8304 22066 8356
rect 23290 8304 23296 8356
rect 23348 8344 23354 8356
rect 23348 8316 24716 8344
rect 23348 8304 23354 8316
rect 22370 8276 22376 8288
rect 19444 8248 22376 8276
rect 22370 8236 22376 8248
rect 22428 8236 22434 8288
rect 24688 8276 24716 8316
rect 24762 8304 24768 8356
rect 24820 8344 24826 8356
rect 25056 8344 25084 8384
rect 28537 8381 28549 8384
rect 28583 8381 28595 8415
rect 28537 8375 28595 8381
rect 28718 8372 28724 8424
rect 28776 8412 28782 8424
rect 29825 8415 29883 8421
rect 29825 8412 29837 8415
rect 28776 8384 29837 8412
rect 28776 8372 28782 8384
rect 29825 8381 29837 8384
rect 29871 8381 29883 8415
rect 29825 8375 29883 8381
rect 27249 8347 27307 8353
rect 27249 8344 27261 8347
rect 24820 8316 25084 8344
rect 25608 8316 27261 8344
rect 24820 8304 24826 8316
rect 25608 8276 25636 8316
rect 27249 8313 27261 8316
rect 27295 8313 27307 8347
rect 27249 8307 27307 8313
rect 28994 8304 29000 8356
rect 29052 8344 29058 8356
rect 30469 8347 30527 8353
rect 30469 8344 30481 8347
rect 29052 8316 30481 8344
rect 29052 8304 29058 8316
rect 30469 8313 30481 8316
rect 30515 8313 30527 8347
rect 30469 8307 30527 8313
rect 24688 8248 25636 8276
rect 26145 8279 26203 8285
rect 26145 8245 26157 8279
rect 26191 8276 26203 8279
rect 26234 8276 26240 8288
rect 26191 8248 26240 8276
rect 26191 8245 26203 8248
rect 26145 8239 26203 8245
rect 26234 8236 26240 8248
rect 26292 8236 26298 8288
rect 26878 8236 26884 8288
rect 26936 8276 26942 8288
rect 29914 8276 29920 8288
rect 26936 8248 29920 8276
rect 26936 8236 26942 8248
rect 29914 8236 29920 8248
rect 29972 8236 29978 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 10226 8032 10232 8084
rect 10284 8072 10290 8084
rect 10873 8075 10931 8081
rect 10873 8072 10885 8075
rect 10284 8044 10885 8072
rect 10284 8032 10290 8044
rect 10873 8041 10885 8044
rect 10919 8072 10931 8075
rect 12066 8072 12072 8084
rect 10919 8044 12072 8072
rect 10919 8041 10931 8044
rect 10873 8035 10931 8041
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 12250 8032 12256 8084
rect 12308 8072 12314 8084
rect 12621 8075 12679 8081
rect 12621 8072 12633 8075
rect 12308 8044 12633 8072
rect 12308 8032 12314 8044
rect 12621 8041 12633 8044
rect 12667 8041 12679 8075
rect 13262 8072 13268 8084
rect 13223 8044 13268 8072
rect 12621 8035 12679 8041
rect 13262 8032 13268 8044
rect 13320 8032 13326 8084
rect 16301 8075 16359 8081
rect 16301 8072 16313 8075
rect 14200 8044 16313 8072
rect 10594 7896 10600 7948
rect 10652 7936 10658 7948
rect 14200 7936 14228 8044
rect 16301 8041 16313 8044
rect 16347 8072 16359 8075
rect 17034 8072 17040 8084
rect 16347 8044 17040 8072
rect 16347 8041 16359 8044
rect 16301 8035 16359 8041
rect 17034 8032 17040 8044
rect 17092 8032 17098 8084
rect 17770 8032 17776 8084
rect 17828 8072 17834 8084
rect 18785 8075 18843 8081
rect 17828 8044 18736 8072
rect 17828 8032 17834 8044
rect 18708 8004 18736 8044
rect 18785 8041 18797 8075
rect 18831 8072 18843 8075
rect 21818 8072 21824 8084
rect 18831 8044 21824 8072
rect 18831 8041 18843 8044
rect 18785 8035 18843 8041
rect 21818 8032 21824 8044
rect 21876 8032 21882 8084
rect 22002 8032 22008 8084
rect 22060 8072 22066 8084
rect 24762 8072 24768 8084
rect 22060 8044 24768 8072
rect 22060 8032 22066 8044
rect 24762 8032 24768 8044
rect 24820 8032 24826 8084
rect 24857 8075 24915 8081
rect 24857 8041 24869 8075
rect 24903 8072 24915 8075
rect 25038 8072 25044 8084
rect 24903 8044 25044 8072
rect 24903 8041 24915 8044
rect 24857 8035 24915 8041
rect 25038 8032 25044 8044
rect 25096 8032 25102 8084
rect 25501 8075 25559 8081
rect 25501 8041 25513 8075
rect 25547 8072 25559 8075
rect 25590 8072 25596 8084
rect 25547 8044 25596 8072
rect 25547 8041 25559 8044
rect 25501 8035 25559 8041
rect 25590 8032 25596 8044
rect 25648 8032 25654 8084
rect 26050 8032 26056 8084
rect 26108 8072 26114 8084
rect 26145 8075 26203 8081
rect 26145 8072 26157 8075
rect 26108 8044 26157 8072
rect 26108 8032 26114 8044
rect 26145 8041 26157 8044
rect 26191 8041 26203 8075
rect 26786 8072 26792 8084
rect 26747 8044 26792 8072
rect 26145 8035 26203 8041
rect 26786 8032 26792 8044
rect 26844 8032 26850 8084
rect 27522 8032 27528 8084
rect 27580 8072 27586 8084
rect 28077 8075 28135 8081
rect 28077 8072 28089 8075
rect 27580 8044 28089 8072
rect 27580 8032 27586 8044
rect 28077 8041 28089 8044
rect 28123 8041 28135 8075
rect 28077 8035 28135 8041
rect 30282 8032 30288 8084
rect 30340 8072 30346 8084
rect 30469 8075 30527 8081
rect 30469 8072 30481 8075
rect 30340 8044 30481 8072
rect 30340 8032 30346 8044
rect 30469 8041 30481 8044
rect 30515 8041 30527 8075
rect 30469 8035 30527 8041
rect 19242 8004 19248 8016
rect 18708 7976 19248 8004
rect 19242 7964 19248 7976
rect 19300 7964 19306 8016
rect 21082 7964 21088 8016
rect 21140 8004 21146 8016
rect 21140 7976 21864 8004
rect 21140 7964 21146 7976
rect 10652 7908 14228 7936
rect 17037 7939 17095 7945
rect 10652 7896 10658 7908
rect 17037 7905 17049 7939
rect 17083 7936 17095 7939
rect 19334 7936 19340 7948
rect 17083 7908 19340 7936
rect 17083 7905 17095 7908
rect 17037 7899 17095 7905
rect 19334 7896 19340 7908
rect 19392 7936 19398 7948
rect 19429 7939 19487 7945
rect 19429 7936 19441 7939
rect 19392 7908 19441 7936
rect 19392 7896 19398 7908
rect 19429 7905 19441 7908
rect 19475 7936 19487 7939
rect 21634 7936 21640 7948
rect 19475 7908 21640 7936
rect 19475 7905 19487 7908
rect 19429 7899 19487 7905
rect 21634 7896 21640 7908
rect 21692 7936 21698 7948
rect 21729 7939 21787 7945
rect 21729 7936 21741 7939
rect 21692 7908 21741 7936
rect 21692 7896 21698 7908
rect 21729 7905 21741 7908
rect 21775 7905 21787 7939
rect 21836 7936 21864 7976
rect 23198 7964 23204 8016
rect 23256 8004 23262 8016
rect 29825 8007 29883 8013
rect 29825 8004 29837 8007
rect 23256 7976 29837 8004
rect 23256 7964 23262 7976
rect 29825 7973 29837 7976
rect 29871 7973 29883 8007
rect 29825 7967 29883 7973
rect 24026 7936 24032 7948
rect 21836 7908 24032 7936
rect 21729 7899 21787 7905
rect 24026 7896 24032 7908
rect 24084 7896 24090 7948
rect 25608 7908 27384 7936
rect 3326 7828 3332 7880
rect 3384 7868 3390 7880
rect 12713 7871 12771 7877
rect 3384 7840 12434 7868
rect 3384 7828 3390 7840
rect 12406 7800 12434 7840
rect 12713 7837 12725 7871
rect 12759 7868 12771 7871
rect 13262 7868 13268 7880
rect 12759 7840 13268 7868
rect 12759 7837 12771 7840
rect 12713 7831 12771 7837
rect 13262 7828 13268 7840
rect 13320 7828 13326 7880
rect 13357 7871 13415 7877
rect 13357 7837 13369 7871
rect 13403 7868 13415 7871
rect 14090 7868 14096 7880
rect 13403 7840 14096 7868
rect 13403 7837 13415 7840
rect 13357 7831 13415 7837
rect 14090 7828 14096 7840
rect 14148 7828 14154 7880
rect 14550 7868 14556 7880
rect 14511 7840 14556 7868
rect 14550 7828 14556 7840
rect 14608 7828 14614 7880
rect 18782 7828 18788 7880
rect 18840 7868 18846 7880
rect 18840 7840 19472 7868
rect 18840 7828 18846 7840
rect 12618 7800 12624 7812
rect 12406 7772 12624 7800
rect 12618 7760 12624 7772
rect 12676 7760 12682 7812
rect 14829 7803 14887 7809
rect 14829 7769 14841 7803
rect 14875 7769 14887 7803
rect 16054 7772 17264 7800
rect 14829 7763 14887 7769
rect 11054 7692 11060 7744
rect 11112 7732 11118 7744
rect 11425 7735 11483 7741
rect 11425 7732 11437 7735
rect 11112 7704 11437 7732
rect 11112 7692 11118 7704
rect 11425 7701 11437 7704
rect 11471 7732 11483 7735
rect 11977 7735 12035 7741
rect 11977 7732 11989 7735
rect 11471 7704 11989 7732
rect 11471 7701 11483 7704
rect 11425 7695 11483 7701
rect 11977 7701 11989 7704
rect 12023 7701 12035 7735
rect 11977 7695 12035 7701
rect 12066 7692 12072 7744
rect 12124 7732 12130 7744
rect 14844 7732 14872 7763
rect 17126 7732 17132 7744
rect 12124 7704 17132 7732
rect 12124 7692 12130 7704
rect 17126 7692 17132 7704
rect 17184 7692 17190 7744
rect 17236 7732 17264 7772
rect 17310 7760 17316 7812
rect 17368 7800 17374 7812
rect 19444 7800 19472 7840
rect 23750 7828 23756 7880
rect 23808 7868 23814 7880
rect 25608 7877 25636 7908
rect 24765 7871 24823 7877
rect 24765 7868 24777 7871
rect 23808 7840 24777 7868
rect 23808 7828 23814 7840
rect 24765 7837 24777 7840
rect 24811 7837 24823 7871
rect 24765 7831 24823 7837
rect 25593 7871 25651 7877
rect 25593 7837 25605 7871
rect 25639 7837 25651 7871
rect 26234 7868 26240 7880
rect 26147 7840 26240 7868
rect 25593 7831 25651 7837
rect 26234 7828 26240 7840
rect 26292 7868 26298 7880
rect 26878 7868 26884 7880
rect 26292 7840 26884 7868
rect 26292 7828 26298 7840
rect 26878 7828 26884 7840
rect 26936 7828 26942 7880
rect 27246 7828 27252 7880
rect 27304 7828 27310 7880
rect 19705 7803 19763 7809
rect 19705 7800 19717 7803
rect 17368 7772 17413 7800
rect 18538 7772 19380 7800
rect 19444 7772 19717 7800
rect 17368 7760 17374 7772
rect 18690 7732 18696 7744
rect 17236 7704 18696 7732
rect 18690 7692 18696 7704
rect 18748 7692 18754 7744
rect 19352 7732 19380 7772
rect 19705 7769 19717 7772
rect 19751 7769 19763 7803
rect 21266 7800 21272 7812
rect 20930 7772 21272 7800
rect 19705 7763 19763 7769
rect 21266 7760 21272 7772
rect 21324 7760 21330 7812
rect 21726 7760 21732 7812
rect 21784 7800 21790 7812
rect 22005 7803 22063 7809
rect 22005 7800 22017 7803
rect 21784 7772 22017 7800
rect 21784 7760 21790 7772
rect 22005 7769 22017 7772
rect 22051 7769 22063 7803
rect 27264 7800 27292 7828
rect 23230 7772 27292 7800
rect 27356 7800 27384 7908
rect 27430 7896 27436 7948
rect 27488 7936 27494 7948
rect 28721 7939 28779 7945
rect 28721 7936 28733 7939
rect 27488 7908 28733 7936
rect 27488 7896 27494 7908
rect 28721 7905 28733 7908
rect 28767 7905 28779 7939
rect 28721 7899 28779 7905
rect 27525 7871 27583 7877
rect 27525 7837 27537 7871
rect 27571 7868 27583 7871
rect 28074 7868 28080 7880
rect 27571 7840 28080 7868
rect 27571 7837 27583 7840
rect 27525 7831 27583 7837
rect 28074 7828 28080 7840
rect 28132 7828 28138 7880
rect 28166 7828 28172 7880
rect 28224 7868 28230 7880
rect 28810 7868 28816 7880
rect 28224 7840 28269 7868
rect 28771 7840 28816 7868
rect 28224 7828 28230 7840
rect 28810 7828 28816 7840
rect 28868 7828 28874 7880
rect 29917 7871 29975 7877
rect 29917 7837 29929 7871
rect 29963 7868 29975 7871
rect 30006 7868 30012 7880
rect 29963 7840 30012 7868
rect 29963 7837 29975 7840
rect 29917 7831 29975 7837
rect 30006 7828 30012 7840
rect 30064 7828 30070 7880
rect 30282 7828 30288 7880
rect 30340 7868 30346 7880
rect 30561 7871 30619 7877
rect 30561 7868 30573 7871
rect 30340 7840 30573 7868
rect 30340 7828 30346 7840
rect 30561 7837 30573 7840
rect 30607 7837 30619 7871
rect 30561 7831 30619 7837
rect 27356 7772 27936 7800
rect 22005 7763 22063 7769
rect 20714 7732 20720 7744
rect 19352 7704 20720 7732
rect 20714 7692 20720 7704
rect 20772 7692 20778 7744
rect 21082 7692 21088 7744
rect 21140 7732 21146 7744
rect 21177 7735 21235 7741
rect 21177 7732 21189 7735
rect 21140 7704 21189 7732
rect 21140 7692 21146 7704
rect 21177 7701 21189 7704
rect 21223 7701 21235 7735
rect 21177 7695 21235 7701
rect 22186 7692 22192 7744
rect 22244 7732 22250 7744
rect 23477 7735 23535 7741
rect 23477 7732 23489 7735
rect 22244 7704 23489 7732
rect 22244 7692 22250 7704
rect 23477 7701 23489 7704
rect 23523 7701 23535 7735
rect 23477 7695 23535 7701
rect 24118 7692 24124 7744
rect 24176 7732 24182 7744
rect 27246 7732 27252 7744
rect 24176 7704 27252 7732
rect 24176 7692 24182 7704
rect 27246 7692 27252 7704
rect 27304 7692 27310 7744
rect 27430 7732 27436 7744
rect 27391 7704 27436 7732
rect 27430 7692 27436 7704
rect 27488 7692 27494 7744
rect 27908 7732 27936 7772
rect 28442 7732 28448 7744
rect 27908 7704 28448 7732
rect 28442 7692 28448 7704
rect 28500 7692 28506 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 13078 7488 13084 7540
rect 13136 7528 13142 7540
rect 13265 7531 13323 7537
rect 13265 7528 13277 7531
rect 13136 7500 13277 7528
rect 13136 7488 13142 7500
rect 13265 7497 13277 7500
rect 13311 7497 13323 7531
rect 13265 7491 13323 7497
rect 15378 7488 15384 7540
rect 15436 7528 15442 7540
rect 16945 7531 17003 7537
rect 16945 7528 16957 7531
rect 15436 7500 16957 7528
rect 15436 7488 15442 7500
rect 16945 7497 16957 7500
rect 16991 7497 17003 7531
rect 16945 7491 17003 7497
rect 17589 7531 17647 7537
rect 17589 7497 17601 7531
rect 17635 7528 17647 7531
rect 17678 7528 17684 7540
rect 17635 7500 17684 7528
rect 17635 7497 17647 7500
rect 17589 7491 17647 7497
rect 17678 7488 17684 7500
rect 17736 7488 17742 7540
rect 18230 7528 18236 7540
rect 18191 7500 18236 7528
rect 18230 7488 18236 7500
rect 18288 7488 18294 7540
rect 18690 7488 18696 7540
rect 18748 7528 18754 7540
rect 22002 7528 22008 7540
rect 18748 7500 22008 7528
rect 18748 7488 18754 7500
rect 22002 7488 22008 7500
rect 22060 7488 22066 7540
rect 23753 7531 23811 7537
rect 23753 7497 23765 7531
rect 23799 7528 23811 7531
rect 23842 7528 23848 7540
rect 23799 7500 23848 7528
rect 23799 7497 23811 7500
rect 23753 7491 23811 7497
rect 23842 7488 23848 7500
rect 23900 7528 23906 7540
rect 25314 7528 25320 7540
rect 23900 7500 25320 7528
rect 23900 7488 23906 7500
rect 25314 7488 25320 7500
rect 25372 7488 25378 7540
rect 25682 7528 25688 7540
rect 25643 7500 25688 7528
rect 25682 7488 25688 7500
rect 25740 7488 25746 7540
rect 26326 7528 26332 7540
rect 26287 7500 26332 7528
rect 26326 7488 26332 7500
rect 26384 7488 26390 7540
rect 27246 7488 27252 7540
rect 27304 7528 27310 7540
rect 28537 7531 28595 7537
rect 28537 7528 28549 7531
rect 27304 7500 28549 7528
rect 27304 7488 27310 7500
rect 28537 7497 28549 7500
rect 28583 7497 28595 7531
rect 28537 7491 28595 7497
rect 28626 7488 28632 7540
rect 28684 7488 28690 7540
rect 29822 7528 29828 7540
rect 29783 7500 29828 7528
rect 29822 7488 29828 7500
rect 29880 7488 29886 7540
rect 1854 7460 1860 7472
rect 1815 7432 1860 7460
rect 1854 7420 1860 7432
rect 1912 7420 1918 7472
rect 10597 7463 10655 7469
rect 10597 7429 10609 7463
rect 10643 7460 10655 7463
rect 14737 7463 14795 7469
rect 14737 7460 14749 7463
rect 10643 7432 14749 7460
rect 10643 7429 10655 7432
rect 10597 7423 10655 7429
rect 14737 7429 14749 7432
rect 14783 7460 14795 7463
rect 15010 7460 15016 7472
rect 14783 7432 15016 7460
rect 14783 7429 14795 7432
rect 14737 7423 14795 7429
rect 15010 7420 15016 7432
rect 15068 7420 15074 7472
rect 16114 7460 16120 7472
rect 15962 7432 16120 7460
rect 16114 7420 16120 7432
rect 16172 7420 16178 7472
rect 17310 7460 17316 7472
rect 16316 7432 17316 7460
rect 1578 7352 1584 7404
rect 1636 7392 1642 7404
rect 1673 7395 1731 7401
rect 1673 7392 1685 7395
rect 1636 7364 1685 7392
rect 1636 7352 1642 7364
rect 1673 7361 1685 7364
rect 1719 7361 1731 7395
rect 13354 7392 13360 7404
rect 13315 7364 13360 7392
rect 1673 7355 1731 7361
rect 13354 7352 13360 7364
rect 13412 7352 13418 7404
rect 14274 7392 14280 7404
rect 13924 7364 14280 7392
rect 11790 7284 11796 7336
rect 11848 7324 11854 7336
rect 13924 7324 13952 7364
rect 14274 7352 14280 7364
rect 14332 7352 14338 7404
rect 11848 7296 13952 7324
rect 14001 7327 14059 7333
rect 11848 7284 11854 7296
rect 14001 7293 14013 7327
rect 14047 7324 14059 7327
rect 14458 7324 14464 7336
rect 14047 7296 14464 7324
rect 14047 7293 14059 7296
rect 14001 7287 14059 7293
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 16316 7324 16344 7432
rect 17310 7420 17316 7432
rect 17368 7420 17374 7472
rect 19334 7460 19340 7472
rect 18800 7432 19340 7460
rect 17037 7395 17095 7401
rect 17037 7361 17049 7395
rect 17083 7392 17095 7395
rect 17402 7392 17408 7404
rect 17083 7364 17408 7392
rect 17083 7361 17095 7364
rect 17037 7355 17095 7361
rect 17402 7352 17408 7364
rect 17460 7352 17466 7404
rect 17497 7395 17555 7401
rect 17497 7361 17509 7395
rect 17543 7392 17555 7395
rect 17678 7392 17684 7404
rect 17543 7364 17684 7392
rect 17543 7361 17555 7364
rect 17497 7355 17555 7361
rect 14568 7296 16344 7324
rect 12713 7259 12771 7265
rect 12713 7225 12725 7259
rect 12759 7256 12771 7259
rect 13814 7256 13820 7268
rect 12759 7228 13820 7256
rect 12759 7225 12771 7228
rect 12713 7219 12771 7225
rect 13814 7216 13820 7228
rect 13872 7256 13878 7268
rect 14568 7256 14596 7296
rect 16850 7284 16856 7336
rect 16908 7324 16914 7336
rect 17512 7324 17540 7355
rect 17678 7352 17684 7364
rect 17736 7352 17742 7404
rect 17862 7352 17868 7404
rect 17920 7392 17926 7404
rect 18800 7401 18828 7432
rect 19334 7420 19340 7432
rect 19392 7420 19398 7472
rect 22554 7460 22560 7472
rect 20286 7432 22560 7460
rect 22554 7420 22560 7432
rect 22612 7420 22618 7472
rect 24210 7420 24216 7472
rect 24268 7460 24274 7472
rect 25590 7460 25596 7472
rect 24268 7432 25596 7460
rect 24268 7420 24274 7432
rect 25590 7420 25596 7432
rect 25648 7420 25654 7472
rect 27890 7460 27896 7472
rect 27851 7432 27896 7460
rect 27890 7420 27896 7432
rect 27948 7420 27954 7472
rect 28644 7460 28672 7488
rect 29178 7460 29184 7472
rect 28000 7432 28672 7460
rect 29139 7432 29184 7460
rect 18325 7395 18383 7401
rect 18325 7392 18337 7395
rect 17920 7364 18337 7392
rect 17920 7352 17926 7364
rect 18325 7361 18337 7364
rect 18371 7361 18383 7395
rect 18325 7355 18383 7361
rect 18785 7395 18843 7401
rect 18785 7361 18797 7395
rect 18831 7361 18843 7395
rect 18785 7355 18843 7361
rect 16908 7296 17540 7324
rect 16908 7284 16914 7296
rect 17770 7284 17776 7336
rect 17828 7324 17834 7336
rect 18800 7324 18828 7355
rect 21174 7352 21180 7404
rect 21232 7392 21238 7404
rect 21453 7395 21511 7401
rect 21453 7392 21465 7395
rect 21232 7364 21465 7392
rect 21232 7352 21238 7364
rect 21453 7361 21465 7364
rect 21499 7392 21511 7395
rect 21634 7392 21640 7404
rect 21499 7364 21640 7392
rect 21499 7361 21511 7364
rect 21453 7355 21511 7361
rect 21634 7352 21640 7364
rect 21692 7392 21698 7404
rect 22005 7395 22063 7401
rect 22005 7392 22017 7395
rect 21692 7364 22017 7392
rect 21692 7352 21698 7364
rect 22005 7361 22017 7364
rect 22051 7361 22063 7395
rect 22005 7355 22063 7361
rect 23382 7352 23388 7404
rect 23440 7352 23446 7404
rect 24489 7395 24547 7401
rect 24489 7361 24501 7395
rect 24535 7392 24547 7395
rect 25133 7395 25191 7401
rect 25133 7392 25145 7395
rect 24535 7364 25145 7392
rect 24535 7361 24547 7364
rect 24489 7355 24547 7361
rect 25133 7361 25145 7364
rect 25179 7361 25191 7395
rect 25133 7355 25191 7361
rect 25777 7395 25835 7401
rect 25777 7361 25789 7395
rect 25823 7390 25835 7395
rect 26234 7392 26240 7404
rect 25884 7390 26240 7392
rect 25823 7364 26240 7390
rect 25823 7362 25912 7364
rect 25823 7361 25835 7362
rect 25777 7355 25835 7361
rect 17828 7296 18828 7324
rect 19061 7327 19119 7333
rect 17828 7284 17834 7296
rect 19061 7293 19073 7327
rect 19107 7324 19119 7327
rect 19610 7324 19616 7336
rect 19107 7296 19616 7324
rect 19107 7293 19119 7296
rect 19061 7287 19119 7293
rect 19610 7284 19616 7296
rect 19668 7284 19674 7336
rect 20254 7284 20260 7336
rect 20312 7324 20318 7336
rect 20533 7327 20591 7333
rect 20533 7324 20545 7327
rect 20312 7296 20545 7324
rect 20312 7284 20318 7296
rect 20533 7293 20545 7296
rect 20579 7293 20591 7327
rect 20533 7287 20591 7293
rect 22281 7327 22339 7333
rect 22281 7293 22293 7327
rect 22327 7324 22339 7327
rect 22370 7324 22376 7336
rect 22327 7296 22376 7324
rect 22327 7293 22339 7296
rect 22281 7287 22339 7293
rect 22370 7284 22376 7296
rect 22428 7284 22434 7336
rect 22646 7284 22652 7336
rect 22704 7324 22710 7336
rect 25148 7324 25176 7355
rect 26234 7352 26240 7364
rect 26292 7352 26298 7404
rect 26418 7392 26424 7404
rect 26379 7364 26424 7392
rect 26418 7352 26424 7364
rect 26476 7352 26482 7404
rect 27341 7395 27399 7401
rect 27341 7361 27353 7395
rect 27387 7392 27399 7395
rect 27522 7392 27528 7404
rect 27387 7364 27528 7392
rect 27387 7361 27399 7364
rect 27341 7355 27399 7361
rect 27522 7352 27528 7364
rect 27580 7392 27586 7404
rect 28000 7401 28028 7432
rect 29178 7420 29184 7432
rect 29236 7420 29242 7472
rect 27985 7395 28043 7401
rect 27985 7392 27997 7395
rect 27580 7364 27997 7392
rect 27580 7352 27586 7364
rect 27985 7361 27997 7364
rect 28031 7361 28043 7395
rect 27985 7355 28043 7361
rect 28074 7352 28080 7404
rect 28132 7392 28138 7404
rect 28629 7395 28687 7401
rect 28629 7392 28641 7395
rect 28132 7364 28641 7392
rect 28132 7352 28138 7364
rect 28629 7361 28641 7364
rect 28675 7392 28687 7395
rect 28810 7392 28816 7404
rect 28675 7364 28816 7392
rect 28675 7361 28687 7364
rect 28629 7355 28687 7361
rect 28810 7352 28816 7364
rect 28868 7352 28874 7404
rect 29273 7395 29331 7401
rect 29273 7392 29285 7395
rect 29196 7364 29285 7392
rect 25682 7324 25688 7336
rect 22704 7296 23336 7324
rect 25148 7296 25688 7324
rect 22704 7284 22710 7296
rect 13872 7228 14596 7256
rect 13872 7216 13878 7228
rect 16114 7216 16120 7268
rect 16172 7256 16178 7268
rect 23308 7256 23336 7296
rect 25682 7284 25688 7296
rect 25740 7324 25746 7336
rect 26436 7324 26464 7352
rect 29196 7336 29224 7364
rect 29273 7361 29285 7364
rect 29319 7361 29331 7395
rect 29273 7355 29331 7361
rect 29917 7395 29975 7401
rect 29917 7361 29929 7395
rect 29963 7392 29975 7395
rect 30006 7392 30012 7404
rect 29963 7364 30012 7392
rect 29963 7361 29975 7364
rect 29917 7355 29975 7361
rect 30006 7352 30012 7364
rect 30064 7352 30070 7404
rect 30561 7395 30619 7401
rect 30561 7361 30573 7395
rect 30607 7361 30619 7395
rect 30561 7355 30619 7361
rect 25740 7296 26464 7324
rect 25740 7284 25746 7296
rect 29178 7284 29184 7336
rect 29236 7324 29242 7336
rect 30282 7324 30288 7336
rect 29236 7296 30288 7324
rect 29236 7284 29242 7296
rect 30282 7284 30288 7296
rect 30340 7324 30346 7336
rect 30576 7324 30604 7355
rect 30340 7296 30604 7324
rect 30340 7284 30346 7296
rect 24397 7259 24455 7265
rect 24397 7256 24409 7259
rect 16172 7228 18920 7256
rect 23308 7228 24409 7256
rect 16172 7216 16178 7228
rect 11054 7188 11060 7200
rect 11015 7160 11060 7188
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 11974 7148 11980 7200
rect 12032 7188 12038 7200
rect 12069 7191 12127 7197
rect 12069 7188 12081 7191
rect 12032 7160 12081 7188
rect 12032 7148 12038 7160
rect 12069 7157 12081 7160
rect 12115 7157 12127 7191
rect 12069 7151 12127 7157
rect 14182 7148 14188 7200
rect 14240 7188 14246 7200
rect 14918 7188 14924 7200
rect 14240 7160 14924 7188
rect 14240 7148 14246 7160
rect 14918 7148 14924 7160
rect 14976 7148 14982 7200
rect 16022 7148 16028 7200
rect 16080 7188 16086 7200
rect 16209 7191 16267 7197
rect 16209 7188 16221 7191
rect 16080 7160 16221 7188
rect 16080 7148 16086 7160
rect 16209 7157 16221 7160
rect 16255 7188 16267 7191
rect 18782 7188 18788 7200
rect 16255 7160 18788 7188
rect 16255 7157 16267 7160
rect 16209 7151 16267 7157
rect 18782 7148 18788 7160
rect 18840 7148 18846 7200
rect 18892 7188 18920 7228
rect 24397 7225 24409 7228
rect 24443 7225 24455 7259
rect 30466 7256 30472 7268
rect 30427 7228 30472 7256
rect 24397 7219 24455 7225
rect 30466 7216 30472 7228
rect 30524 7216 30530 7268
rect 21266 7188 21272 7200
rect 18892 7160 21272 7188
rect 21266 7148 21272 7160
rect 21324 7148 21330 7200
rect 25038 7188 25044 7200
rect 24999 7160 25044 7188
rect 25038 7148 25044 7160
rect 25096 7148 25102 7200
rect 27246 7188 27252 7200
rect 27207 7160 27252 7188
rect 27246 7148 27252 7160
rect 27304 7148 27310 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1578 6984 1584 6996
rect 1539 6956 1584 6984
rect 1578 6944 1584 6956
rect 1636 6944 1642 6996
rect 12084 6956 14044 6984
rect 9674 6808 9680 6860
rect 9732 6848 9738 6860
rect 10321 6851 10379 6857
rect 10321 6848 10333 6851
rect 9732 6820 10333 6848
rect 9732 6808 9738 6820
rect 10321 6817 10333 6820
rect 10367 6848 10379 6851
rect 12084 6848 12112 6956
rect 14016 6916 14044 6956
rect 14090 6944 14096 6996
rect 14148 6984 14154 6996
rect 15562 6984 15568 6996
rect 14148 6956 15568 6984
rect 14148 6944 14154 6956
rect 15562 6944 15568 6956
rect 15620 6944 15626 6996
rect 21082 6984 21088 6996
rect 15672 6956 21088 6984
rect 15672 6916 15700 6956
rect 21082 6944 21088 6956
rect 21140 6944 21146 6996
rect 21266 6944 21272 6996
rect 21324 6984 21330 6996
rect 27246 6984 27252 6996
rect 21324 6956 27252 6984
rect 21324 6944 21330 6956
rect 27246 6944 27252 6956
rect 27304 6944 27310 6996
rect 14016 6888 15700 6916
rect 17126 6876 17132 6928
rect 17184 6916 17190 6928
rect 17313 6919 17371 6925
rect 17313 6916 17325 6919
rect 17184 6888 17325 6916
rect 17184 6876 17190 6888
rect 17313 6885 17325 6888
rect 17359 6916 17371 6919
rect 17586 6916 17592 6928
rect 17359 6888 17592 6916
rect 17359 6885 17371 6888
rect 17313 6879 17371 6885
rect 17586 6876 17592 6888
rect 17644 6876 17650 6928
rect 17678 6876 17684 6928
rect 17736 6916 17742 6928
rect 18782 6916 18788 6928
rect 17736 6888 18788 6916
rect 17736 6876 17742 6888
rect 18782 6876 18788 6888
rect 18840 6916 18846 6928
rect 18840 6888 21312 6916
rect 18840 6876 18846 6888
rect 12253 6851 12311 6857
rect 12253 6848 12265 6851
rect 10367 6820 12265 6848
rect 10367 6817 10379 6820
rect 10321 6811 10379 6817
rect 12253 6817 12265 6820
rect 12299 6817 12311 6851
rect 12253 6811 12311 6817
rect 12894 6808 12900 6860
rect 12952 6848 12958 6860
rect 12952 6820 13492 6848
rect 12952 6808 12958 6820
rect 11974 6780 11980 6792
rect 11935 6752 11980 6780
rect 11974 6740 11980 6752
rect 12032 6740 12038 6792
rect 13464 6780 13492 6820
rect 14550 6808 14556 6860
rect 14608 6848 14614 6860
rect 15105 6851 15163 6857
rect 15105 6848 15117 6851
rect 14608 6820 15117 6848
rect 14608 6808 14614 6820
rect 15105 6817 15117 6820
rect 15151 6848 15163 6851
rect 15565 6851 15623 6857
rect 15565 6848 15577 6851
rect 15151 6820 15577 6848
rect 15151 6817 15163 6820
rect 15105 6811 15163 6817
rect 15565 6817 15577 6820
rect 15611 6848 15623 6851
rect 17770 6848 17776 6860
rect 15611 6820 17776 6848
rect 15611 6817 15623 6820
rect 15565 6811 15623 6817
rect 17770 6808 17776 6820
rect 17828 6808 17834 6860
rect 17954 6848 17960 6860
rect 17915 6820 17960 6848
rect 17954 6808 17960 6820
rect 18012 6808 18018 6860
rect 19521 6851 19579 6857
rect 19521 6848 19533 6851
rect 18800 6820 19533 6848
rect 15010 6780 15016 6792
rect 13464 6752 15016 6780
rect 15010 6740 15016 6752
rect 15068 6740 15074 6792
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 18800 6780 18828 6820
rect 19521 6817 19533 6820
rect 19567 6817 19579 6851
rect 19521 6811 19579 6817
rect 20165 6851 20223 6857
rect 20165 6817 20177 6851
rect 20211 6848 20223 6851
rect 20622 6848 20628 6860
rect 20211 6820 20628 6848
rect 20211 6817 20223 6820
rect 20165 6811 20223 6817
rect 20622 6808 20628 6820
rect 20680 6848 20686 6860
rect 20717 6851 20775 6857
rect 20717 6848 20729 6851
rect 20680 6820 20729 6848
rect 20680 6808 20686 6820
rect 20717 6817 20729 6820
rect 20763 6848 20775 6851
rect 21174 6848 21180 6860
rect 20763 6820 21180 6848
rect 20763 6817 20775 6820
rect 20717 6811 20775 6817
rect 21174 6808 21180 6820
rect 21232 6808 21238 6860
rect 21284 6848 21312 6888
rect 22462 6876 22468 6928
rect 22520 6916 22526 6928
rect 25038 6916 25044 6928
rect 22520 6888 25044 6916
rect 22520 6876 22526 6888
rect 25038 6876 25044 6888
rect 25096 6876 25102 6928
rect 25590 6876 25596 6928
rect 25648 6916 25654 6928
rect 26697 6919 26755 6925
rect 26697 6916 26709 6919
rect 25648 6888 26709 6916
rect 25648 6876 25654 6888
rect 26697 6885 26709 6888
rect 26743 6885 26755 6919
rect 26697 6879 26755 6885
rect 21453 6851 21511 6857
rect 21453 6848 21465 6851
rect 21284 6820 21465 6848
rect 21453 6817 21465 6820
rect 21499 6817 21511 6851
rect 21453 6811 21511 6817
rect 21910 6808 21916 6860
rect 21968 6848 21974 6860
rect 22925 6851 22983 6857
rect 22925 6848 22937 6851
rect 21968 6820 22937 6848
rect 21968 6808 21974 6820
rect 22925 6817 22937 6820
rect 22971 6817 22983 6851
rect 22925 6811 22983 6817
rect 24949 6851 25007 6857
rect 24949 6817 24961 6851
rect 24995 6848 25007 6851
rect 25130 6848 25136 6860
rect 24995 6820 25136 6848
rect 24995 6817 25007 6820
rect 24949 6811 25007 6817
rect 25130 6808 25136 6820
rect 25188 6808 25194 6860
rect 29089 6851 29147 6857
rect 26804 6820 28120 6848
rect 17276 6752 18828 6780
rect 17276 6740 17282 6752
rect 18874 6740 18880 6792
rect 18932 6780 18938 6792
rect 19610 6780 19616 6792
rect 18932 6752 18977 6780
rect 19571 6752 19616 6780
rect 18932 6740 18938 6752
rect 19610 6740 19616 6752
rect 19668 6740 19674 6792
rect 23198 6740 23204 6792
rect 23256 6780 23262 6792
rect 23658 6780 23664 6792
rect 23256 6752 23664 6780
rect 23256 6740 23262 6752
rect 23658 6740 23664 6752
rect 23716 6740 23722 6792
rect 24029 6783 24087 6789
rect 24029 6749 24041 6783
rect 24075 6780 24087 6783
rect 24486 6780 24492 6792
rect 24075 6752 24492 6780
rect 24075 6749 24087 6752
rect 24029 6743 24087 6749
rect 24486 6740 24492 6752
rect 24544 6740 24550 6792
rect 24762 6740 24768 6792
rect 24820 6780 24826 6792
rect 24865 6783 24923 6789
rect 24865 6780 24877 6783
rect 24820 6752 24877 6780
rect 24820 6740 24826 6752
rect 24865 6749 24877 6752
rect 24911 6749 24923 6783
rect 25590 6780 25596 6792
rect 25551 6752 25596 6780
rect 24865 6743 24923 6749
rect 25590 6740 25596 6752
rect 25648 6740 25654 6792
rect 25682 6740 25688 6792
rect 25740 6780 25746 6792
rect 26804 6789 26832 6820
rect 28092 6792 28120 6820
rect 29089 6817 29101 6851
rect 29135 6848 29147 6851
rect 29270 6848 29276 6860
rect 29135 6820 29276 6848
rect 29135 6817 29147 6820
rect 29089 6811 29147 6817
rect 29270 6808 29276 6820
rect 29328 6808 29334 6860
rect 26789 6783 26847 6789
rect 25740 6752 25785 6780
rect 25740 6740 25746 6752
rect 26789 6749 26801 6783
rect 26835 6749 26847 6783
rect 26789 6743 26847 6749
rect 26878 6740 26884 6792
rect 26936 6780 26942 6792
rect 27433 6783 27491 6789
rect 27433 6780 27445 6783
rect 26936 6752 27445 6780
rect 26936 6740 26942 6752
rect 27433 6749 27445 6752
rect 27479 6749 27491 6783
rect 28074 6780 28080 6792
rect 28035 6752 28080 6780
rect 27433 6743 27491 6749
rect 28074 6740 28080 6752
rect 28132 6740 28138 6792
rect 29178 6780 29184 6792
rect 29139 6752 29184 6780
rect 29178 6740 29184 6752
rect 29236 6740 29242 6792
rect 13478 6684 15700 6712
rect 10965 6647 11023 6653
rect 10965 6613 10977 6647
rect 11011 6644 11023 6647
rect 11054 6644 11060 6656
rect 11011 6616 11060 6644
rect 11011 6613 11023 6616
rect 10965 6607 11023 6613
rect 11054 6604 11060 6616
rect 11112 6644 11118 6656
rect 11425 6647 11483 6653
rect 11425 6644 11437 6647
rect 11112 6616 11437 6644
rect 11112 6604 11118 6616
rect 11425 6613 11437 6616
rect 11471 6613 11483 6647
rect 11425 6607 11483 6613
rect 12434 6604 12440 6656
rect 12492 6644 12498 6656
rect 13538 6644 13544 6656
rect 12492 6616 13544 6644
rect 12492 6604 12498 6616
rect 13538 6604 13544 6616
rect 13596 6644 13602 6656
rect 13725 6647 13783 6653
rect 13725 6644 13737 6647
rect 13596 6616 13737 6644
rect 13596 6604 13602 6616
rect 13725 6613 13737 6616
rect 13771 6613 13783 6647
rect 13725 6607 13783 6613
rect 14553 6647 14611 6653
rect 14553 6613 14565 6647
rect 14599 6644 14611 6647
rect 15286 6644 15292 6656
rect 14599 6616 15292 6644
rect 14599 6613 14611 6616
rect 14553 6607 14611 6613
rect 15286 6604 15292 6616
rect 15344 6604 15350 6656
rect 15672 6644 15700 6684
rect 15746 6672 15752 6724
rect 15804 6712 15810 6724
rect 15841 6715 15899 6721
rect 15841 6712 15853 6715
rect 15804 6684 15853 6712
rect 15804 6672 15810 6684
rect 15841 6681 15853 6684
rect 15887 6681 15899 6715
rect 19242 6712 19248 6724
rect 17066 6684 19248 6712
rect 15841 6675 15899 6681
rect 19242 6672 19248 6684
rect 19300 6672 19306 6724
rect 20162 6712 20168 6724
rect 19352 6684 20168 6712
rect 17218 6644 17224 6656
rect 15672 6616 17224 6644
rect 17218 6604 17224 6616
rect 17276 6604 17282 6656
rect 17586 6604 17592 6656
rect 17644 6644 17650 6656
rect 19352 6644 19380 6684
rect 20162 6672 20168 6684
rect 20220 6672 20226 6724
rect 27246 6712 27252 6724
rect 22678 6684 27252 6712
rect 27246 6672 27252 6684
rect 27304 6672 27310 6724
rect 17644 6616 19380 6644
rect 17644 6604 17650 6616
rect 19978 6604 19984 6656
rect 20036 6644 20042 6656
rect 23658 6644 23664 6656
rect 20036 6616 23664 6644
rect 20036 6604 20042 6616
rect 23658 6604 23664 6616
rect 23716 6604 23722 6656
rect 23937 6647 23995 6653
rect 23937 6613 23949 6647
rect 23983 6644 23995 6647
rect 26510 6644 26516 6656
rect 23983 6616 26516 6644
rect 23983 6613 23995 6616
rect 23937 6607 23995 6613
rect 26510 6604 26516 6616
rect 26568 6604 26574 6656
rect 27338 6644 27344 6656
rect 27299 6616 27344 6644
rect 27338 6604 27344 6616
rect 27396 6604 27402 6656
rect 27982 6644 27988 6656
rect 27943 6616 27988 6644
rect 27982 6604 27988 6616
rect 28040 6604 28046 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 12618 6400 12624 6452
rect 12676 6440 12682 6452
rect 18138 6440 18144 6452
rect 12676 6412 18144 6440
rect 12676 6400 12682 6412
rect 18138 6400 18144 6412
rect 18196 6400 18202 6452
rect 20622 6440 20628 6452
rect 18432 6412 20484 6440
rect 20583 6412 20628 6440
rect 10597 6375 10655 6381
rect 10597 6341 10609 6375
rect 10643 6372 10655 6375
rect 12894 6372 12900 6384
rect 10643 6344 12900 6372
rect 10643 6341 10655 6344
rect 10597 6335 10655 6341
rect 12894 6332 12900 6344
rect 12952 6332 12958 6384
rect 14829 6375 14887 6381
rect 14829 6341 14841 6375
rect 14875 6372 14887 6375
rect 15102 6372 15108 6384
rect 14875 6344 15108 6372
rect 14875 6341 14887 6344
rect 14829 6335 14887 6341
rect 15102 6332 15108 6344
rect 15160 6332 15166 6384
rect 18432 6372 18460 6412
rect 16054 6344 18460 6372
rect 19334 6332 19340 6384
rect 19392 6372 19398 6384
rect 20070 6372 20076 6384
rect 19392 6344 20076 6372
rect 19392 6332 19398 6344
rect 20070 6332 20076 6344
rect 20128 6332 20134 6384
rect 20456 6372 20484 6412
rect 20622 6400 20628 6412
rect 20680 6400 20686 6452
rect 27982 6440 27988 6452
rect 22066 6412 27988 6440
rect 22066 6372 22094 6412
rect 27982 6400 27988 6412
rect 28040 6400 28046 6452
rect 27893 6375 27951 6381
rect 27893 6372 27905 6375
rect 20456 6344 22094 6372
rect 23138 6344 27905 6372
rect 27893 6341 27905 6344
rect 27939 6341 27951 6375
rect 27893 6335 27951 6341
rect 29638 6332 29644 6384
rect 29696 6372 29702 6384
rect 38013 6375 38071 6381
rect 38013 6372 38025 6375
rect 29696 6344 38025 6372
rect 29696 6332 29702 6344
rect 38013 6341 38025 6344
rect 38059 6341 38071 6375
rect 38013 6335 38071 6341
rect 11698 6264 11704 6316
rect 11756 6304 11762 6316
rect 12250 6304 12256 6316
rect 11756 6276 12256 6304
rect 11756 6264 11762 6276
rect 12250 6264 12256 6276
rect 12308 6264 12314 6316
rect 13722 6264 13728 6316
rect 13780 6264 13786 6316
rect 16114 6264 16120 6316
rect 16172 6304 16178 6316
rect 17221 6307 17279 6313
rect 16172 6276 16988 6304
rect 16172 6264 16178 6276
rect 11882 6236 11888 6248
rect 11843 6208 11888 6236
rect 11882 6196 11888 6208
rect 11940 6196 11946 6248
rect 11974 6196 11980 6248
rect 12032 6236 12038 6248
rect 12345 6239 12403 6245
rect 12345 6236 12357 6239
rect 12032 6208 12357 6236
rect 12032 6196 12038 6208
rect 12345 6205 12357 6208
rect 12391 6205 12403 6239
rect 12621 6239 12679 6245
rect 12621 6236 12633 6239
rect 12345 6199 12403 6205
rect 12452 6208 12633 6236
rect 10410 6128 10416 6180
rect 10468 6168 10474 6180
rect 12452 6168 12480 6208
rect 12621 6205 12633 6208
rect 12667 6236 12679 6239
rect 14550 6236 14556 6248
rect 12667 6208 14412 6236
rect 14511 6208 14556 6236
rect 12667 6205 12679 6208
rect 12621 6199 12679 6205
rect 10468 6140 12480 6168
rect 14384 6168 14412 6208
rect 14550 6196 14556 6208
rect 14608 6196 14614 6248
rect 16301 6239 16359 6245
rect 14660 6208 15884 6236
rect 14660 6168 14688 6208
rect 14384 6140 14688 6168
rect 15856 6168 15884 6208
rect 16301 6205 16313 6239
rect 16347 6236 16359 6239
rect 16482 6236 16488 6248
rect 16347 6208 16488 6236
rect 16347 6205 16359 6208
rect 16301 6199 16359 6205
rect 16482 6196 16488 6208
rect 16540 6196 16546 6248
rect 16960 6236 16988 6276
rect 17221 6273 17233 6307
rect 17267 6304 17279 6307
rect 17770 6304 17776 6316
rect 17267 6276 17776 6304
rect 17267 6273 17279 6276
rect 17221 6267 17279 6273
rect 17770 6264 17776 6276
rect 17828 6264 17834 6316
rect 19150 6264 19156 6316
rect 19208 6264 19214 6316
rect 22278 6304 22284 6316
rect 19260 6276 22284 6304
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 16960 6208 18061 6236
rect 18049 6205 18061 6208
rect 18095 6236 18107 6239
rect 18598 6236 18604 6248
rect 18095 6208 18604 6236
rect 18095 6205 18107 6208
rect 18049 6199 18107 6205
rect 18598 6196 18604 6208
rect 18656 6196 18662 6248
rect 19260 6236 19288 6276
rect 22278 6264 22284 6276
rect 22336 6264 22342 6316
rect 24949 6307 25007 6313
rect 24949 6273 24961 6307
rect 24995 6273 25007 6307
rect 24949 6267 25007 6273
rect 19076 6208 19288 6236
rect 16666 6168 16672 6180
rect 15856 6140 16672 6168
rect 10468 6128 10474 6140
rect 16666 6128 16672 6140
rect 16724 6128 16730 6180
rect 9858 6060 9864 6112
rect 9916 6100 9922 6112
rect 9953 6103 10011 6109
rect 9953 6100 9965 6103
rect 9916 6072 9965 6100
rect 9916 6060 9922 6072
rect 9953 6069 9965 6072
rect 9999 6100 10011 6103
rect 11054 6100 11060 6112
rect 9999 6072 11060 6100
rect 9999 6069 10011 6072
rect 9953 6063 10011 6069
rect 11054 6060 11060 6072
rect 11112 6060 11118 6112
rect 12250 6060 12256 6112
rect 12308 6100 12314 6112
rect 14093 6103 14151 6109
rect 14093 6100 14105 6103
rect 12308 6072 14105 6100
rect 12308 6060 12314 6072
rect 14093 6069 14105 6072
rect 14139 6100 14151 6103
rect 15194 6100 15200 6112
rect 14139 6072 15200 6100
rect 14139 6069 14151 6072
rect 14093 6063 14151 6069
rect 15194 6060 15200 6072
rect 15252 6060 15258 6112
rect 15286 6060 15292 6112
rect 15344 6100 15350 6112
rect 17126 6100 17132 6112
rect 15344 6072 17132 6100
rect 15344 6060 15350 6072
rect 17126 6060 17132 6072
rect 17184 6060 17190 6112
rect 17218 6060 17224 6112
rect 17276 6100 17282 6112
rect 19076 6100 19104 6208
rect 19426 6196 19432 6248
rect 19484 6236 19490 6248
rect 19521 6239 19579 6245
rect 19521 6236 19533 6239
rect 19484 6208 19533 6236
rect 19484 6196 19490 6208
rect 19521 6205 19533 6208
rect 19567 6205 19579 6239
rect 19521 6199 19579 6205
rect 21726 6196 21732 6248
rect 21784 6236 21790 6248
rect 22097 6239 22155 6245
rect 22097 6236 22109 6239
rect 21784 6208 22109 6236
rect 21784 6196 21790 6208
rect 22097 6205 22109 6208
rect 22143 6205 22155 6239
rect 22097 6199 22155 6205
rect 23566 6196 23572 6248
rect 23624 6236 23630 6248
rect 23842 6236 23848 6248
rect 23624 6208 23669 6236
rect 23803 6208 23848 6236
rect 23624 6196 23630 6208
rect 23842 6196 23848 6208
rect 23900 6196 23906 6248
rect 24964 6236 24992 6267
rect 25222 6264 25228 6316
rect 25280 6304 25286 6316
rect 26145 6307 26203 6313
rect 26145 6304 26157 6307
rect 25280 6276 26157 6304
rect 25280 6264 25286 6276
rect 26145 6273 26157 6276
rect 26191 6273 26203 6307
rect 26145 6267 26203 6273
rect 26237 6307 26295 6313
rect 26237 6273 26249 6307
rect 26283 6273 26295 6307
rect 27246 6304 27252 6316
rect 27207 6276 27252 6304
rect 26237 6267 26295 6273
rect 25682 6236 25688 6248
rect 24964 6208 25688 6236
rect 25682 6196 25688 6208
rect 25740 6196 25746 6248
rect 26252 6236 26280 6267
rect 27246 6264 27252 6276
rect 27304 6264 27310 6316
rect 27341 6307 27399 6313
rect 27341 6273 27353 6307
rect 27387 6304 27399 6307
rect 27798 6304 27804 6316
rect 27387 6276 27804 6304
rect 27387 6273 27399 6276
rect 27341 6267 27399 6273
rect 27798 6264 27804 6276
rect 27856 6264 27862 6316
rect 27985 6307 28043 6313
rect 27985 6273 27997 6307
rect 28031 6304 28043 6307
rect 28166 6304 28172 6316
rect 28031 6276 28172 6304
rect 28031 6273 28043 6276
rect 27985 6267 28043 6273
rect 28166 6264 28172 6276
rect 28224 6264 28230 6316
rect 37553 6307 37611 6313
rect 37553 6273 37565 6307
rect 37599 6304 37611 6307
rect 38194 6304 38200 6316
rect 37599 6276 38200 6304
rect 37599 6273 37611 6276
rect 37553 6267 37611 6273
rect 38194 6264 38200 6276
rect 38252 6264 38258 6316
rect 33134 6236 33140 6248
rect 26252 6208 33140 6236
rect 33134 6196 33140 6208
rect 33192 6196 33198 6248
rect 19242 6128 19248 6180
rect 19300 6168 19306 6180
rect 22554 6168 22560 6180
rect 19300 6140 22560 6168
rect 19300 6128 19306 6140
rect 22554 6128 22560 6140
rect 22612 6128 22618 6180
rect 24762 6128 24768 6180
rect 24820 6168 24826 6180
rect 27338 6168 27344 6180
rect 24820 6140 27344 6168
rect 24820 6128 24826 6140
rect 27338 6128 27344 6140
rect 27396 6128 27402 6180
rect 27890 6128 27896 6180
rect 27948 6168 27954 6180
rect 28537 6171 28595 6177
rect 28537 6168 28549 6171
rect 27948 6140 28549 6168
rect 27948 6128 27954 6140
rect 28537 6137 28549 6140
rect 28583 6168 28595 6171
rect 29089 6171 29147 6177
rect 29089 6168 29101 6171
rect 28583 6140 29101 6168
rect 28583 6137 28595 6140
rect 28537 6131 28595 6137
rect 29089 6137 29101 6140
rect 29135 6168 29147 6171
rect 29641 6171 29699 6177
rect 29641 6168 29653 6171
rect 29135 6140 29653 6168
rect 29135 6137 29147 6140
rect 29089 6131 29147 6137
rect 29641 6137 29653 6140
rect 29687 6168 29699 6171
rect 30374 6168 30380 6180
rect 29687 6140 30380 6168
rect 29687 6137 29699 6140
rect 29641 6131 29699 6137
rect 30374 6128 30380 6140
rect 30432 6128 30438 6180
rect 17276 6072 19104 6100
rect 17276 6060 17282 6072
rect 20898 6060 20904 6112
rect 20956 6100 20962 6112
rect 21085 6103 21143 6109
rect 21085 6100 21097 6103
rect 20956 6072 21097 6100
rect 20956 6060 20962 6072
rect 21085 6069 21097 6072
rect 21131 6069 21143 6103
rect 21085 6063 21143 6069
rect 24857 6103 24915 6109
rect 24857 6069 24869 6103
rect 24903 6100 24915 6103
rect 24946 6100 24952 6112
rect 24903 6072 24952 6100
rect 24903 6069 24915 6072
rect 24857 6063 24915 6069
rect 24946 6060 24952 6072
rect 25004 6060 25010 6112
rect 25406 6100 25412 6112
rect 25367 6072 25412 6100
rect 25406 6060 25412 6072
rect 25464 6060 25470 6112
rect 27430 6060 27436 6112
rect 27488 6100 27494 6112
rect 30101 6103 30159 6109
rect 30101 6100 30113 6103
rect 27488 6072 30113 6100
rect 27488 6060 27494 6072
rect 30101 6069 30113 6072
rect 30147 6069 30159 6103
rect 30101 6063 30159 6069
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 10410 5896 10416 5908
rect 10371 5868 10416 5896
rect 10410 5856 10416 5868
rect 10468 5856 10474 5908
rect 13722 5856 13728 5908
rect 13780 5896 13786 5908
rect 20254 5896 20260 5908
rect 13780 5868 20260 5896
rect 13780 5856 13786 5868
rect 20254 5856 20260 5868
rect 20312 5856 20318 5908
rect 20349 5899 20407 5905
rect 20349 5865 20361 5899
rect 20395 5896 20407 5899
rect 20622 5896 20628 5908
rect 20395 5868 20628 5896
rect 20395 5865 20407 5868
rect 20349 5859 20407 5865
rect 20622 5856 20628 5868
rect 20680 5896 20686 5908
rect 20993 5899 21051 5905
rect 20993 5896 21005 5899
rect 20680 5868 21005 5896
rect 20680 5856 20686 5868
rect 20993 5865 21005 5868
rect 21039 5865 21051 5899
rect 20993 5859 21051 5865
rect 9950 5788 9956 5840
rect 10008 5828 10014 5840
rect 10318 5828 10324 5840
rect 10008 5800 10324 5828
rect 10008 5788 10014 5800
rect 10318 5788 10324 5800
rect 10376 5828 10382 5840
rect 12250 5828 12256 5840
rect 10376 5800 12256 5828
rect 10376 5788 10382 5800
rect 12250 5788 12256 5800
rect 12308 5788 12314 5840
rect 16666 5828 16672 5840
rect 16627 5800 16672 5828
rect 16666 5788 16672 5800
rect 16724 5788 16730 5840
rect 18414 5788 18420 5840
rect 18472 5828 18478 5840
rect 19705 5831 19763 5837
rect 19705 5828 19717 5831
rect 18472 5800 19717 5828
rect 18472 5788 18478 5800
rect 19705 5797 19717 5800
rect 19751 5797 19763 5831
rect 19705 5791 19763 5797
rect 11974 5720 11980 5772
rect 12032 5760 12038 5772
rect 13725 5763 13783 5769
rect 13725 5760 13737 5763
rect 12032 5732 13737 5760
rect 12032 5720 12038 5732
rect 13725 5729 13737 5732
rect 13771 5760 13783 5763
rect 14461 5763 14519 5769
rect 14461 5760 14473 5763
rect 13771 5732 14473 5760
rect 13771 5729 13783 5732
rect 13725 5723 13783 5729
rect 14461 5729 14473 5732
rect 14507 5760 14519 5763
rect 14550 5760 14556 5772
rect 14507 5732 14556 5760
rect 14507 5729 14519 5732
rect 14461 5723 14519 5729
rect 14550 5720 14556 5732
rect 14608 5760 14614 5772
rect 14921 5763 14979 5769
rect 14921 5760 14933 5763
rect 14608 5732 14933 5760
rect 14608 5720 14614 5732
rect 14921 5729 14933 5732
rect 14967 5729 14979 5763
rect 15194 5760 15200 5772
rect 15155 5732 15200 5760
rect 14921 5723 14979 5729
rect 15194 5720 15200 5732
rect 15252 5720 15258 5772
rect 17129 5763 17187 5769
rect 17129 5729 17141 5763
rect 17175 5760 17187 5763
rect 17770 5760 17776 5772
rect 17175 5732 17776 5760
rect 17175 5729 17187 5732
rect 17129 5723 17187 5729
rect 17770 5720 17776 5732
rect 17828 5720 17834 5772
rect 18138 5720 18144 5772
rect 18196 5760 18202 5772
rect 18877 5763 18935 5769
rect 18877 5760 18889 5763
rect 18196 5732 18889 5760
rect 18196 5720 18202 5732
rect 18877 5729 18889 5732
rect 18923 5760 18935 5763
rect 19426 5760 19432 5772
rect 18923 5732 19432 5760
rect 18923 5729 18935 5732
rect 18877 5723 18935 5729
rect 19426 5720 19432 5732
rect 19484 5720 19490 5772
rect 19720 5760 19748 5791
rect 20898 5760 20904 5772
rect 19720 5732 20904 5760
rect 20898 5720 20904 5732
rect 20956 5720 20962 5772
rect 21008 5760 21036 5859
rect 23106 5856 23112 5908
rect 23164 5896 23170 5908
rect 23293 5899 23351 5905
rect 23293 5896 23305 5899
rect 23164 5868 23305 5896
rect 23164 5856 23170 5868
rect 23293 5865 23305 5868
rect 23339 5865 23351 5899
rect 23293 5859 23351 5865
rect 25866 5856 25872 5908
rect 25924 5896 25930 5908
rect 27522 5896 27528 5908
rect 25924 5868 27528 5896
rect 25924 5856 25930 5868
rect 27522 5856 27528 5868
rect 27580 5856 27586 5908
rect 27890 5896 27896 5908
rect 27851 5868 27896 5896
rect 27890 5856 27896 5868
rect 27948 5856 27954 5908
rect 23382 5788 23388 5840
rect 23440 5828 23446 5840
rect 29086 5828 29092 5840
rect 23440 5800 29092 5828
rect 23440 5788 23446 5800
rect 29086 5788 29092 5800
rect 29144 5788 29150 5840
rect 21545 5763 21603 5769
rect 21545 5760 21557 5763
rect 21008 5732 21557 5760
rect 21545 5729 21557 5732
rect 21591 5729 21603 5763
rect 26694 5760 26700 5772
rect 26655 5732 26700 5760
rect 21545 5723 21603 5729
rect 26694 5720 26700 5732
rect 26752 5720 26758 5772
rect 12342 5652 12348 5704
rect 12400 5652 12406 5704
rect 21266 5692 21272 5704
rect 18538 5664 21272 5692
rect 21266 5652 21272 5664
rect 21324 5652 21330 5704
rect 24578 5692 24584 5704
rect 24539 5664 24584 5692
rect 24578 5652 24584 5664
rect 24636 5652 24642 5704
rect 24670 5652 24676 5704
rect 24728 5692 24734 5704
rect 25866 5692 25872 5704
rect 24728 5664 24773 5692
rect 25827 5664 25872 5692
rect 24728 5652 24734 5664
rect 25866 5652 25872 5664
rect 25924 5652 25930 5704
rect 26789 5695 26847 5701
rect 26789 5661 26801 5695
rect 26835 5694 26847 5695
rect 26835 5692 26924 5694
rect 28166 5692 28172 5704
rect 26835 5666 28172 5692
rect 26835 5661 26847 5666
rect 26896 5664 28172 5666
rect 26789 5655 26847 5661
rect 28166 5652 28172 5664
rect 28224 5652 28230 5704
rect 28905 5695 28963 5701
rect 28905 5661 28917 5695
rect 28951 5692 28963 5695
rect 29178 5692 29184 5704
rect 28951 5664 29184 5692
rect 28951 5661 28963 5664
rect 28905 5655 28963 5661
rect 29178 5652 29184 5664
rect 29236 5652 29242 5704
rect 11425 5627 11483 5633
rect 11425 5593 11437 5627
rect 11471 5593 11483 5627
rect 11425 5587 11483 5593
rect 13449 5627 13507 5633
rect 13449 5593 13461 5627
rect 13495 5624 13507 5627
rect 13722 5624 13728 5636
rect 13495 5596 13728 5624
rect 13495 5593 13507 5596
rect 13449 5587 13507 5593
rect 9858 5556 9864 5568
rect 9819 5528 9864 5556
rect 9858 5516 9864 5528
rect 9916 5556 9922 5568
rect 10965 5559 11023 5565
rect 10965 5556 10977 5559
rect 9916 5528 10977 5556
rect 9916 5516 9922 5528
rect 10965 5525 10977 5528
rect 11011 5556 11023 5559
rect 11440 5556 11468 5587
rect 13722 5584 13728 5596
rect 13780 5584 13786 5636
rect 16422 5596 17356 5624
rect 11011 5528 11468 5556
rect 11011 5525 11023 5528
rect 10965 5519 11023 5525
rect 11514 5516 11520 5568
rect 11572 5556 11578 5568
rect 11977 5559 12035 5565
rect 11977 5556 11989 5559
rect 11572 5528 11989 5556
rect 11572 5516 11578 5528
rect 11977 5525 11989 5528
rect 12023 5525 12035 5559
rect 17328 5556 17356 5596
rect 17402 5584 17408 5636
rect 17460 5624 17466 5636
rect 19978 5624 19984 5636
rect 17460 5596 17505 5624
rect 18708 5596 19984 5624
rect 17460 5584 17466 5596
rect 18708 5556 18736 5596
rect 19978 5584 19984 5596
rect 20036 5584 20042 5636
rect 21821 5627 21879 5633
rect 21821 5593 21833 5627
rect 21867 5624 21879 5627
rect 23382 5624 23388 5636
rect 21867 5596 22094 5624
rect 23046 5596 23388 5624
rect 21867 5593 21879 5596
rect 21821 5587 21879 5593
rect 17328 5528 18736 5556
rect 11977 5519 12035 5525
rect 20346 5516 20352 5568
rect 20404 5556 20410 5568
rect 20530 5556 20536 5568
rect 20404 5528 20536 5556
rect 20404 5516 20410 5528
rect 20530 5516 20536 5528
rect 20588 5516 20594 5568
rect 22066 5556 22094 5596
rect 23382 5584 23388 5596
rect 23440 5584 23446 5636
rect 23658 5584 23664 5636
rect 23716 5624 23722 5636
rect 23716 5596 24348 5624
rect 23716 5584 23722 5596
rect 23198 5556 23204 5568
rect 22066 5528 23204 5556
rect 23198 5516 23204 5528
rect 23256 5516 23262 5568
rect 23845 5559 23903 5565
rect 23845 5525 23857 5559
rect 23891 5556 23903 5559
rect 24026 5556 24032 5568
rect 23891 5528 24032 5556
rect 23891 5525 23903 5528
rect 23845 5519 23903 5525
rect 24026 5516 24032 5528
rect 24084 5516 24090 5568
rect 24320 5556 24348 5596
rect 25406 5584 25412 5636
rect 25464 5624 25470 5636
rect 28813 5627 28871 5633
rect 28813 5624 28825 5627
rect 25464 5596 28825 5624
rect 25464 5584 25470 5596
rect 28813 5593 28825 5596
rect 28859 5593 28871 5627
rect 28813 5587 28871 5593
rect 25498 5556 25504 5568
rect 24320 5528 25504 5556
rect 25498 5516 25504 5528
rect 25556 5516 25562 5568
rect 25774 5556 25780 5568
rect 25735 5528 25780 5556
rect 25774 5516 25780 5528
rect 25832 5516 25838 5568
rect 25958 5516 25964 5568
rect 26016 5556 26022 5568
rect 27249 5559 27307 5565
rect 27249 5556 27261 5559
rect 26016 5528 27261 5556
rect 26016 5516 26022 5528
rect 27249 5525 27261 5528
rect 27295 5525 27307 5559
rect 27249 5519 27307 5525
rect 29825 5559 29883 5565
rect 29825 5525 29837 5559
rect 29871 5556 29883 5559
rect 30374 5556 30380 5568
rect 29871 5528 30380 5556
rect 29871 5525 29883 5528
rect 29825 5519 29883 5525
rect 30374 5516 30380 5528
rect 30432 5516 30438 5568
rect 30834 5556 30840 5568
rect 30795 5528 30840 5556
rect 30834 5516 30840 5528
rect 30892 5516 30898 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 8754 5312 8760 5364
rect 8812 5352 8818 5364
rect 14093 5355 14151 5361
rect 8812 5324 14044 5352
rect 8812 5312 8818 5324
rect 11514 5244 11520 5296
rect 11572 5284 11578 5296
rect 12621 5287 12679 5293
rect 12621 5284 12633 5287
rect 11572 5256 12633 5284
rect 11572 5244 11578 5256
rect 12621 5253 12633 5256
rect 12667 5253 12679 5287
rect 14016 5284 14044 5324
rect 14093 5321 14105 5355
rect 14139 5352 14151 5355
rect 14734 5352 14740 5364
rect 14139 5324 14740 5352
rect 14139 5321 14151 5324
rect 14093 5315 14151 5321
rect 14734 5312 14740 5324
rect 14792 5312 14798 5364
rect 14918 5312 14924 5364
rect 14976 5352 14982 5364
rect 20162 5352 20168 5364
rect 14976 5324 20168 5352
rect 14976 5312 14982 5324
rect 20162 5312 20168 5324
rect 20220 5312 20226 5364
rect 25774 5352 25780 5364
rect 20272 5324 25780 5352
rect 14458 5284 14464 5296
rect 14016 5256 14464 5284
rect 12621 5247 12679 5253
rect 14458 5244 14464 5256
rect 14516 5244 14522 5296
rect 14826 5244 14832 5296
rect 14884 5284 14890 5296
rect 16482 5284 16488 5296
rect 14884 5256 14929 5284
rect 16054 5256 16488 5284
rect 14884 5244 14890 5256
rect 16482 5244 16488 5256
rect 16540 5244 16546 5296
rect 17770 5284 17776 5296
rect 17420 5256 17776 5284
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5216 1915 5219
rect 2774 5216 2780 5228
rect 1903 5188 2780 5216
rect 1903 5185 1915 5188
rect 1857 5179 1915 5185
rect 2774 5176 2780 5188
rect 2832 5176 2838 5228
rect 11974 5176 11980 5228
rect 12032 5216 12038 5228
rect 12345 5219 12403 5225
rect 12345 5216 12357 5219
rect 12032 5188 12357 5216
rect 12032 5176 12038 5188
rect 12345 5185 12357 5188
rect 12391 5185 12403 5219
rect 12345 5179 12403 5185
rect 13722 5176 13728 5228
rect 13780 5176 13786 5228
rect 14550 5216 14556 5228
rect 14511 5188 14556 5216
rect 14550 5176 14556 5188
rect 14608 5176 14614 5228
rect 16945 5219 17003 5225
rect 16945 5185 16957 5219
rect 16991 5216 17003 5219
rect 17126 5216 17132 5228
rect 16991 5188 17132 5216
rect 16991 5185 17003 5188
rect 16945 5179 17003 5185
rect 17126 5176 17132 5188
rect 17184 5216 17190 5228
rect 17420 5225 17448 5256
rect 17770 5244 17776 5256
rect 17828 5244 17834 5296
rect 20272 5284 20300 5324
rect 25774 5312 25780 5324
rect 25832 5312 25838 5364
rect 27246 5352 27252 5364
rect 27207 5324 27252 5352
rect 27246 5312 27252 5324
rect 27304 5312 27310 5364
rect 28534 5312 28540 5364
rect 28592 5352 28598 5364
rect 31205 5355 31263 5361
rect 31205 5352 31217 5355
rect 28592 5324 31217 5352
rect 28592 5312 28598 5324
rect 31205 5321 31217 5324
rect 31251 5321 31263 5355
rect 31205 5315 31263 5321
rect 22370 5284 22376 5296
rect 18906 5256 20300 5284
rect 21114 5256 22376 5284
rect 22370 5244 22376 5256
rect 22428 5244 22434 5296
rect 24762 5284 24768 5296
rect 23506 5256 24768 5284
rect 24762 5244 24768 5256
rect 24820 5244 24826 5296
rect 30101 5287 30159 5293
rect 30101 5284 30113 5287
rect 24872 5256 30113 5284
rect 17405 5219 17463 5225
rect 17405 5216 17417 5219
rect 17184 5188 17417 5216
rect 17184 5176 17190 5188
rect 17405 5185 17417 5188
rect 17451 5185 17463 5219
rect 17405 5179 17463 5185
rect 24394 5176 24400 5228
rect 24452 5216 24458 5228
rect 24872 5216 24900 5256
rect 30101 5253 30113 5256
rect 30147 5253 30159 5287
rect 30101 5247 30159 5253
rect 24452 5188 24900 5216
rect 24452 5176 24458 5188
rect 25038 5176 25044 5228
rect 25096 5216 25102 5228
rect 26513 5219 26571 5225
rect 25096 5188 25544 5216
rect 25096 5176 25102 5188
rect 9493 5151 9551 5157
rect 9493 5117 9505 5151
rect 9539 5148 9551 5151
rect 13814 5148 13820 5160
rect 9539 5120 13820 5148
rect 9539 5117 9551 5120
rect 9493 5111 9551 5117
rect 13814 5108 13820 5120
rect 13872 5148 13878 5160
rect 16298 5148 16304 5160
rect 13872 5120 16304 5148
rect 13872 5108 13878 5120
rect 16298 5108 16304 5120
rect 16356 5108 16362 5160
rect 17034 5108 17040 5160
rect 17092 5148 17098 5160
rect 17681 5151 17739 5157
rect 17681 5148 17693 5151
rect 17092 5120 17693 5148
rect 17092 5108 17098 5120
rect 17681 5117 17693 5120
rect 17727 5117 17739 5151
rect 17681 5111 17739 5117
rect 18046 5108 18052 5160
rect 18104 5148 18110 5160
rect 19610 5148 19616 5160
rect 18104 5120 18736 5148
rect 19571 5120 19616 5148
rect 18104 5108 18110 5120
rect 14550 5080 14556 5092
rect 13648 5052 14556 5080
rect 1670 5012 1676 5024
rect 1631 4984 1676 5012
rect 1670 4972 1676 4984
rect 1728 4972 1734 5024
rect 9306 4972 9312 5024
rect 9364 5012 9370 5024
rect 9858 5012 9864 5024
rect 9364 4984 9864 5012
rect 9364 4972 9370 4984
rect 9858 4972 9864 4984
rect 9916 5012 9922 5024
rect 9953 5015 10011 5021
rect 9953 5012 9965 5015
rect 9916 4984 9965 5012
rect 9916 4972 9922 4984
rect 9953 4981 9965 4984
rect 9999 5012 10011 5015
rect 10505 5015 10563 5021
rect 10505 5012 10517 5015
rect 9999 4984 10517 5012
rect 9999 4981 10011 4984
rect 9953 4975 10011 4981
rect 10505 4981 10517 4984
rect 10551 5012 10563 5015
rect 11054 5012 11060 5024
rect 10551 4984 11060 5012
rect 10551 4981 10563 4984
rect 10505 4975 10563 4981
rect 11054 4972 11060 4984
rect 11112 4972 11118 5024
rect 11885 5015 11943 5021
rect 11885 4981 11897 5015
rect 11931 5012 11943 5015
rect 13648 5012 13676 5052
rect 14550 5040 14556 5052
rect 14608 5040 14614 5092
rect 18708 5080 18736 5120
rect 19610 5108 19616 5120
rect 19668 5108 19674 5160
rect 19889 5151 19947 5157
rect 19889 5148 19901 5151
rect 19720 5120 19901 5148
rect 19058 5080 19064 5092
rect 15856 5052 16436 5080
rect 18708 5052 19064 5080
rect 11931 4984 13676 5012
rect 11931 4981 11943 4984
rect 11885 4975 11943 4981
rect 13722 4972 13728 5024
rect 13780 5012 13786 5024
rect 15856 5012 15884 5052
rect 13780 4984 15884 5012
rect 13780 4972 13786 4984
rect 16114 4972 16120 5024
rect 16172 5012 16178 5024
rect 16301 5015 16359 5021
rect 16301 5012 16313 5015
rect 16172 4984 16313 5012
rect 16172 4972 16178 4984
rect 16301 4981 16313 4984
rect 16347 4981 16359 5015
rect 16408 5012 16436 5052
rect 19058 5040 19064 5052
rect 19116 5080 19122 5092
rect 19720 5080 19748 5120
rect 19889 5117 19901 5120
rect 19935 5117 19947 5151
rect 19889 5111 19947 5117
rect 20622 5108 20628 5160
rect 20680 5148 20686 5160
rect 21818 5148 21824 5160
rect 20680 5120 21824 5148
rect 20680 5108 20686 5120
rect 21818 5108 21824 5120
rect 21876 5148 21882 5160
rect 22005 5151 22063 5157
rect 22005 5148 22017 5151
rect 21876 5120 22017 5148
rect 21876 5108 21882 5120
rect 22005 5117 22017 5120
rect 22051 5117 22063 5151
rect 22278 5148 22284 5160
rect 22239 5120 22284 5148
rect 22005 5111 22063 5117
rect 22278 5108 22284 5120
rect 22336 5108 22342 5160
rect 22370 5108 22376 5160
rect 22428 5148 22434 5160
rect 25406 5148 25412 5160
rect 22428 5120 25412 5148
rect 22428 5108 22434 5120
rect 25406 5108 25412 5120
rect 25464 5108 25470 5160
rect 25516 5148 25544 5188
rect 26513 5185 26525 5219
rect 26559 5216 26571 5219
rect 26878 5216 26884 5228
rect 26559 5188 26884 5216
rect 26559 5185 26571 5188
rect 26513 5179 26571 5185
rect 26878 5176 26884 5188
rect 26936 5176 26942 5228
rect 27341 5219 27399 5225
rect 27341 5185 27353 5219
rect 27387 5216 27399 5219
rect 27522 5216 27528 5228
rect 27387 5188 27528 5216
rect 27387 5185 27399 5188
rect 27341 5179 27399 5185
rect 27522 5176 27528 5188
rect 27580 5176 27586 5228
rect 27982 5216 27988 5228
rect 27943 5188 27988 5216
rect 27982 5176 27988 5188
rect 28040 5176 28046 5228
rect 28074 5176 28080 5228
rect 28132 5216 28138 5228
rect 28905 5219 28963 5225
rect 28905 5216 28917 5219
rect 28132 5188 28917 5216
rect 28132 5176 28138 5188
rect 28905 5185 28917 5188
rect 28951 5216 28963 5219
rect 29549 5219 29607 5225
rect 29549 5216 29561 5219
rect 28951 5188 29561 5216
rect 28951 5185 28963 5188
rect 28905 5179 28963 5185
rect 29549 5185 29561 5188
rect 29595 5216 29607 5219
rect 29914 5216 29920 5228
rect 29595 5188 29920 5216
rect 29595 5185 29607 5188
rect 29549 5179 29607 5185
rect 29914 5176 29920 5188
rect 29972 5176 29978 5228
rect 30006 5176 30012 5228
rect 30064 5216 30070 5228
rect 30193 5219 30251 5225
rect 30193 5216 30205 5219
rect 30064 5188 30205 5216
rect 30064 5176 30070 5188
rect 30193 5185 30205 5188
rect 30239 5185 30251 5219
rect 30193 5179 30251 5185
rect 29457 5151 29515 5157
rect 29457 5148 29469 5151
rect 25516 5120 29469 5148
rect 29457 5117 29469 5120
rect 29503 5117 29515 5151
rect 38010 5148 38016 5160
rect 37971 5120 38016 5148
rect 29457 5111 29515 5117
rect 38010 5108 38016 5120
rect 38068 5108 38074 5160
rect 38286 5148 38292 5160
rect 38247 5120 38292 5148
rect 38286 5108 38292 5120
rect 38344 5108 38350 5160
rect 21910 5080 21916 5092
rect 19116 5052 19748 5080
rect 21192 5052 21916 5080
rect 19116 5040 19122 5052
rect 19153 5015 19211 5021
rect 19153 5012 19165 5015
rect 16408 4984 19165 5012
rect 16301 4975 16359 4981
rect 19153 4981 19165 4984
rect 19199 4981 19211 5015
rect 19153 4975 19211 4981
rect 19242 4972 19248 5024
rect 19300 5012 19306 5024
rect 21192 5012 21220 5052
rect 21910 5040 21916 5052
rect 21968 5040 21974 5092
rect 23566 5040 23572 5092
rect 23624 5080 23630 5092
rect 27893 5083 27951 5089
rect 27893 5080 27905 5083
rect 23624 5052 27905 5080
rect 23624 5040 23630 5052
rect 27893 5049 27905 5052
rect 27939 5049 27951 5083
rect 27893 5043 27951 5049
rect 30374 5040 30380 5092
rect 30432 5080 30438 5092
rect 30745 5083 30803 5089
rect 30745 5080 30757 5083
rect 30432 5052 30757 5080
rect 30432 5040 30438 5052
rect 30745 5049 30757 5052
rect 30791 5080 30803 5083
rect 33594 5080 33600 5092
rect 30791 5052 33600 5080
rect 30791 5049 30803 5052
rect 30745 5043 30803 5049
rect 33594 5040 33600 5052
rect 33652 5040 33658 5092
rect 21358 5012 21364 5024
rect 19300 4984 21220 5012
rect 21319 4984 21364 5012
rect 19300 4972 19306 4984
rect 21358 4972 21364 4984
rect 21416 4972 21422 5024
rect 21450 4972 21456 5024
rect 21508 5012 21514 5024
rect 23474 5012 23480 5024
rect 21508 4984 23480 5012
rect 21508 4972 21514 4984
rect 23474 4972 23480 4984
rect 23532 4972 23538 5024
rect 23750 5012 23756 5024
rect 23711 4984 23756 5012
rect 23750 4972 23756 4984
rect 23808 4972 23814 5024
rect 24305 5015 24363 5021
rect 24305 4981 24317 5015
rect 24351 5012 24363 5015
rect 24762 5012 24768 5024
rect 24351 4984 24768 5012
rect 24351 4981 24363 4984
rect 24305 4975 24363 4981
rect 24762 4972 24768 4984
rect 24820 5012 24826 5024
rect 25317 5015 25375 5021
rect 25317 5012 25329 5015
rect 24820 4984 25329 5012
rect 24820 4972 24826 4984
rect 25317 4981 25329 4984
rect 25363 4981 25375 5015
rect 26418 5012 26424 5024
rect 26379 4984 26424 5012
rect 25317 4975 25375 4981
rect 26418 4972 26424 4984
rect 26476 4972 26482 5024
rect 28810 5012 28816 5024
rect 28771 4984 28816 5012
rect 28810 4972 28816 4984
rect 28868 4972 28874 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 11054 4768 11060 4820
rect 11112 4808 11118 4820
rect 11425 4811 11483 4817
rect 11425 4808 11437 4811
rect 11112 4780 11437 4808
rect 11112 4768 11118 4780
rect 11425 4777 11437 4780
rect 11471 4777 11483 4811
rect 11425 4771 11483 4777
rect 11532 4780 18644 4808
rect 10502 4700 10508 4752
rect 10560 4740 10566 4752
rect 11532 4740 11560 4780
rect 14918 4740 14924 4752
rect 10560 4712 11560 4740
rect 13648 4712 14924 4740
rect 10560 4700 10566 4712
rect 11054 4632 11060 4684
rect 11112 4672 11118 4684
rect 11974 4672 11980 4684
rect 11112 4644 11980 4672
rect 11112 4632 11118 4644
rect 11974 4632 11980 4644
rect 12032 4632 12038 4684
rect 12253 4675 12311 4681
rect 12253 4641 12265 4675
rect 12299 4672 12311 4675
rect 13648 4672 13676 4712
rect 14918 4700 14924 4712
rect 14976 4700 14982 4752
rect 16850 4740 16856 4752
rect 16316 4712 16856 4740
rect 12299 4644 13676 4672
rect 13725 4675 13783 4681
rect 12299 4641 12311 4644
rect 12253 4635 12311 4641
rect 13725 4641 13737 4675
rect 13771 4672 13783 4675
rect 16316 4672 16344 4712
rect 16850 4700 16856 4712
rect 16908 4700 16914 4752
rect 18616 4740 18644 4780
rect 18782 4768 18788 4820
rect 18840 4808 18846 4820
rect 18877 4811 18935 4817
rect 18877 4808 18889 4811
rect 18840 4780 18889 4808
rect 18840 4768 18846 4780
rect 18877 4777 18889 4780
rect 18923 4777 18935 4811
rect 18877 4771 18935 4777
rect 19334 4768 19340 4820
rect 19392 4808 19398 4820
rect 19521 4811 19579 4817
rect 19521 4808 19533 4811
rect 19392 4780 19533 4808
rect 19392 4768 19398 4780
rect 19521 4777 19533 4780
rect 19567 4808 19579 4811
rect 19610 4808 19616 4820
rect 19567 4780 19616 4808
rect 19567 4777 19579 4780
rect 19521 4771 19579 4777
rect 19610 4768 19616 4780
rect 19668 4808 19674 4820
rect 20622 4808 20628 4820
rect 19668 4780 20628 4808
rect 19668 4768 19674 4780
rect 20622 4768 20628 4780
rect 20680 4808 20686 4820
rect 20809 4811 20867 4817
rect 20809 4808 20821 4811
rect 20680 4780 20821 4808
rect 20680 4768 20686 4780
rect 20809 4777 20821 4780
rect 20855 4777 20867 4811
rect 20809 4771 20867 4777
rect 21174 4768 21180 4820
rect 21232 4808 21238 4820
rect 23566 4808 23572 4820
rect 21232 4780 23572 4808
rect 21232 4768 21238 4780
rect 23566 4768 23572 4780
rect 23624 4768 23630 4820
rect 23661 4811 23719 4817
rect 23661 4777 23673 4811
rect 23707 4808 23719 4811
rect 23842 4808 23848 4820
rect 23707 4780 23848 4808
rect 23707 4777 23719 4780
rect 23661 4771 23719 4777
rect 18616 4712 21588 4740
rect 13771 4644 16344 4672
rect 16393 4675 16451 4681
rect 13771 4641 13783 4644
rect 13725 4635 13783 4641
rect 16393 4641 16405 4675
rect 16439 4672 16451 4675
rect 17126 4672 17132 4684
rect 16439 4644 17132 4672
rect 16439 4641 16451 4644
rect 16393 4635 16451 4641
rect 17126 4632 17132 4644
rect 17184 4632 17190 4684
rect 20070 4672 20076 4684
rect 20031 4644 20076 4672
rect 20070 4632 20076 4644
rect 20128 4632 20134 4684
rect 9861 4607 9919 4613
rect 9861 4573 9873 4607
rect 9907 4604 9919 4607
rect 13630 4604 13636 4616
rect 9907 4576 12020 4604
rect 13386 4576 13636 4604
rect 9907 4573 9919 4576
rect 9861 4567 9919 4573
rect 11992 4536 12020 4576
rect 13630 4564 13636 4576
rect 13688 4564 13694 4616
rect 21174 4604 21180 4616
rect 18538 4576 21180 4604
rect 21174 4564 21180 4576
rect 21232 4564 21238 4616
rect 12342 4536 12348 4548
rect 11992 4508 12348 4536
rect 12342 4496 12348 4508
rect 12400 4496 12406 4548
rect 14826 4536 14832 4548
rect 13924 4508 14832 4536
rect 9306 4468 9312 4480
rect 9267 4440 9312 4468
rect 9306 4428 9312 4440
rect 9364 4468 9370 4480
rect 10413 4471 10471 4477
rect 10413 4468 10425 4471
rect 9364 4440 10425 4468
rect 9364 4428 9370 4440
rect 10413 4437 10425 4440
rect 10459 4437 10471 4471
rect 10413 4431 10471 4437
rect 10965 4471 11023 4477
rect 10965 4437 10977 4471
rect 11011 4468 11023 4471
rect 13924 4468 13952 4508
rect 14826 4496 14832 4508
rect 14884 4496 14890 4548
rect 16117 4539 16175 4545
rect 15686 4508 16068 4536
rect 14642 4468 14648 4480
rect 11011 4440 13952 4468
rect 14603 4440 14648 4468
rect 11011 4437 11023 4440
rect 10965 4431 11023 4437
rect 14642 4428 14648 4440
rect 14700 4428 14706 4480
rect 16040 4468 16068 4508
rect 16117 4505 16129 4539
rect 16163 4536 16175 4539
rect 16206 4536 16212 4548
rect 16163 4508 16212 4536
rect 16163 4505 16175 4508
rect 16117 4499 16175 4505
rect 16206 4496 16212 4508
rect 16264 4496 16270 4548
rect 16666 4496 16672 4548
rect 16724 4536 16730 4548
rect 17405 4539 17463 4545
rect 17405 4536 17417 4539
rect 16724 4508 17417 4536
rect 16724 4496 16730 4508
rect 17405 4505 17417 4508
rect 17451 4505 17463 4539
rect 21450 4536 21456 4548
rect 17405 4499 17463 4505
rect 18708 4508 21456 4536
rect 18708 4468 18736 4508
rect 21450 4496 21456 4508
rect 21508 4496 21514 4548
rect 16040 4440 18736 4468
rect 21361 4471 21419 4477
rect 21361 4437 21373 4471
rect 21407 4468 21419 4471
rect 21560 4468 21588 4712
rect 21818 4632 21824 4684
rect 21876 4672 21882 4684
rect 23109 4675 23167 4681
rect 23109 4672 23121 4675
rect 21876 4644 23121 4672
rect 21876 4632 21882 4644
rect 23109 4641 23121 4644
rect 23155 4672 23167 4675
rect 23676 4672 23704 4771
rect 23842 4768 23848 4780
rect 23900 4808 23906 4820
rect 24673 4811 24731 4817
rect 24673 4808 24685 4811
rect 23900 4780 24685 4808
rect 23900 4768 23906 4780
rect 24673 4777 24685 4780
rect 24719 4808 24731 4811
rect 24762 4808 24768 4820
rect 24719 4780 24768 4808
rect 24719 4777 24731 4780
rect 24673 4771 24731 4777
rect 24762 4768 24768 4780
rect 24820 4808 24826 4820
rect 25225 4811 25283 4817
rect 25225 4808 25237 4811
rect 24820 4780 25237 4808
rect 24820 4768 24826 4780
rect 25225 4777 25237 4780
rect 25271 4808 25283 4811
rect 25777 4811 25835 4817
rect 25777 4808 25789 4811
rect 25271 4780 25789 4808
rect 25271 4777 25283 4780
rect 25225 4771 25283 4777
rect 25777 4777 25789 4780
rect 25823 4808 25835 4811
rect 26234 4808 26240 4820
rect 25823 4780 26240 4808
rect 25823 4777 25835 4780
rect 25777 4771 25835 4777
rect 26234 4768 26240 4780
rect 26292 4808 26298 4820
rect 26329 4811 26387 4817
rect 26329 4808 26341 4811
rect 26292 4780 26341 4808
rect 26292 4768 26298 4780
rect 26329 4777 26341 4780
rect 26375 4808 26387 4811
rect 27706 4808 27712 4820
rect 26375 4780 27712 4808
rect 26375 4777 26387 4780
rect 26329 4771 26387 4777
rect 27706 4768 27712 4780
rect 27764 4768 27770 4820
rect 28626 4768 28632 4820
rect 28684 4808 28690 4820
rect 29089 4811 29147 4817
rect 29089 4808 29101 4811
rect 28684 4780 29101 4808
rect 28684 4768 28690 4780
rect 29089 4777 29101 4780
rect 29135 4777 29147 4811
rect 33042 4808 33048 4820
rect 33003 4780 33048 4808
rect 29089 4771 29147 4777
rect 33042 4768 33048 4780
rect 33100 4768 33106 4820
rect 38286 4808 38292 4820
rect 38247 4780 38292 4808
rect 38286 4768 38292 4780
rect 38344 4768 38350 4820
rect 27154 4700 27160 4752
rect 27212 4740 27218 4752
rect 29825 4743 29883 4749
rect 29825 4740 29837 4743
rect 27212 4712 29837 4740
rect 27212 4700 27218 4712
rect 29825 4709 29837 4712
rect 29871 4709 29883 4743
rect 29825 4703 29883 4709
rect 31021 4675 31079 4681
rect 31021 4672 31033 4675
rect 23155 4644 23704 4672
rect 23768 4644 31033 4672
rect 23155 4641 23167 4644
rect 23109 4635 23167 4641
rect 23474 4564 23480 4616
rect 23532 4604 23538 4616
rect 23768 4604 23796 4644
rect 31021 4641 31033 4644
rect 31067 4641 31079 4675
rect 38010 4672 38016 4684
rect 31021 4635 31079 4641
rect 35866 4644 38016 4672
rect 27062 4604 27068 4616
rect 23532 4576 23796 4604
rect 27023 4576 27068 4604
rect 23532 4564 23538 4576
rect 27062 4564 27068 4576
rect 27120 4564 27126 4616
rect 27157 4607 27215 4613
rect 27157 4573 27169 4607
rect 27203 4604 27215 4607
rect 27430 4604 27436 4616
rect 27203 4576 27436 4604
rect 27203 4573 27215 4576
rect 27157 4567 27215 4573
rect 27430 4564 27436 4576
rect 27488 4604 27494 4616
rect 28166 4604 28172 4616
rect 27488 4576 28172 4604
rect 27488 4564 27494 4576
rect 28166 4564 28172 4576
rect 28224 4564 28230 4616
rect 28442 4604 28448 4616
rect 28403 4576 28448 4604
rect 28442 4564 28448 4576
rect 28500 4564 28506 4616
rect 29178 4604 29184 4616
rect 29091 4576 29184 4604
rect 29178 4564 29184 4576
rect 29236 4604 29242 4616
rect 29917 4607 29975 4613
rect 29917 4604 29929 4607
rect 29236 4576 29929 4604
rect 29236 4564 29242 4576
rect 29917 4573 29929 4576
rect 29963 4604 29975 4607
rect 30561 4607 30619 4613
rect 30561 4604 30573 4607
rect 29963 4576 30573 4604
rect 29963 4573 29975 4576
rect 29917 4567 29975 4573
rect 30561 4573 30573 4576
rect 30607 4604 30619 4607
rect 31202 4604 31208 4616
rect 30607 4576 31208 4604
rect 30607 4573 30619 4576
rect 30561 4567 30619 4573
rect 31202 4564 31208 4576
rect 31260 4604 31266 4616
rect 31846 4604 31852 4616
rect 31260 4576 31852 4604
rect 31260 4564 31266 4576
rect 31846 4564 31852 4576
rect 31904 4604 31910 4616
rect 32217 4607 32275 4613
rect 32217 4604 32229 4607
rect 31904 4576 32229 4604
rect 31904 4564 31910 4576
rect 32217 4573 32229 4576
rect 32263 4573 32275 4607
rect 32217 4567 32275 4573
rect 32493 4607 32551 4613
rect 32493 4573 32505 4607
rect 32539 4604 32551 4607
rect 33042 4604 33048 4616
rect 32539 4576 33048 4604
rect 32539 4573 32551 4576
rect 32493 4567 32551 4573
rect 33042 4564 33048 4576
rect 33100 4564 33106 4616
rect 22833 4539 22891 4545
rect 22402 4508 22784 4536
rect 22094 4468 22100 4480
rect 21407 4440 22100 4468
rect 21407 4437 21419 4440
rect 21361 4431 21419 4437
rect 22094 4428 22100 4440
rect 22152 4428 22158 4480
rect 22756 4468 22784 4508
rect 22833 4505 22845 4539
rect 22879 4536 22891 4539
rect 23106 4536 23112 4548
rect 22879 4508 23112 4536
rect 22879 4505 22891 4508
rect 22833 4499 22891 4505
rect 23106 4496 23112 4508
rect 23164 4496 23170 4548
rect 23198 4496 23204 4548
rect 23256 4536 23262 4548
rect 25590 4536 25596 4548
rect 23256 4508 25596 4536
rect 23256 4496 23262 4508
rect 25590 4496 25596 4508
rect 25648 4496 25654 4548
rect 26326 4496 26332 4548
rect 26384 4536 26390 4548
rect 30469 4539 30527 4545
rect 30469 4536 30481 4539
rect 26384 4508 30481 4536
rect 26384 4496 26390 4508
rect 30469 4505 30481 4508
rect 30515 4505 30527 4539
rect 30469 4499 30527 4505
rect 26970 4468 26976 4480
rect 22756 4440 26976 4468
rect 26970 4428 26976 4440
rect 27028 4428 27034 4480
rect 27062 4428 27068 4480
rect 27120 4468 27126 4480
rect 28261 4471 28319 4477
rect 28261 4468 28273 4471
rect 27120 4440 28273 4468
rect 27120 4428 27126 4440
rect 28261 4437 28273 4440
rect 28307 4437 28319 4471
rect 28261 4431 28319 4437
rect 28442 4428 28448 4480
rect 28500 4468 28506 4480
rect 35866 4468 35894 4644
rect 38010 4632 38016 4644
rect 38068 4632 38074 4684
rect 28500 4440 35894 4468
rect 28500 4428 28506 4440
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 10042 4264 10048 4276
rect 10003 4236 10048 4264
rect 10042 4224 10048 4236
rect 10100 4224 10106 4276
rect 11054 4264 11060 4276
rect 11015 4236 11060 4264
rect 11054 4224 11060 4236
rect 11112 4224 11118 4276
rect 12069 4267 12127 4273
rect 12069 4233 12081 4267
rect 12115 4264 12127 4267
rect 12526 4264 12532 4276
rect 12115 4236 12532 4264
rect 12115 4233 12127 4236
rect 12069 4227 12127 4233
rect 12526 4224 12532 4236
rect 12584 4224 12590 4276
rect 20530 4264 20536 4276
rect 13464 4236 20536 4264
rect 13464 4196 13492 4236
rect 20530 4224 20536 4236
rect 20588 4224 20594 4276
rect 20622 4224 20628 4276
rect 20680 4264 20686 4276
rect 21361 4267 21419 4273
rect 21361 4264 21373 4267
rect 20680 4236 21373 4264
rect 20680 4224 20686 4236
rect 21361 4233 21373 4236
rect 21407 4233 21419 4267
rect 21361 4227 21419 4233
rect 21450 4224 21456 4276
rect 21508 4264 21514 4276
rect 26418 4264 26424 4276
rect 21508 4236 26424 4264
rect 21508 4224 21514 4236
rect 26418 4224 26424 4236
rect 26476 4224 26482 4276
rect 26970 4224 26976 4276
rect 27028 4264 27034 4276
rect 30374 4264 30380 4276
rect 27028 4236 30380 4264
rect 27028 4224 27034 4236
rect 30374 4224 30380 4236
rect 30432 4224 30438 4276
rect 13110 4168 13492 4196
rect 13541 4199 13599 4205
rect 13541 4165 13553 4199
rect 13587 4196 13599 4199
rect 13814 4196 13820 4208
rect 13587 4168 13820 4196
rect 13587 4165 13599 4168
rect 13541 4159 13599 4165
rect 13814 4156 13820 4168
rect 13872 4156 13878 4208
rect 16206 4196 16212 4208
rect 15778 4168 16212 4196
rect 16206 4156 16212 4168
rect 16264 4156 16270 4208
rect 16298 4156 16304 4208
rect 16356 4196 16362 4208
rect 16356 4168 16401 4196
rect 16356 4156 16362 4168
rect 16482 4156 16488 4208
rect 16540 4196 16546 4208
rect 19150 4196 19156 4208
rect 16540 4168 19156 4196
rect 16540 4156 16546 4168
rect 19150 4156 19156 4168
rect 19208 4156 19214 4208
rect 22186 4196 22192 4208
rect 20102 4168 22192 4196
rect 22186 4156 22192 4168
rect 22244 4156 22250 4208
rect 24394 4196 24400 4208
rect 23046 4168 24400 4196
rect 24394 4156 24400 4168
rect 24452 4156 24458 4208
rect 24486 4156 24492 4208
rect 24544 4196 24550 4208
rect 28810 4196 28816 4208
rect 24544 4168 24589 4196
rect 25714 4168 28816 4196
rect 24544 4156 24550 4168
rect 28810 4156 28816 4168
rect 28868 4156 28874 4208
rect 30006 4196 30012 4208
rect 29288 4168 30012 4196
rect 16850 4128 16856 4140
rect 16811 4100 16856 4128
rect 16850 4088 16856 4100
rect 16908 4088 16914 4140
rect 21266 4128 21272 4140
rect 20088 4100 21272 4128
rect 13817 4063 13875 4069
rect 13817 4029 13829 4063
rect 13863 4060 13875 4063
rect 14277 4063 14335 4069
rect 14277 4060 14289 4063
rect 13863 4032 14289 4060
rect 13863 4029 13875 4032
rect 13817 4023 13875 4029
rect 14277 4029 14289 4032
rect 14323 4029 14335 4063
rect 14550 4060 14556 4072
rect 14511 4032 14556 4060
rect 14277 4023 14335 4029
rect 8018 3884 8024 3936
rect 8076 3924 8082 3936
rect 8297 3927 8355 3933
rect 8297 3924 8309 3927
rect 8076 3896 8309 3924
rect 8076 3884 8082 3896
rect 8297 3893 8309 3896
rect 8343 3924 8355 3927
rect 8849 3927 8907 3933
rect 8849 3924 8861 3927
rect 8343 3896 8861 3924
rect 8343 3893 8355 3896
rect 8297 3887 8355 3893
rect 8849 3893 8861 3896
rect 8895 3924 8907 3927
rect 9306 3924 9312 3936
rect 8895 3896 9312 3924
rect 8895 3893 8907 3896
rect 8849 3887 8907 3893
rect 9306 3884 9312 3896
rect 9364 3924 9370 3936
rect 9401 3927 9459 3933
rect 9401 3924 9413 3927
rect 9364 3896 9413 3924
rect 9364 3884 9370 3896
rect 9401 3893 9413 3896
rect 9447 3893 9459 3927
rect 9401 3887 9459 3893
rect 10597 3927 10655 3933
rect 10597 3893 10609 3927
rect 10643 3924 10655 3927
rect 12066 3924 12072 3936
rect 10643 3896 12072 3924
rect 10643 3893 10655 3896
rect 10597 3887 10655 3893
rect 12066 3884 12072 3896
rect 12124 3884 12130 3936
rect 14292 3924 14320 4023
rect 14550 4020 14556 4032
rect 14608 4020 14614 4072
rect 17126 4060 17132 4072
rect 17087 4032 17132 4060
rect 17126 4020 17132 4032
rect 17184 4020 17190 4072
rect 17218 4020 17224 4072
rect 17276 4060 17282 4072
rect 17862 4060 17868 4072
rect 17276 4032 17868 4060
rect 17276 4020 17282 4032
rect 17862 4020 17868 4032
rect 17920 4020 17926 4072
rect 18601 4063 18659 4069
rect 18601 4029 18613 4063
rect 18647 4029 18659 4063
rect 18874 4060 18880 4072
rect 18835 4032 18880 4060
rect 18601 4023 18659 4029
rect 18506 3992 18512 4004
rect 15580 3964 18512 3992
rect 14550 3924 14556 3936
rect 14292 3896 14556 3924
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 15580 3924 15608 3964
rect 18506 3952 18512 3964
rect 18564 3952 18570 4004
rect 18616 3992 18644 4023
rect 18874 4020 18880 4032
rect 18932 4020 18938 4072
rect 18966 4020 18972 4072
rect 19024 4060 19030 4072
rect 20088 4060 20116 4100
rect 21266 4088 21272 4100
rect 21324 4088 21330 4140
rect 23753 4131 23811 4137
rect 23753 4097 23765 4131
rect 23799 4128 23811 4131
rect 23842 4128 23848 4140
rect 23799 4100 23848 4128
rect 23799 4097 23811 4100
rect 23753 4091 23811 4097
rect 23842 4088 23848 4100
rect 23900 4128 23906 4140
rect 24213 4131 24271 4137
rect 24213 4128 24225 4131
rect 23900 4100 24225 4128
rect 23900 4088 23906 4100
rect 24213 4097 24225 4100
rect 24259 4097 24271 4131
rect 24213 4091 24271 4097
rect 25774 4088 25780 4140
rect 25832 4128 25838 4140
rect 27525 4131 27583 4137
rect 27525 4128 27537 4131
rect 25832 4100 27537 4128
rect 25832 4088 25838 4100
rect 27525 4097 27537 4100
rect 27571 4097 27583 4131
rect 27525 4091 27583 4097
rect 27617 4131 27675 4137
rect 27617 4097 27629 4131
rect 27663 4128 27675 4131
rect 27982 4128 27988 4140
rect 27663 4100 27988 4128
rect 27663 4097 27675 4100
rect 27617 4091 27675 4097
rect 27982 4088 27988 4100
rect 28040 4088 28046 4140
rect 28166 4088 28172 4140
rect 28224 4128 28230 4140
rect 28261 4131 28319 4137
rect 28261 4128 28273 4131
rect 28224 4100 28273 4128
rect 28224 4088 28230 4100
rect 28261 4097 28273 4100
rect 28307 4128 28319 4131
rect 28994 4128 29000 4140
rect 28307 4100 29000 4128
rect 28307 4097 28319 4100
rect 28261 4091 28319 4097
rect 28994 4088 29000 4100
rect 29052 4088 29058 4140
rect 29086 4088 29092 4140
rect 29144 4128 29150 4140
rect 29288 4137 29316 4168
rect 30006 4156 30012 4168
rect 30064 4156 30070 4208
rect 29181 4131 29239 4137
rect 29181 4128 29193 4131
rect 29144 4100 29193 4128
rect 29144 4088 29150 4100
rect 29181 4097 29193 4100
rect 29227 4097 29239 4131
rect 29181 4091 29239 4097
rect 29273 4131 29331 4137
rect 29273 4097 29285 4131
rect 29319 4097 29331 4131
rect 29273 4091 29331 4097
rect 29822 4088 29828 4140
rect 29880 4128 29886 4140
rect 29917 4131 29975 4137
rect 29917 4128 29929 4131
rect 29880 4100 29929 4128
rect 29880 4088 29886 4100
rect 29917 4097 29929 4100
rect 29963 4128 29975 4131
rect 30282 4128 30288 4140
rect 29963 4100 30288 4128
rect 29963 4097 29975 4100
rect 29917 4091 29975 4097
rect 30282 4088 30288 4100
rect 30340 4088 30346 4140
rect 30377 4131 30435 4137
rect 30377 4097 30389 4131
rect 30423 4128 30435 4131
rect 30558 4128 30564 4140
rect 30423 4100 30564 4128
rect 30423 4097 30435 4100
rect 30377 4091 30435 4097
rect 30558 4088 30564 4100
rect 30616 4088 30622 4140
rect 31202 4128 31208 4140
rect 31163 4100 31208 4128
rect 31202 4088 31208 4100
rect 31260 4088 31266 4140
rect 32309 4131 32367 4137
rect 32309 4097 32321 4131
rect 32355 4128 32367 4131
rect 33042 4128 33048 4140
rect 32355 4100 33048 4128
rect 32355 4097 32367 4100
rect 32309 4091 32367 4097
rect 33042 4088 33048 4100
rect 33100 4128 33106 4140
rect 33229 4131 33287 4137
rect 33229 4128 33241 4131
rect 33100 4100 33241 4128
rect 33100 4088 33106 4100
rect 33229 4097 33241 4100
rect 33275 4097 33287 4131
rect 33229 4091 33287 4097
rect 19024 4032 20116 4060
rect 19024 4020 19030 4032
rect 20346 4020 20352 4072
rect 20404 4060 20410 4072
rect 20625 4063 20683 4069
rect 20625 4060 20637 4063
rect 20404 4032 20637 4060
rect 20404 4020 20410 4032
rect 20625 4029 20637 4032
rect 20671 4029 20683 4063
rect 20625 4023 20683 4029
rect 20806 4020 20812 4072
rect 20864 4060 20870 4072
rect 22005 4063 22063 4069
rect 22005 4060 22017 4063
rect 20864 4032 22017 4060
rect 20864 4020 20870 4032
rect 22005 4029 22017 4032
rect 22051 4029 22063 4063
rect 22005 4023 22063 4029
rect 22094 4020 22100 4072
rect 22152 4060 22158 4072
rect 23474 4060 23480 4072
rect 22152 4032 23480 4060
rect 22152 4020 22158 4032
rect 23474 4020 23480 4032
rect 23532 4020 23538 4072
rect 26326 4060 26332 4072
rect 24320 4032 26332 4060
rect 18616 3964 18736 3992
rect 14792 3896 15608 3924
rect 14792 3884 14798 3896
rect 15654 3884 15660 3936
rect 15712 3924 15718 3936
rect 15930 3924 15936 3936
rect 15712 3896 15936 3924
rect 15712 3884 15718 3896
rect 15930 3884 15936 3896
rect 15988 3884 15994 3936
rect 16942 3884 16948 3936
rect 17000 3924 17006 3936
rect 18598 3924 18604 3936
rect 17000 3896 18604 3924
rect 17000 3884 17006 3896
rect 18598 3884 18604 3896
rect 18656 3884 18662 3936
rect 18708 3924 18736 3964
rect 19886 3952 19892 4004
rect 19944 3992 19950 4004
rect 22370 3992 22376 4004
rect 19944 3964 22376 3992
rect 19944 3952 19950 3964
rect 22370 3952 22376 3964
rect 22428 3952 22434 4004
rect 19334 3924 19340 3936
rect 18708 3896 19340 3924
rect 19334 3884 19340 3896
rect 19392 3884 19398 3936
rect 20346 3884 20352 3936
rect 20404 3924 20410 3936
rect 24320 3924 24348 4032
rect 26326 4020 26332 4032
rect 26384 4020 26390 4072
rect 26418 4020 26424 4072
rect 26476 4060 26482 4072
rect 31665 4063 31723 4069
rect 31665 4060 31677 4063
rect 26476 4032 31677 4060
rect 26476 4020 26482 4032
rect 31665 4029 31677 4032
rect 31711 4029 31723 4063
rect 32490 4060 32496 4072
rect 32451 4032 32496 4060
rect 31665 4023 31723 4029
rect 32490 4020 32496 4032
rect 32548 4020 32554 4072
rect 26510 3952 26516 4004
rect 26568 3992 26574 4004
rect 26568 3964 26613 3992
rect 26568 3952 26574 3964
rect 27430 3952 27436 4004
rect 27488 3992 27494 4004
rect 30469 3995 30527 4001
rect 30469 3992 30481 3995
rect 27488 3964 30481 3992
rect 27488 3952 27494 3964
rect 30469 3961 30481 3964
rect 30515 3961 30527 3995
rect 31110 3992 31116 4004
rect 31071 3964 31116 3992
rect 30469 3955 30527 3961
rect 31110 3952 31116 3964
rect 31168 3952 31174 4004
rect 31754 3952 31760 4004
rect 31812 3992 31818 4004
rect 38010 3992 38016 4004
rect 31812 3964 38016 3992
rect 31812 3952 31818 3964
rect 38010 3952 38016 3964
rect 38068 3952 38074 4004
rect 20404 3896 24348 3924
rect 20404 3884 20410 3896
rect 24578 3884 24584 3936
rect 24636 3924 24642 3936
rect 25961 3927 26019 3933
rect 25961 3924 25973 3927
rect 24636 3896 25973 3924
rect 24636 3884 24642 3896
rect 25961 3893 25973 3896
rect 26007 3893 26019 3927
rect 28166 3924 28172 3936
rect 28127 3896 28172 3924
rect 25961 3887 26019 3893
rect 28166 3884 28172 3896
rect 28224 3884 28230 3936
rect 28442 3884 28448 3936
rect 28500 3924 28506 3936
rect 29825 3927 29883 3933
rect 29825 3924 29837 3927
rect 28500 3896 29837 3924
rect 28500 3884 28506 3896
rect 29825 3893 29837 3896
rect 29871 3893 29883 3927
rect 29825 3887 29883 3893
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 9217 3723 9275 3729
rect 9217 3689 9229 3723
rect 9263 3720 9275 3723
rect 12434 3720 12440 3732
rect 9263 3692 12440 3720
rect 9263 3689 9275 3692
rect 9217 3683 9275 3689
rect 12434 3680 12440 3692
rect 12492 3680 12498 3732
rect 12618 3680 12624 3732
rect 12676 3720 12682 3732
rect 17126 3720 17132 3732
rect 12676 3692 17132 3720
rect 12676 3680 12682 3692
rect 17126 3680 17132 3692
rect 17184 3680 17190 3732
rect 17218 3680 17224 3732
rect 17276 3720 17282 3732
rect 20257 3723 20315 3729
rect 20257 3720 20269 3723
rect 17276 3692 20269 3720
rect 17276 3680 17282 3692
rect 20257 3689 20269 3692
rect 20303 3689 20315 3723
rect 20257 3683 20315 3689
rect 23290 3680 23296 3732
rect 23348 3720 23354 3732
rect 28166 3720 28172 3732
rect 23348 3692 28172 3720
rect 23348 3680 23354 3692
rect 28166 3680 28172 3692
rect 28224 3680 28230 3732
rect 28718 3680 28724 3732
rect 28776 3720 28782 3732
rect 28813 3723 28871 3729
rect 28813 3720 28825 3723
rect 28776 3692 28825 3720
rect 28776 3680 28782 3692
rect 28813 3689 28825 3692
rect 28859 3689 28871 3723
rect 28813 3683 28871 3689
rect 30374 3680 30380 3732
rect 30432 3720 30438 3732
rect 32401 3723 32459 3729
rect 32401 3720 32413 3723
rect 30432 3692 32413 3720
rect 30432 3680 30438 3692
rect 32401 3689 32413 3692
rect 32447 3689 32459 3723
rect 32401 3683 32459 3689
rect 34790 3680 34796 3732
rect 34848 3720 34854 3732
rect 34885 3723 34943 3729
rect 34885 3720 34897 3723
rect 34848 3692 34897 3720
rect 34848 3680 34854 3692
rect 34885 3689 34897 3692
rect 34931 3689 34943 3723
rect 34885 3683 34943 3689
rect 4430 3612 4436 3664
rect 4488 3652 4494 3664
rect 4801 3655 4859 3661
rect 4801 3652 4813 3655
rect 4488 3624 4813 3652
rect 4488 3612 4494 3624
rect 4801 3621 4813 3624
rect 4847 3652 4859 3655
rect 8110 3652 8116 3664
rect 4847 3624 8116 3652
rect 4847 3621 4859 3624
rect 4801 3615 4859 3621
rect 8110 3612 8116 3624
rect 8168 3652 8174 3664
rect 11974 3652 11980 3664
rect 8168 3624 11980 3652
rect 8168 3612 8174 3624
rect 11974 3612 11980 3624
rect 12032 3612 12038 3664
rect 13262 3612 13268 3664
rect 13320 3652 13326 3664
rect 13725 3655 13783 3661
rect 13725 3652 13737 3655
rect 13320 3624 13737 3652
rect 13320 3612 13326 3624
rect 13725 3621 13737 3624
rect 13771 3621 13783 3655
rect 13725 3615 13783 3621
rect 14642 3612 14648 3664
rect 14700 3652 14706 3664
rect 14700 3624 14780 3652
rect 14700 3612 14706 3624
rect 8570 3584 8576 3596
rect 8483 3556 8576 3584
rect 8570 3544 8576 3556
rect 8628 3584 8634 3596
rect 11882 3584 11888 3596
rect 8628 3556 11888 3584
rect 8628 3544 8634 3556
rect 11882 3544 11888 3556
rect 11940 3544 11946 3596
rect 12250 3584 12256 3596
rect 12211 3556 12256 3584
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 12710 3544 12716 3596
rect 12768 3584 12774 3596
rect 14752 3584 14780 3624
rect 18782 3612 18788 3664
rect 18840 3652 18846 3664
rect 20346 3652 20352 3664
rect 18840 3624 20352 3652
rect 18840 3612 18846 3624
rect 20346 3612 20352 3624
rect 20404 3612 20410 3664
rect 23750 3612 23756 3664
rect 23808 3652 23814 3664
rect 26329 3655 26387 3661
rect 23808 3624 24716 3652
rect 23808 3612 23814 3624
rect 14921 3587 14979 3593
rect 14921 3584 14933 3587
rect 12768 3556 13584 3584
rect 14752 3556 14933 3584
rect 12768 3544 12774 3556
rect 1578 3516 1584 3528
rect 1539 3488 1584 3516
rect 1578 3476 1584 3488
rect 1636 3516 1642 3528
rect 2225 3519 2283 3525
rect 2225 3516 2237 3519
rect 1636 3488 2237 3516
rect 1636 3476 1642 3488
rect 2225 3485 2237 3488
rect 2271 3485 2283 3519
rect 2225 3479 2283 3485
rect 8202 3476 8208 3528
rect 8260 3516 8266 3528
rect 11425 3519 11483 3525
rect 11425 3516 11437 3519
rect 8260 3488 11437 3516
rect 8260 3476 8266 3488
rect 11425 3485 11437 3488
rect 11471 3485 11483 3519
rect 11425 3479 11483 3485
rect 11517 3519 11575 3525
rect 11517 3485 11529 3519
rect 11563 3516 11575 3519
rect 11790 3516 11796 3528
rect 11563 3488 11796 3516
rect 11563 3485 11575 3488
rect 11517 3479 11575 3485
rect 11790 3476 11796 3488
rect 11848 3476 11854 3528
rect 11977 3519 12035 3525
rect 11977 3485 11989 3519
rect 12023 3485 12035 3519
rect 11977 3479 12035 3485
rect 8570 3448 8576 3460
rect 1780 3420 8576 3448
rect 1780 3389 1808 3420
rect 8570 3408 8576 3420
rect 8628 3408 8634 3460
rect 11992 3448 12020 3479
rect 13354 3476 13360 3528
rect 13412 3476 13418 3528
rect 12342 3448 12348 3460
rect 11808 3420 12348 3448
rect 1765 3383 1823 3389
rect 1765 3349 1777 3383
rect 1811 3349 1823 3383
rect 7466 3380 7472 3392
rect 7427 3352 7472 3380
rect 1765 3343 1823 3349
rect 7466 3340 7472 3352
rect 7524 3340 7530 3392
rect 8018 3380 8024 3392
rect 7979 3352 8024 3380
rect 8018 3340 8024 3352
rect 8076 3340 8082 3392
rect 9769 3383 9827 3389
rect 9769 3349 9781 3383
rect 9815 3380 9827 3383
rect 10229 3383 10287 3389
rect 10229 3380 10241 3383
rect 9815 3352 10241 3380
rect 9815 3349 9827 3352
rect 9769 3343 9827 3349
rect 10229 3349 10241 3352
rect 10275 3380 10287 3383
rect 10781 3383 10839 3389
rect 10781 3380 10793 3383
rect 10275 3352 10793 3380
rect 10275 3349 10287 3352
rect 10229 3343 10287 3349
rect 10781 3349 10793 3352
rect 10827 3380 10839 3383
rect 11808 3380 11836 3420
rect 12342 3408 12348 3420
rect 12400 3408 12406 3460
rect 13556 3448 13584 3556
rect 14921 3553 14933 3556
rect 14967 3553 14979 3587
rect 14921 3547 14979 3553
rect 15010 3544 15016 3596
rect 15068 3584 15074 3596
rect 16853 3587 16911 3593
rect 15068 3556 16344 3584
rect 15068 3544 15074 3556
rect 14550 3476 14556 3528
rect 14608 3516 14614 3528
rect 14645 3519 14703 3525
rect 14645 3516 14657 3519
rect 14608 3488 14657 3516
rect 14608 3476 14614 3488
rect 14645 3485 14657 3488
rect 14691 3485 14703 3519
rect 14645 3479 14703 3485
rect 15194 3448 15200 3460
rect 13556 3420 15200 3448
rect 15194 3408 15200 3420
rect 15252 3408 15258 3460
rect 16206 3448 16212 3460
rect 16146 3420 16212 3448
rect 16206 3408 16212 3420
rect 16264 3408 16270 3460
rect 16316 3448 16344 3556
rect 16853 3553 16865 3587
rect 16899 3584 16911 3587
rect 17126 3584 17132 3596
rect 16899 3556 17132 3584
rect 16899 3553 16911 3556
rect 16853 3547 16911 3553
rect 17126 3544 17132 3556
rect 17184 3544 17190 3596
rect 19886 3584 19892 3596
rect 18248 3556 19892 3584
rect 18248 3502 18276 3556
rect 19886 3544 19892 3556
rect 19944 3544 19950 3596
rect 20622 3544 20628 3596
rect 20680 3584 20686 3596
rect 20993 3587 21051 3593
rect 20993 3584 21005 3587
rect 20680 3556 21005 3584
rect 20680 3544 20686 3556
rect 20993 3553 21005 3556
rect 21039 3553 21051 3587
rect 20993 3547 21051 3553
rect 23842 3544 23848 3596
rect 23900 3584 23906 3596
rect 24581 3587 24639 3593
rect 24581 3584 24593 3587
rect 23900 3556 24593 3584
rect 23900 3544 23906 3556
rect 24581 3553 24593 3556
rect 24627 3553 24639 3587
rect 24688 3584 24716 3624
rect 26329 3621 26341 3655
rect 26375 3652 26387 3655
rect 26418 3652 26424 3664
rect 26375 3624 26424 3652
rect 26375 3621 26387 3624
rect 26329 3615 26387 3621
rect 26418 3612 26424 3624
rect 26476 3652 26482 3664
rect 26602 3652 26608 3664
rect 26476 3624 26608 3652
rect 26476 3612 26482 3624
rect 26602 3612 26608 3624
rect 26660 3612 26666 3664
rect 26973 3655 27031 3661
rect 26973 3621 26985 3655
rect 27019 3652 27031 3655
rect 31754 3652 31760 3664
rect 27019 3624 31760 3652
rect 27019 3621 27031 3624
rect 26973 3615 27031 3621
rect 31754 3612 31760 3624
rect 31812 3612 31818 3664
rect 37918 3612 37924 3664
rect 37976 3652 37982 3664
rect 38013 3655 38071 3661
rect 38013 3652 38025 3655
rect 37976 3624 38025 3652
rect 37976 3612 37982 3624
rect 38013 3621 38025 3624
rect 38059 3621 38071 3655
rect 38013 3615 38071 3621
rect 24857 3587 24915 3593
rect 24857 3584 24869 3587
rect 24688 3556 24869 3584
rect 24581 3547 24639 3553
rect 24857 3553 24869 3556
rect 24903 3553 24915 3587
rect 24857 3547 24915 3553
rect 25498 3544 25504 3596
rect 25556 3584 25562 3596
rect 29825 3587 29883 3593
rect 29825 3584 29837 3587
rect 25556 3556 29837 3584
rect 25556 3544 25562 3556
rect 29825 3553 29837 3556
rect 29871 3553 29883 3587
rect 29825 3547 29883 3553
rect 30006 3544 30012 3596
rect 30064 3584 30070 3596
rect 32950 3584 32956 3596
rect 30064 3556 31248 3584
rect 32911 3556 32956 3584
rect 30064 3544 30070 3556
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 18524 3488 19441 3516
rect 17129 3451 17187 3457
rect 17129 3448 17141 3451
rect 16316 3420 17141 3448
rect 17129 3417 17141 3420
rect 17175 3417 17187 3451
rect 17129 3411 17187 3417
rect 10827 3352 11836 3380
rect 10827 3349 10839 3352
rect 10781 3343 10839 3349
rect 14826 3340 14832 3392
rect 14884 3380 14890 3392
rect 16393 3383 16451 3389
rect 16393 3380 16405 3383
rect 14884 3352 16405 3380
rect 14884 3340 14890 3352
rect 16393 3349 16405 3352
rect 16439 3380 16451 3383
rect 17310 3380 17316 3392
rect 16439 3352 17316 3380
rect 16439 3349 16451 3352
rect 16393 3343 16451 3349
rect 17310 3340 17316 3352
rect 17368 3340 17374 3392
rect 17494 3340 17500 3392
rect 17552 3380 17558 3392
rect 18524 3380 18552 3488
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 20438 3516 20444 3528
rect 20399 3488 20444 3516
rect 19429 3479 19487 3485
rect 20438 3476 20444 3488
rect 20496 3476 20502 3528
rect 23198 3516 23204 3528
rect 22402 3488 23204 3516
rect 23198 3476 23204 3488
rect 23256 3476 23262 3528
rect 23753 3519 23811 3525
rect 23753 3485 23765 3519
rect 23799 3516 23811 3519
rect 23934 3516 23940 3528
rect 23799 3488 23940 3516
rect 23799 3485 23811 3488
rect 23753 3479 23811 3485
rect 23934 3476 23940 3488
rect 23992 3476 23998 3528
rect 26786 3516 26792 3528
rect 26699 3488 26792 3516
rect 26786 3476 26792 3488
rect 26844 3516 26850 3528
rect 27338 3516 27344 3528
rect 26844 3488 27344 3516
rect 26844 3476 26850 3488
rect 27338 3476 27344 3488
rect 27396 3476 27402 3528
rect 27522 3516 27528 3528
rect 27483 3488 27528 3516
rect 27522 3476 27528 3488
rect 27580 3476 27586 3528
rect 27617 3519 27675 3525
rect 27617 3485 27629 3519
rect 27663 3516 27675 3519
rect 28074 3516 28080 3528
rect 27663 3488 28080 3516
rect 27663 3485 27675 3488
rect 27617 3479 27675 3485
rect 28074 3476 28080 3488
rect 28132 3476 28138 3528
rect 28261 3519 28319 3525
rect 28261 3485 28273 3519
rect 28307 3516 28319 3519
rect 28307 3488 28672 3516
rect 28307 3485 28319 3488
rect 28261 3479 28319 3485
rect 18598 3408 18604 3460
rect 18656 3448 18662 3460
rect 18877 3451 18935 3457
rect 18877 3448 18889 3451
rect 18656 3420 18889 3448
rect 18656 3408 18662 3420
rect 18877 3417 18889 3420
rect 18923 3417 18935 3451
rect 18877 3411 18935 3417
rect 18966 3408 18972 3460
rect 19024 3448 19030 3460
rect 21174 3448 21180 3460
rect 19024 3420 21180 3448
rect 19024 3408 19030 3420
rect 21174 3408 21180 3420
rect 21232 3408 21238 3460
rect 21269 3451 21327 3457
rect 21269 3417 21281 3451
rect 21315 3448 21327 3451
rect 21358 3448 21364 3460
rect 21315 3420 21364 3448
rect 21315 3417 21327 3420
rect 21269 3411 21327 3417
rect 21358 3408 21364 3420
rect 21416 3408 21422 3460
rect 22922 3408 22928 3460
rect 22980 3448 22986 3460
rect 23017 3451 23075 3457
rect 23017 3448 23029 3451
rect 22980 3420 23029 3448
rect 22980 3408 22986 3420
rect 23017 3417 23029 3420
rect 23063 3417 23075 3451
rect 28442 3448 28448 3460
rect 26082 3420 28448 3448
rect 23017 3411 23075 3417
rect 28442 3408 28448 3420
rect 28500 3408 28506 3460
rect 28644 3448 28672 3488
rect 28810 3476 28816 3528
rect 28868 3516 28874 3528
rect 28913 3519 28971 3525
rect 28913 3516 28925 3519
rect 28868 3488 28925 3516
rect 28868 3476 28874 3488
rect 28913 3485 28925 3488
rect 28959 3485 28971 3519
rect 29914 3516 29920 3528
rect 29875 3488 29920 3516
rect 28913 3479 28971 3485
rect 29914 3476 29920 3488
rect 29972 3476 29978 3528
rect 30282 3476 30288 3528
rect 30340 3516 30346 3528
rect 30561 3519 30619 3525
rect 30561 3516 30573 3519
rect 30340 3488 30573 3516
rect 30340 3476 30346 3488
rect 30561 3485 30573 3488
rect 30607 3485 30619 3519
rect 30561 3479 30619 3485
rect 31018 3476 31024 3528
rect 31076 3516 31082 3528
rect 31220 3525 31248 3556
rect 32950 3544 32956 3556
rect 33008 3544 33014 3596
rect 31113 3519 31171 3525
rect 31113 3516 31125 3519
rect 31076 3488 31125 3516
rect 31076 3476 31082 3488
rect 31113 3485 31125 3488
rect 31159 3485 31171 3519
rect 31113 3479 31171 3485
rect 31205 3519 31263 3525
rect 31205 3485 31217 3519
rect 31251 3516 31263 3519
rect 31846 3516 31852 3528
rect 31251 3488 31754 3516
rect 31807 3488 31852 3516
rect 31251 3485 31263 3488
rect 31205 3479 31263 3485
rect 31294 3448 31300 3460
rect 28644 3420 31300 3448
rect 31294 3408 31300 3420
rect 31352 3408 31358 3460
rect 31726 3448 31754 3488
rect 31846 3476 31852 3488
rect 31904 3476 31910 3528
rect 32490 3516 32496 3528
rect 32403 3488 32496 3516
rect 32490 3476 32496 3488
rect 32548 3476 32554 3528
rect 32508 3448 32536 3476
rect 31726 3420 32536 3448
rect 37553 3451 37611 3457
rect 37553 3417 37565 3451
rect 37599 3448 37611 3451
rect 38197 3451 38255 3457
rect 38197 3448 38209 3451
rect 37599 3420 38209 3448
rect 37599 3417 37611 3420
rect 37553 3411 37611 3417
rect 38197 3417 38209 3420
rect 38243 3448 38255 3451
rect 39298 3448 39304 3460
rect 38243 3420 39304 3448
rect 38243 3417 38255 3420
rect 38197 3411 38255 3417
rect 39298 3408 39304 3420
rect 39356 3408 39362 3460
rect 17552 3352 18552 3380
rect 17552 3340 17558 3352
rect 18690 3340 18696 3392
rect 18748 3380 18754 3392
rect 19613 3383 19671 3389
rect 19613 3380 19625 3383
rect 18748 3352 19625 3380
rect 18748 3340 18754 3352
rect 19613 3349 19625 3352
rect 19659 3349 19671 3383
rect 19613 3343 19671 3349
rect 21910 3340 21916 3392
rect 21968 3380 21974 3392
rect 23569 3383 23627 3389
rect 23569 3380 23581 3383
rect 21968 3352 23581 3380
rect 21968 3340 21974 3352
rect 23569 3349 23581 3352
rect 23615 3349 23627 3383
rect 23569 3343 23627 3349
rect 28169 3383 28227 3389
rect 28169 3349 28181 3383
rect 28215 3380 28227 3383
rect 28258 3380 28264 3392
rect 28215 3352 28264 3380
rect 28215 3349 28227 3352
rect 28169 3343 28227 3349
rect 28258 3340 28264 3352
rect 28316 3340 28322 3392
rect 30466 3380 30472 3392
rect 30427 3352 30472 3380
rect 30466 3340 30472 3352
rect 30524 3340 30530 3392
rect 31754 3380 31760 3392
rect 31715 3352 31760 3380
rect 31754 3340 31760 3352
rect 31812 3340 31818 3392
rect 33594 3380 33600 3392
rect 33555 3352 33600 3380
rect 33594 3340 33600 3352
rect 33652 3340 33658 3392
rect 34054 3380 34060 3392
rect 34015 3352 34060 3380
rect 34054 3340 34060 3352
rect 34112 3340 34118 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 2777 3179 2835 3185
rect 2777 3145 2789 3179
rect 2823 3176 2835 3179
rect 2866 3176 2872 3188
rect 2823 3148 2872 3176
rect 2823 3145 2835 3148
rect 2777 3139 2835 3145
rect 2866 3136 2872 3148
rect 2924 3136 2930 3188
rect 3326 3176 3332 3188
rect 3287 3148 3332 3176
rect 3326 3136 3332 3148
rect 3384 3136 3390 3188
rect 7193 3179 7251 3185
rect 7193 3145 7205 3179
rect 7239 3176 7251 3179
rect 11146 3176 11152 3188
rect 7239 3148 11152 3176
rect 7239 3145 7251 3148
rect 7193 3139 7251 3145
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 11793 3179 11851 3185
rect 11793 3145 11805 3179
rect 11839 3176 11851 3179
rect 12158 3176 12164 3188
rect 11839 3148 12164 3176
rect 11839 3145 11851 3148
rect 11793 3139 11851 3145
rect 12158 3136 12164 3148
rect 12216 3136 12222 3188
rect 12250 3136 12256 3188
rect 12308 3176 12314 3188
rect 12308 3148 12756 3176
rect 12308 3136 12314 3148
rect 10042 3108 10048 3120
rect 5276 3080 10048 3108
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3009 1915 3043
rect 4430 3040 4436 3052
rect 4391 3012 4436 3040
rect 1857 3003 1915 3009
rect 1872 2972 1900 3003
rect 4430 3000 4436 3012
rect 4488 3000 4494 3052
rect 5276 3049 5304 3080
rect 10042 3068 10048 3080
rect 10100 3068 10106 3120
rect 10318 3108 10324 3120
rect 10279 3080 10324 3108
rect 10318 3068 10324 3080
rect 10376 3068 10382 3120
rect 11606 3068 11612 3120
rect 11664 3108 11670 3120
rect 12621 3111 12679 3117
rect 12621 3108 12633 3111
rect 11664 3080 12633 3108
rect 11664 3068 11670 3080
rect 12621 3077 12633 3080
rect 12667 3077 12679 3111
rect 12728 3108 12756 3148
rect 12802 3136 12808 3188
rect 12860 3176 12866 3188
rect 16301 3179 16359 3185
rect 16301 3176 16313 3179
rect 12860 3148 16313 3176
rect 12860 3136 12866 3148
rect 16301 3145 16313 3148
rect 16347 3145 16359 3179
rect 16301 3139 16359 3145
rect 12894 3108 12900 3120
rect 12728 3080 12900 3108
rect 12621 3071 12679 3077
rect 12894 3068 12900 3080
rect 12952 3068 12958 3120
rect 13906 3068 13912 3120
rect 13964 3108 13970 3120
rect 14829 3111 14887 3117
rect 14829 3108 14841 3111
rect 13964 3080 14841 3108
rect 13964 3068 13970 3080
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 7466 3000 7472 3052
rect 7524 3040 7530 3052
rect 9309 3043 9367 3049
rect 9309 3040 9321 3043
rect 7524 3012 9321 3040
rect 7524 3000 7530 3012
rect 9309 3009 9321 3012
rect 9355 3009 9367 3043
rect 9309 3003 9367 3009
rect 9401 3043 9459 3049
rect 9401 3009 9413 3043
rect 9447 3040 9459 3043
rect 10873 3043 10931 3049
rect 10873 3040 10885 3043
rect 9447 3012 10885 3040
rect 9447 3009 9459 3012
rect 9401 3003 9459 3009
rect 10873 3009 10885 3012
rect 10919 3009 10931 3043
rect 10873 3003 10931 3009
rect 8849 2975 8907 2981
rect 1872 2944 2774 2972
rect 2746 2904 2774 2944
rect 8849 2941 8861 2975
rect 8895 2972 8907 2975
rect 8938 2972 8944 2984
rect 8895 2944 8944 2972
rect 8895 2941 8907 2944
rect 8849 2935 8907 2941
rect 8938 2932 8944 2944
rect 8996 2932 9002 2984
rect 9324 2972 9352 3003
rect 10962 3000 10968 3052
rect 11020 3040 11026 3052
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 11020 3012 11713 3040
rect 11020 3000 11026 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 12342 3040 12348 3052
rect 12303 3012 12348 3040
rect 11701 3003 11759 3009
rect 12342 3000 12348 3012
rect 12400 3000 12406 3052
rect 13722 3000 13728 3052
rect 13780 3000 13786 3052
rect 12710 2972 12716 2984
rect 9324 2944 12716 2972
rect 12710 2932 12716 2944
rect 12768 2932 12774 2984
rect 12986 2932 12992 2984
rect 13044 2972 13050 2984
rect 14090 2972 14096 2984
rect 13044 2944 13768 2972
rect 14051 2944 14096 2972
rect 13044 2932 13050 2944
rect 5077 2907 5135 2913
rect 5077 2904 5089 2907
rect 2746 2876 5089 2904
rect 5077 2873 5089 2876
rect 5123 2873 5135 2907
rect 5077 2867 5135 2873
rect 6641 2907 6699 2913
rect 6641 2873 6653 2907
rect 6687 2904 6699 2907
rect 9858 2904 9864 2916
rect 6687 2876 9864 2904
rect 6687 2873 6699 2876
rect 6641 2867 6699 2873
rect 9858 2864 9864 2876
rect 9916 2864 9922 2916
rect 10042 2864 10048 2916
rect 10100 2904 10106 2916
rect 10962 2904 10968 2916
rect 10100 2876 10968 2904
rect 10100 2864 10106 2876
rect 10962 2864 10968 2876
rect 11020 2864 11026 2916
rect 11146 2864 11152 2916
rect 11204 2904 11210 2916
rect 11204 2876 11744 2904
rect 11204 2864 11210 2876
rect 1670 2836 1676 2848
rect 1631 2808 1676 2836
rect 1670 2796 1676 2808
rect 1728 2796 1734 2848
rect 4614 2836 4620 2848
rect 4575 2808 4620 2836
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 7745 2839 7803 2845
rect 7745 2805 7757 2839
rect 7791 2836 7803 2839
rect 8018 2836 8024 2848
rect 7791 2808 8024 2836
rect 7791 2805 7803 2808
rect 7745 2799 7803 2805
rect 8018 2796 8024 2808
rect 8076 2836 8082 2848
rect 8205 2839 8263 2845
rect 8205 2836 8217 2839
rect 8076 2808 8217 2836
rect 8076 2796 8082 2808
rect 8205 2805 8217 2808
rect 8251 2805 8263 2839
rect 8205 2799 8263 2805
rect 8938 2796 8944 2848
rect 8996 2836 9002 2848
rect 10870 2836 10876 2848
rect 8996 2808 10876 2836
rect 8996 2796 9002 2808
rect 10870 2796 10876 2808
rect 10928 2796 10934 2848
rect 11057 2839 11115 2845
rect 11057 2805 11069 2839
rect 11103 2836 11115 2839
rect 11606 2836 11612 2848
rect 11103 2808 11612 2836
rect 11103 2805 11115 2808
rect 11057 2799 11115 2805
rect 11606 2796 11612 2808
rect 11664 2796 11670 2848
rect 11716 2836 11744 2876
rect 13630 2836 13636 2848
rect 11716 2808 13636 2836
rect 13630 2796 13636 2808
rect 13688 2796 13694 2848
rect 13740 2836 13768 2944
rect 14090 2932 14096 2944
rect 14148 2932 14154 2984
rect 14384 2904 14412 3080
rect 14829 3077 14841 3080
rect 14875 3077 14887 3111
rect 16316 3108 16344 3139
rect 17126 3136 17132 3188
rect 17184 3176 17190 3188
rect 19334 3176 19340 3188
rect 17184 3148 19340 3176
rect 17184 3136 17190 3148
rect 16316 3080 17172 3108
rect 14829 3071 14887 3077
rect 15962 3012 17080 3040
rect 14550 2972 14556 2984
rect 14511 2944 14556 2972
rect 14550 2932 14556 2944
rect 14608 2932 14614 2984
rect 16942 2972 16948 2984
rect 14660 2944 16948 2972
rect 14660 2904 14688 2944
rect 16942 2932 16948 2944
rect 17000 2932 17006 2984
rect 14384 2876 14688 2904
rect 16114 2836 16120 2848
rect 13740 2808 16120 2836
rect 16114 2796 16120 2808
rect 16172 2796 16178 2848
rect 17052 2836 17080 3012
rect 17144 2972 17172 3080
rect 17236 3049 17264 3148
rect 19334 3136 19340 3148
rect 19392 3136 19398 3188
rect 19794 3136 19800 3188
rect 19852 3176 19858 3188
rect 32401 3179 32459 3185
rect 32401 3176 32413 3179
rect 19852 3148 32413 3176
rect 19852 3136 19858 3148
rect 32401 3145 32413 3148
rect 32447 3145 32459 3179
rect 32401 3139 32459 3145
rect 18782 3108 18788 3120
rect 18722 3080 18788 3108
rect 18782 3068 18788 3080
rect 18840 3068 18846 3120
rect 19610 3068 19616 3120
rect 19668 3108 19674 3120
rect 19705 3111 19763 3117
rect 19705 3108 19717 3111
rect 19668 3080 19717 3108
rect 19668 3068 19674 3080
rect 19705 3077 19717 3080
rect 19751 3077 19763 3111
rect 22462 3108 22468 3120
rect 20930 3080 22468 3108
rect 19705 3071 19763 3077
rect 22462 3068 22468 3080
rect 22520 3068 22526 3120
rect 23290 3068 23296 3120
rect 23348 3068 23354 3120
rect 23842 3068 23848 3120
rect 23900 3108 23906 3120
rect 23900 3080 24072 3108
rect 23900 3068 23906 3080
rect 17221 3043 17279 3049
rect 17221 3009 17233 3043
rect 17267 3009 17279 3043
rect 17221 3003 17279 3009
rect 19334 3000 19340 3052
rect 19392 3040 19398 3052
rect 24044 3049 24072 3080
rect 25498 3068 25504 3120
rect 25556 3068 25562 3120
rect 28442 3108 28448 3120
rect 28092 3080 28448 3108
rect 19429 3043 19487 3049
rect 19429 3040 19441 3043
rect 19392 3012 19441 3040
rect 19392 3000 19398 3012
rect 19429 3009 19441 3012
rect 19475 3009 19487 3043
rect 19429 3003 19487 3009
rect 24029 3043 24087 3049
rect 24029 3009 24041 3043
rect 24075 3009 24087 3043
rect 24029 3003 24087 3009
rect 26234 3000 26240 3052
rect 26292 3040 26298 3052
rect 27430 3040 27436 3052
rect 26292 3012 26337 3040
rect 27391 3012 27436 3040
rect 26292 3000 26298 3012
rect 27430 3000 27436 3012
rect 27488 3000 27494 3052
rect 28092 3049 28120 3080
rect 28442 3068 28448 3080
rect 28500 3068 28506 3120
rect 28626 3068 28632 3120
rect 28684 3108 28690 3120
rect 33045 3111 33103 3117
rect 33045 3108 33057 3111
rect 28684 3080 33057 3108
rect 28684 3068 28690 3080
rect 33045 3077 33057 3080
rect 33091 3077 33103 3111
rect 33045 3071 33103 3077
rect 28077 3043 28135 3049
rect 28077 3009 28089 3043
rect 28123 3009 28135 3043
rect 28534 3040 28540 3052
rect 28495 3012 28540 3040
rect 28077 3003 28135 3009
rect 28534 3000 28540 3012
rect 28592 3040 28598 3052
rect 28592 3012 28764 3040
rect 28592 3000 28598 3012
rect 17497 2975 17555 2981
rect 17497 2972 17509 2975
rect 17144 2944 17509 2972
rect 17497 2941 17509 2944
rect 17543 2941 17555 2975
rect 17497 2935 17555 2941
rect 17586 2932 17592 2984
rect 17644 2972 17650 2984
rect 18969 2975 19027 2981
rect 18969 2972 18981 2975
rect 17644 2944 18981 2972
rect 17644 2932 17650 2944
rect 18969 2941 18981 2944
rect 19015 2941 19027 2975
rect 18969 2935 19027 2941
rect 19150 2932 19156 2984
rect 19208 2972 19214 2984
rect 21453 2975 21511 2981
rect 21453 2972 21465 2975
rect 19208 2944 21465 2972
rect 19208 2932 19214 2944
rect 21453 2941 21465 2944
rect 21499 2941 21511 2975
rect 21453 2935 21511 2941
rect 22005 2975 22063 2981
rect 22005 2941 22017 2975
rect 22051 2941 22063 2975
rect 23382 2972 23388 2984
rect 22005 2935 22063 2941
rect 22388 2944 23388 2972
rect 20714 2864 20720 2916
rect 20772 2904 20778 2916
rect 22020 2904 22048 2935
rect 20772 2876 22048 2904
rect 20772 2864 20778 2876
rect 19794 2836 19800 2848
rect 17052 2808 19800 2836
rect 19794 2796 19800 2808
rect 19852 2796 19858 2848
rect 20438 2796 20444 2848
rect 20496 2836 20502 2848
rect 22388 2836 22416 2944
rect 23382 2932 23388 2944
rect 23440 2932 23446 2984
rect 23750 2972 23756 2984
rect 23663 2944 23756 2972
rect 23750 2932 23756 2944
rect 23808 2972 23814 2984
rect 24486 2972 24492 2984
rect 23808 2944 24164 2972
rect 24447 2944 24492 2972
rect 23808 2932 23814 2944
rect 24136 2904 24164 2944
rect 24486 2932 24492 2944
rect 24544 2932 24550 2984
rect 25222 2932 25228 2984
rect 25280 2972 25286 2984
rect 25961 2975 26019 2981
rect 25961 2972 25973 2975
rect 25280 2944 25973 2972
rect 25280 2932 25286 2944
rect 25961 2941 25973 2944
rect 26007 2972 26019 2975
rect 28626 2972 28632 2984
rect 26007 2944 28632 2972
rect 26007 2941 26019 2944
rect 25961 2935 26019 2941
rect 28626 2932 28632 2944
rect 28684 2932 28690 2984
rect 24854 2904 24860 2916
rect 24136 2876 24860 2904
rect 24854 2864 24860 2876
rect 24912 2864 24918 2916
rect 28736 2904 28764 3012
rect 28902 3000 28908 3052
rect 28960 3044 28966 3052
rect 29181 3044 29239 3049
rect 28960 3043 29239 3044
rect 28960 3016 29193 3043
rect 28960 3012 28994 3016
rect 28960 3000 28966 3012
rect 29181 3009 29193 3016
rect 29227 3009 29239 3043
rect 29181 3003 29239 3009
rect 29270 3000 29276 3052
rect 29328 3040 29334 3052
rect 29730 3040 29736 3052
rect 29328 3012 29736 3040
rect 29328 3000 29334 3012
rect 29730 3000 29736 3012
rect 29788 3040 29794 3052
rect 29825 3043 29883 3049
rect 29825 3040 29837 3043
rect 29788 3012 29837 3040
rect 29788 3000 29794 3012
rect 29825 3009 29837 3012
rect 29871 3009 29883 3043
rect 29825 3003 29883 3009
rect 30282 3000 30288 3052
rect 30340 3040 30346 3052
rect 30653 3043 30711 3049
rect 30653 3040 30665 3043
rect 30340 3012 30665 3040
rect 30340 3000 30346 3012
rect 30653 3009 30665 3012
rect 30699 3040 30711 3043
rect 31297 3043 31355 3049
rect 31297 3040 31309 3043
rect 30699 3012 31309 3040
rect 30699 3009 30711 3012
rect 30653 3003 30711 3009
rect 31297 3009 31309 3012
rect 31343 3009 31355 3043
rect 32490 3040 32496 3052
rect 32451 3012 32496 3040
rect 31297 3003 31355 3009
rect 32490 3000 32496 3012
rect 32548 3040 32554 3052
rect 32953 3043 33011 3049
rect 32953 3040 32965 3043
rect 32548 3012 32965 3040
rect 32548 3000 32554 3012
rect 32953 3009 32965 3012
rect 32999 3009 33011 3043
rect 32953 3003 33011 3009
rect 33134 3000 33140 3052
rect 33192 3040 33198 3052
rect 33597 3043 33655 3049
rect 33597 3040 33609 3043
rect 33192 3012 33609 3040
rect 33192 3000 33198 3012
rect 33597 3009 33609 3012
rect 33643 3009 33655 3043
rect 38010 3040 38016 3052
rect 37971 3012 38016 3040
rect 33597 3003 33655 3009
rect 38010 3000 38016 3012
rect 38068 3000 38074 3052
rect 31018 2932 31024 2984
rect 31076 2972 31082 2984
rect 34241 2975 34299 2981
rect 34241 2972 34253 2975
rect 31076 2944 34253 2972
rect 31076 2932 31082 2944
rect 34241 2941 34253 2944
rect 34287 2941 34299 2975
rect 34241 2935 34299 2941
rect 34330 2932 34336 2984
rect 34388 2972 34394 2984
rect 35345 2975 35403 2981
rect 35345 2972 35357 2975
rect 34388 2944 35357 2972
rect 34388 2932 34394 2944
rect 35345 2941 35357 2944
rect 35391 2941 35403 2975
rect 35345 2935 35403 2941
rect 30834 2904 30840 2916
rect 28736 2876 30840 2904
rect 30834 2864 30840 2876
rect 30892 2864 30898 2916
rect 33781 2907 33839 2913
rect 33781 2873 33793 2907
rect 33827 2904 33839 2907
rect 36630 2904 36636 2916
rect 33827 2876 36636 2904
rect 33827 2873 33839 2876
rect 33781 2867 33839 2873
rect 36630 2864 36636 2876
rect 36688 2864 36694 2916
rect 20496 2808 22416 2836
rect 20496 2796 20502 2808
rect 27062 2796 27068 2848
rect 27120 2836 27126 2848
rect 27249 2839 27307 2845
rect 27249 2836 27261 2839
rect 27120 2808 27261 2836
rect 27120 2796 27126 2808
rect 27249 2805 27261 2808
rect 27295 2805 27307 2839
rect 27890 2836 27896 2848
rect 27851 2808 27896 2836
rect 27249 2799 27307 2805
rect 27890 2796 27896 2808
rect 27948 2796 27954 2848
rect 28721 2839 28779 2845
rect 28721 2805 28733 2839
rect 28767 2836 28779 2839
rect 28902 2836 28908 2848
rect 28767 2808 28908 2836
rect 28767 2805 28779 2808
rect 28721 2799 28779 2805
rect 28902 2796 28908 2808
rect 28960 2796 28966 2848
rect 29270 2836 29276 2848
rect 29231 2808 29276 2836
rect 29270 2796 29276 2808
rect 29328 2796 29334 2848
rect 29914 2836 29920 2848
rect 29875 2808 29920 2836
rect 29914 2796 29920 2808
rect 29972 2796 29978 2848
rect 30558 2836 30564 2848
rect 30519 2808 30564 2836
rect 30558 2796 30564 2808
rect 30616 2796 30622 2848
rect 31202 2836 31208 2848
rect 31163 2808 31208 2836
rect 31202 2796 31208 2808
rect 31260 2796 31266 2848
rect 32306 2796 32312 2848
rect 32364 2836 32370 2848
rect 34793 2839 34851 2845
rect 34793 2836 34805 2839
rect 32364 2808 34805 2836
rect 32364 2796 32370 2808
rect 34793 2805 34805 2808
rect 34839 2805 34851 2839
rect 34793 2799 34851 2805
rect 35434 2796 35440 2848
rect 35492 2836 35498 2848
rect 35897 2839 35955 2845
rect 35897 2836 35909 2839
rect 35492 2808 35909 2836
rect 35492 2796 35498 2808
rect 35897 2805 35909 2808
rect 35943 2805 35955 2839
rect 38194 2836 38200 2848
rect 38155 2808 38200 2836
rect 35897 2799 35955 2805
rect 38194 2796 38200 2808
rect 38252 2796 38258 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 2130 2592 2136 2644
rect 2188 2632 2194 2644
rect 3237 2635 3295 2641
rect 3237 2632 3249 2635
rect 2188 2604 3249 2632
rect 2188 2592 2194 2604
rect 3237 2601 3249 2604
rect 3283 2601 3295 2635
rect 3237 2595 3295 2601
rect 7469 2635 7527 2641
rect 7469 2601 7481 2635
rect 7515 2632 7527 2635
rect 8018 2632 8024 2644
rect 7515 2604 8024 2632
rect 7515 2601 7527 2604
rect 7469 2595 7527 2601
rect 8018 2592 8024 2604
rect 8076 2592 8082 2644
rect 10042 2632 10048 2644
rect 10003 2604 10048 2632
rect 10042 2592 10048 2604
rect 10100 2592 10106 2644
rect 11698 2592 11704 2644
rect 11756 2632 11762 2644
rect 11977 2635 12035 2641
rect 11977 2632 11989 2635
rect 11756 2604 11989 2632
rect 11756 2592 11762 2604
rect 11977 2601 11989 2604
rect 12023 2601 12035 2635
rect 11977 2595 12035 2601
rect 13262 2592 13268 2644
rect 13320 2632 13326 2644
rect 14810 2635 14868 2641
rect 14810 2632 14822 2635
rect 13320 2604 14822 2632
rect 13320 2592 13326 2604
rect 14810 2601 14822 2604
rect 14856 2601 14868 2635
rect 22002 2632 22008 2644
rect 14810 2595 14868 2601
rect 18524 2604 22008 2632
rect 14 2524 20 2576
rect 72 2564 78 2576
rect 2409 2567 2467 2573
rect 2409 2564 2421 2567
rect 72 2536 2421 2564
rect 72 2524 78 2536
rect 2409 2533 2421 2536
rect 2455 2533 2467 2567
rect 2409 2527 2467 2533
rect 3326 2524 3332 2576
rect 3384 2524 3390 2576
rect 10778 2524 10784 2576
rect 10836 2564 10842 2576
rect 10873 2567 10931 2573
rect 10873 2564 10885 2567
rect 10836 2536 10885 2564
rect 10836 2524 10842 2536
rect 10873 2533 10885 2536
rect 10919 2533 10931 2567
rect 10873 2527 10931 2533
rect 12342 2524 12348 2576
rect 12400 2564 12406 2576
rect 12400 2536 12480 2564
rect 12400 2524 12406 2536
rect 3344 2496 3372 2524
rect 7190 2496 7196 2508
rect 1872 2468 3372 2496
rect 4908 2468 7196 2496
rect 1872 2437 1900 2468
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2397 1915 2431
rect 1857 2391 1915 2397
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2428 2651 2431
rect 2866 2428 2872 2440
rect 2639 2400 2872 2428
rect 2639 2397 2651 2400
rect 2593 2391 2651 2397
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 4908 2437 4936 2468
rect 7190 2456 7196 2468
rect 7248 2456 7254 2508
rect 12452 2496 12480 2536
rect 13725 2499 13783 2505
rect 13725 2496 13737 2499
rect 12452 2468 13737 2496
rect 13725 2465 13737 2468
rect 13771 2496 13783 2499
rect 14550 2496 14556 2508
rect 13771 2468 14556 2496
rect 13771 2465 13783 2468
rect 13725 2459 13783 2465
rect 14550 2456 14556 2468
rect 14608 2496 14614 2508
rect 17126 2496 17132 2508
rect 14608 2468 17132 2496
rect 14608 2456 14614 2468
rect 17126 2456 17132 2468
rect 17184 2456 17190 2508
rect 3329 2431 3387 2437
rect 3329 2428 3341 2431
rect 3292 2400 3341 2428
rect 3292 2388 3298 2400
rect 3329 2397 3341 2400
rect 3375 2428 3387 2431
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3375 2400 3985 2428
rect 3375 2397 3387 2400
rect 3329 2391 3387 2397
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 6825 2431 6883 2437
rect 6825 2397 6837 2431
rect 6871 2428 6883 2431
rect 8202 2428 8208 2440
rect 6871 2400 8208 2428
rect 6871 2397 6883 2400
rect 6825 2391 6883 2397
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 9858 2428 9864 2440
rect 9819 2400 9864 2428
rect 9858 2388 9864 2400
rect 9916 2388 9922 2440
rect 11057 2431 11115 2437
rect 11057 2397 11069 2431
rect 11103 2428 11115 2431
rect 11146 2428 11152 2440
rect 11103 2400 11152 2428
rect 11103 2397 11115 2400
rect 11057 2391 11115 2397
rect 11146 2388 11152 2400
rect 11204 2388 11210 2440
rect 12342 2388 12348 2440
rect 12400 2388 12406 2440
rect 18524 2414 18552 2604
rect 22002 2592 22008 2604
rect 22060 2592 22066 2644
rect 27985 2635 28043 2641
rect 27985 2601 27997 2635
rect 28031 2632 28043 2635
rect 29546 2632 29552 2644
rect 28031 2604 29552 2632
rect 28031 2601 28043 2604
rect 27985 2595 28043 2601
rect 29546 2592 29552 2604
rect 29604 2592 29610 2644
rect 31294 2592 31300 2644
rect 31352 2632 31358 2644
rect 32953 2635 33011 2641
rect 32953 2632 32965 2635
rect 31352 2604 32965 2632
rect 31352 2592 31358 2604
rect 32953 2601 32965 2604
rect 32999 2601 33011 2635
rect 32953 2595 33011 2601
rect 33594 2592 33600 2644
rect 33652 2632 33658 2644
rect 34149 2635 34207 2641
rect 34149 2632 34161 2635
rect 33652 2604 34161 2632
rect 33652 2592 33658 2604
rect 34149 2601 34161 2604
rect 34195 2601 34207 2635
rect 34149 2595 34207 2601
rect 23474 2524 23480 2576
rect 23532 2564 23538 2576
rect 24581 2567 24639 2573
rect 24581 2564 24593 2567
rect 23532 2536 24593 2564
rect 23532 2524 23538 2536
rect 24581 2533 24593 2536
rect 24627 2533 24639 2567
rect 24581 2527 24639 2533
rect 26510 2524 26516 2576
rect 26568 2564 26574 2576
rect 29270 2564 29276 2576
rect 26568 2536 29276 2564
rect 26568 2524 26574 2536
rect 29270 2524 29276 2536
rect 29328 2524 29334 2576
rect 30926 2524 30932 2576
rect 30984 2564 30990 2576
rect 35621 2567 35679 2573
rect 35621 2564 35633 2567
rect 30984 2536 35633 2564
rect 30984 2524 30990 2536
rect 35621 2533 35633 2536
rect 35667 2533 35679 2567
rect 35621 2527 35679 2533
rect 18598 2456 18604 2508
rect 18656 2496 18662 2508
rect 19705 2499 19763 2505
rect 19705 2496 19717 2499
rect 18656 2468 19717 2496
rect 18656 2456 18662 2468
rect 19705 2465 19717 2468
rect 19751 2465 19763 2499
rect 19705 2459 19763 2465
rect 22281 2499 22339 2505
rect 22281 2465 22293 2499
rect 22327 2496 22339 2499
rect 24394 2496 24400 2508
rect 22327 2468 24400 2496
rect 22327 2465 22339 2468
rect 22281 2459 22339 2465
rect 24394 2456 24400 2468
rect 24452 2456 24458 2508
rect 25038 2496 25044 2508
rect 24504 2468 25044 2496
rect 19426 2428 19432 2440
rect 19339 2400 19432 2428
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 22005 2431 22063 2437
rect 22005 2397 22017 2431
rect 22051 2397 22063 2431
rect 24504 2428 24532 2468
rect 25038 2456 25044 2468
rect 25096 2456 25102 2508
rect 26326 2496 26332 2508
rect 26287 2468 26332 2496
rect 26326 2456 26332 2468
rect 26384 2456 26390 2508
rect 29822 2496 29828 2508
rect 29783 2468 29828 2496
rect 29822 2456 29828 2468
rect 29880 2456 29886 2508
rect 34054 2496 34060 2508
rect 29932 2468 31248 2496
rect 23414 2400 24532 2428
rect 27433 2431 27491 2437
rect 22005 2391 22063 2397
rect 27433 2397 27445 2431
rect 27479 2428 27491 2431
rect 27890 2428 27896 2440
rect 27479 2400 27896 2428
rect 27479 2397 27491 2400
rect 27433 2391 27491 2397
rect 5997 2363 6055 2369
rect 5997 2329 6009 2363
rect 6043 2360 6055 2363
rect 8386 2360 8392 2372
rect 6043 2332 8392 2360
rect 6043 2329 6055 2332
rect 5997 2323 6055 2329
rect 8386 2320 8392 2332
rect 8444 2360 8450 2372
rect 9217 2363 9275 2369
rect 9217 2360 9229 2363
rect 8444 2332 9229 2360
rect 8444 2320 8450 2332
rect 9217 2329 9229 2332
rect 9263 2329 9275 2363
rect 9217 2323 9275 2329
rect 13449 2363 13507 2369
rect 13449 2329 13461 2363
rect 13495 2360 13507 2363
rect 13538 2360 13544 2372
rect 13495 2332 13544 2360
rect 13495 2329 13507 2332
rect 13449 2323 13507 2329
rect 13538 2320 13544 2332
rect 13596 2320 13602 2372
rect 17310 2360 17316 2372
rect 16054 2332 17316 2360
rect 17310 2320 17316 2332
rect 17368 2320 17374 2372
rect 17405 2363 17463 2369
rect 17405 2329 17417 2363
rect 17451 2360 17463 2363
rect 17678 2360 17684 2372
rect 17451 2332 17684 2360
rect 17451 2329 17463 2332
rect 17405 2323 17463 2329
rect 17678 2320 17684 2332
rect 17736 2320 17742 2372
rect 19444 2360 19472 2388
rect 19978 2360 19984 2372
rect 19444 2332 19984 2360
rect 19978 2320 19984 2332
rect 20036 2320 20042 2372
rect 21358 2360 21364 2372
rect 20930 2332 21364 2360
rect 21358 2320 21364 2332
rect 21416 2320 21422 2372
rect 21450 2320 21456 2372
rect 21508 2360 21514 2372
rect 21508 2332 21553 2360
rect 21508 2320 21514 2332
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 1360 2264 1685 2292
rect 1360 2252 1366 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 4522 2252 4528 2304
rect 4580 2292 4586 2304
rect 4709 2295 4767 2301
rect 4709 2292 4721 2295
rect 4580 2264 4721 2292
rect 4580 2252 4586 2264
rect 4709 2261 4721 2264
rect 4755 2261 4767 2295
rect 4709 2255 4767 2261
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6641 2295 6699 2301
rect 6641 2292 6653 2295
rect 6512 2264 6653 2292
rect 6512 2252 6518 2264
rect 6641 2261 6653 2264
rect 6687 2261 6699 2295
rect 8570 2292 8576 2304
rect 8531 2264 8576 2292
rect 6641 2255 6699 2261
rect 8570 2252 8576 2264
rect 8628 2252 8634 2304
rect 9306 2292 9312 2304
rect 9267 2264 9312 2292
rect 9306 2252 9312 2264
rect 9364 2252 9370 2304
rect 11330 2252 11336 2304
rect 11388 2292 11394 2304
rect 16301 2295 16359 2301
rect 16301 2292 16313 2295
rect 11388 2264 16313 2292
rect 11388 2252 11394 2264
rect 16301 2261 16313 2264
rect 16347 2292 16359 2295
rect 18414 2292 18420 2304
rect 16347 2264 18420 2292
rect 16347 2261 16359 2264
rect 16301 2255 16359 2261
rect 18414 2252 18420 2264
rect 18472 2252 18478 2304
rect 18877 2295 18935 2301
rect 18877 2261 18889 2295
rect 18923 2292 18935 2295
rect 19886 2292 19892 2304
rect 18923 2264 19892 2292
rect 18923 2261 18935 2264
rect 18877 2255 18935 2261
rect 19886 2252 19892 2264
rect 19944 2252 19950 2304
rect 19996 2292 20024 2320
rect 22020 2292 22048 2391
rect 27890 2388 27896 2400
rect 27948 2388 27954 2440
rect 27982 2388 27988 2440
rect 28040 2428 28046 2440
rect 28810 2428 28816 2440
rect 28040 2400 28816 2428
rect 28040 2388 28046 2400
rect 28810 2388 28816 2400
rect 28868 2388 28874 2440
rect 29730 2428 29736 2440
rect 29691 2400 29736 2428
rect 29730 2388 29736 2400
rect 29788 2388 29794 2440
rect 25590 2320 25596 2372
rect 25648 2320 25654 2372
rect 26053 2363 26111 2369
rect 26053 2329 26065 2363
rect 26099 2360 26111 2363
rect 26418 2360 26424 2372
rect 26099 2332 26424 2360
rect 26099 2329 26111 2332
rect 26053 2323 26111 2329
rect 26418 2320 26424 2332
rect 26476 2320 26482 2372
rect 28074 2360 28080 2372
rect 28035 2332 28080 2360
rect 28074 2320 28080 2332
rect 28132 2360 28138 2372
rect 29932 2360 29960 2468
rect 30653 2431 30711 2437
rect 30653 2397 30665 2431
rect 30699 2428 30711 2431
rect 30699 2400 31156 2428
rect 30699 2397 30711 2400
rect 30653 2391 30711 2397
rect 28132 2332 29960 2360
rect 28132 2320 28138 2332
rect 23750 2292 23756 2304
rect 19996 2264 22048 2292
rect 23711 2264 23756 2292
rect 23750 2252 23756 2264
rect 23808 2252 23814 2304
rect 23842 2252 23848 2304
rect 23900 2292 23906 2304
rect 27249 2295 27307 2301
rect 27249 2292 27261 2295
rect 23900 2264 27261 2292
rect 23900 2252 23906 2264
rect 27249 2261 27261 2264
rect 27295 2261 27307 2295
rect 28718 2292 28724 2304
rect 28679 2264 28724 2292
rect 27249 2255 27307 2261
rect 28718 2252 28724 2264
rect 28776 2252 28782 2304
rect 30282 2252 30288 2304
rect 30340 2292 30346 2304
rect 31128 2301 31156 2400
rect 31220 2360 31248 2468
rect 31726 2468 34060 2496
rect 31294 2388 31300 2440
rect 31352 2428 31358 2440
rect 31352 2400 31397 2428
rect 31352 2388 31358 2400
rect 31726 2360 31754 2468
rect 34054 2456 34060 2468
rect 34112 2456 34118 2508
rect 32306 2428 32312 2440
rect 32267 2400 32312 2428
rect 32306 2388 32312 2400
rect 32364 2388 32370 2440
rect 33137 2431 33195 2437
rect 33137 2397 33149 2431
rect 33183 2428 33195 2431
rect 34330 2428 34336 2440
rect 33183 2400 34336 2428
rect 33183 2397 33195 2400
rect 33137 2391 33195 2397
rect 31220 2332 31754 2360
rect 32214 2320 32220 2372
rect 32272 2360 32278 2372
rect 33152 2360 33180 2391
rect 34330 2388 34336 2400
rect 34388 2388 34394 2440
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34848 2400 34897 2428
rect 34848 2388 34854 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 36630 2428 36636 2440
rect 36591 2400 36636 2428
rect 34885 2391 34943 2397
rect 36630 2388 36636 2400
rect 36688 2388 36694 2440
rect 37458 2428 37464 2440
rect 37419 2400 37464 2428
rect 37458 2388 37464 2400
rect 37516 2388 37522 2440
rect 32272 2332 33180 2360
rect 32272 2320 32278 2332
rect 35434 2320 35440 2372
rect 35492 2360 35498 2372
rect 35805 2363 35863 2369
rect 35805 2360 35817 2363
rect 35492 2332 35817 2360
rect 35492 2320 35498 2332
rect 35805 2329 35817 2332
rect 35851 2329 35863 2363
rect 35805 2323 35863 2329
rect 30469 2295 30527 2301
rect 30469 2292 30481 2295
rect 30340 2264 30481 2292
rect 30340 2252 30346 2264
rect 30469 2261 30481 2264
rect 30515 2261 30527 2295
rect 30469 2255 30527 2261
rect 31113 2295 31171 2301
rect 31113 2261 31125 2295
rect 31159 2261 31171 2295
rect 31113 2255 31171 2261
rect 32493 2295 32551 2301
rect 32493 2261 32505 2295
rect 32539 2292 32551 2295
rect 33134 2292 33140 2304
rect 32539 2264 33140 2292
rect 32539 2261 32551 2264
rect 32493 2255 32551 2261
rect 33134 2252 33140 2264
rect 33192 2252 33198 2304
rect 33594 2292 33600 2304
rect 33555 2264 33600 2292
rect 33594 2252 33600 2264
rect 33652 2252 33658 2304
rect 34146 2252 34152 2304
rect 34204 2292 34210 2304
rect 35069 2295 35127 2301
rect 35069 2292 35081 2295
rect 34204 2264 35081 2292
rect 34204 2252 34210 2264
rect 35069 2261 35081 2264
rect 35115 2261 35127 2295
rect 35069 2255 35127 2261
rect 36817 2295 36875 2301
rect 36817 2261 36829 2295
rect 36863 2292 36875 2295
rect 37182 2292 37188 2304
rect 36863 2264 37188 2292
rect 36863 2261 36875 2264
rect 36817 2255 36875 2261
rect 37182 2252 37188 2264
rect 37240 2252 37246 2304
rect 37366 2252 37372 2304
rect 37424 2292 37430 2304
rect 37645 2295 37703 2301
rect 37645 2292 37657 2295
rect 37424 2264 37657 2292
rect 37424 2252 37430 2264
rect 37645 2261 37657 2264
rect 37691 2261 37703 2295
rect 37645 2255 37703 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 17310 2048 17316 2100
rect 17368 2088 17374 2100
rect 17368 2060 22140 2088
rect 17368 2048 17374 2060
rect 8570 1980 8576 2032
rect 8628 2020 8634 2032
rect 18598 2020 18604 2032
rect 8628 1992 18604 2020
rect 8628 1980 8634 1992
rect 18598 1980 18604 1992
rect 18656 1980 18662 2032
rect 18874 1980 18880 2032
rect 18932 2020 18938 2032
rect 21450 2020 21456 2032
rect 18932 1992 21456 2020
rect 18932 1980 18938 1992
rect 21450 1980 21456 1992
rect 21508 1980 21514 2032
rect 22112 2020 22140 2060
rect 22186 2048 22192 2100
rect 22244 2088 22250 2100
rect 28718 2088 28724 2100
rect 22244 2060 28724 2088
rect 22244 2048 22250 2060
rect 28718 2048 28724 2060
rect 28776 2048 28782 2100
rect 28902 2048 28908 2100
rect 28960 2088 28966 2100
rect 37458 2088 37464 2100
rect 28960 2060 37464 2088
rect 28960 2048 28966 2060
rect 37458 2048 37464 2060
rect 37516 2048 37522 2100
rect 31202 2020 31208 2032
rect 22112 1992 31208 2020
rect 31202 1980 31208 1992
rect 31260 1980 31266 2032
rect 16206 1912 16212 1964
rect 16264 1952 16270 1964
rect 31754 1952 31760 1964
rect 16264 1924 31760 1952
rect 16264 1912 16270 1924
rect 31754 1912 31760 1924
rect 31812 1912 31818 1964
rect 13354 1844 13360 1896
rect 13412 1884 13418 1896
rect 25498 1884 25504 1896
rect 13412 1856 25504 1884
rect 13412 1844 13418 1856
rect 25498 1844 25504 1856
rect 25556 1844 25562 1896
rect 25590 1844 25596 1896
rect 25648 1884 25654 1896
rect 30558 1884 30564 1896
rect 25648 1856 30564 1884
rect 25648 1844 25654 1856
rect 30558 1844 30564 1856
rect 30616 1844 30622 1896
rect 21358 1776 21364 1828
rect 21416 1816 21422 1828
rect 33594 1816 33600 1828
rect 21416 1788 33600 1816
rect 21416 1776 21422 1788
rect 33594 1776 33600 1788
rect 33652 1776 33658 1828
rect 25130 1708 25136 1760
rect 25188 1748 25194 1760
rect 28074 1748 28080 1760
rect 25188 1720 28080 1748
rect 25188 1708 25194 1720
rect 28074 1708 28080 1720
rect 28132 1708 28138 1760
rect 28994 1708 29000 1760
rect 29052 1748 29058 1760
rect 32306 1748 32312 1760
rect 29052 1720 32312 1748
rect 29052 1708 29058 1720
rect 32306 1708 32312 1720
rect 32364 1708 32370 1760
rect 9306 1640 9312 1692
rect 9364 1680 9370 1692
rect 26786 1680 26792 1692
rect 9364 1652 26792 1680
rect 9364 1640 9370 1652
rect 26786 1640 26792 1652
rect 26844 1640 26850 1692
rect 25498 1572 25504 1624
rect 25556 1612 25562 1624
rect 30466 1612 30472 1624
rect 25556 1584 30472 1612
rect 25556 1572 25562 1584
rect 30466 1572 30472 1584
rect 30524 1572 30530 1624
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 18052 37408 18104 37460
rect 2320 37204 2372 37256
rect 5448 37204 5500 37256
rect 7288 37204 7340 37256
rect 7748 37204 7800 37256
rect 6736 37136 6788 37188
rect 12072 37204 12124 37256
rect 14832 37272 14884 37324
rect 16672 37272 16724 37324
rect 16764 37272 16816 37324
rect 18144 37315 18196 37324
rect 18144 37281 18153 37315
rect 18153 37281 18187 37315
rect 18187 37281 18196 37315
rect 18144 37272 18196 37281
rect 21916 37272 21968 37324
rect 35440 37272 35492 37324
rect 38292 37315 38344 37324
rect 38292 37281 38301 37315
rect 38301 37281 38335 37315
rect 38335 37281 38344 37315
rect 38292 37272 38344 37281
rect 13268 37247 13320 37256
rect 13268 37213 13277 37247
rect 13277 37213 13311 37247
rect 13311 37213 13320 37247
rect 13268 37204 13320 37213
rect 13360 37204 13412 37256
rect 18052 37204 18104 37256
rect 20076 37247 20128 37256
rect 20076 37213 20085 37247
rect 20085 37213 20119 37247
rect 20119 37213 20128 37247
rect 20076 37204 20128 37213
rect 20536 37204 20588 37256
rect 23020 37204 23072 37256
rect 23296 37247 23348 37256
rect 23296 37213 23305 37247
rect 23305 37213 23339 37247
rect 23339 37213 23348 37247
rect 23296 37204 23348 37213
rect 13176 37136 13228 37188
rect 20720 37136 20772 37188
rect 25872 37204 25924 37256
rect 27436 37204 27488 37256
rect 30472 37204 30524 37256
rect 30840 37204 30892 37256
rect 33600 37247 33652 37256
rect 33600 37213 33609 37247
rect 33609 37213 33643 37247
rect 33643 37213 33652 37247
rect 33600 37204 33652 37213
rect 35808 37247 35860 37256
rect 35808 37213 35817 37247
rect 35817 37213 35851 37247
rect 35851 37213 35860 37247
rect 35808 37204 35860 37213
rect 37832 37204 37884 37256
rect 1308 37068 1360 37120
rect 2780 37111 2832 37120
rect 2780 37077 2789 37111
rect 2789 37077 2823 37111
rect 2823 37077 2832 37111
rect 2780 37068 2832 37077
rect 4620 37068 4672 37120
rect 5448 37111 5500 37120
rect 5448 37077 5457 37111
rect 5457 37077 5491 37111
rect 5491 37077 5500 37111
rect 5448 37068 5500 37077
rect 6460 37068 6512 37120
rect 8024 37111 8076 37120
rect 8024 37077 8033 37111
rect 8033 37077 8067 37111
rect 8067 37077 8076 37111
rect 8024 37068 8076 37077
rect 9680 37068 9732 37120
rect 11612 37068 11664 37120
rect 12900 37068 12952 37120
rect 19984 37068 20036 37120
rect 23204 37068 23256 37120
rect 25136 37068 25188 37120
rect 27068 37068 27120 37120
rect 28356 37068 28408 37120
rect 30380 37068 30432 37120
rect 32220 37068 32272 37120
rect 33508 37068 33560 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 5448 36864 5500 36916
rect 22100 36864 22152 36916
rect 23296 36864 23348 36916
rect 33600 36864 33652 36916
rect 37372 36864 37424 36916
rect 2872 36796 2924 36848
rect 2964 36728 3016 36780
rect 13360 36728 13412 36780
rect 22284 36728 22336 36780
rect 22744 36728 22796 36780
rect 23020 36728 23072 36780
rect 37740 36771 37792 36780
rect 37740 36737 37749 36771
rect 37749 36737 37783 36771
rect 37783 36737 37792 36771
rect 37740 36728 37792 36737
rect 37924 36660 37976 36712
rect 16304 36592 16356 36644
rect 2504 36567 2556 36576
rect 2504 36533 2513 36567
rect 2513 36533 2547 36567
rect 2547 36533 2556 36567
rect 2504 36524 2556 36533
rect 7288 36524 7340 36576
rect 22744 36567 22796 36576
rect 22744 36533 22753 36567
rect 22753 36533 22787 36567
rect 22787 36533 22796 36567
rect 22744 36524 22796 36533
rect 38016 36524 38068 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2872 36320 2924 36372
rect 22744 36320 22796 36372
rect 35808 36320 35860 36372
rect 37188 36320 37240 36372
rect 38660 36320 38712 36372
rect 1860 36159 1912 36168
rect 1860 36125 1869 36159
rect 1869 36125 1903 36159
rect 1903 36125 1912 36159
rect 1860 36116 1912 36125
rect 38016 36159 38068 36168
rect 38016 36125 38025 36159
rect 38025 36125 38059 36159
rect 38059 36125 38068 36159
rect 38016 36116 38068 36125
rect 1676 36023 1728 36032
rect 1676 35989 1685 36023
rect 1685 35989 1719 36023
rect 1719 35989 1728 36023
rect 1676 35980 1728 35989
rect 36728 36023 36780 36032
rect 36728 35989 36737 36023
rect 36737 35989 36771 36023
rect 36771 35989 36780 36023
rect 36728 35980 36780 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 1860 35776 1912 35828
rect 37924 35572 37976 35624
rect 38292 35615 38344 35624
rect 38292 35581 38301 35615
rect 38301 35581 38335 35615
rect 38335 35581 38344 35615
rect 38292 35572 38344 35581
rect 3424 35436 3476 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 20720 35232 20772 35284
rect 30472 35232 30524 35284
rect 38292 35275 38344 35284
rect 38292 35241 38301 35275
rect 38301 35241 38335 35275
rect 38335 35241 38344 35275
rect 38292 35232 38344 35241
rect 19984 35028 20036 35080
rect 29644 35028 29696 35080
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 2228 34484 2280 34536
rect 1676 34391 1728 34400
rect 1676 34357 1685 34391
rect 1685 34357 1719 34391
rect 1719 34357 1728 34391
rect 1676 34348 1728 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 6736 34144 6788 34196
rect 7104 33983 7156 33992
rect 7104 33949 7113 33983
rect 7113 33949 7147 33983
rect 7147 33949 7156 33983
rect 7104 33940 7156 33949
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 12716 33464 12768 33516
rect 38200 33371 38252 33380
rect 38200 33337 38209 33371
rect 38209 33337 38243 33371
rect 38243 33337 38252 33371
rect 38200 33328 38252 33337
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 1584 32376 1636 32428
rect 12992 32172 13044 32224
rect 19984 32376 20036 32428
rect 29644 32376 29696 32428
rect 38292 32351 38344 32360
rect 38292 32317 38301 32351
rect 38301 32317 38335 32351
rect 38335 32317 38344 32351
rect 38292 32308 38344 32317
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 1584 32011 1636 32020
rect 1584 31977 1593 32011
rect 1593 31977 1627 32011
rect 1627 31977 1636 32011
rect 1584 31968 1636 31977
rect 38292 32011 38344 32020
rect 38292 31977 38301 32011
rect 38301 31977 38335 32011
rect 38335 31977 38344 32011
rect 38292 31968 38344 31977
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 27436 30923 27488 30932
rect 27436 30889 27445 30923
rect 27445 30889 27479 30923
rect 27479 30889 27488 30923
rect 27436 30880 27488 30889
rect 30840 30923 30892 30932
rect 30840 30889 30849 30923
rect 30849 30889 30883 30923
rect 30883 30889 30892 30923
rect 30840 30880 30892 30889
rect 1676 30651 1728 30660
rect 1676 30617 1685 30651
rect 1685 30617 1719 30651
rect 1719 30617 1728 30651
rect 1676 30608 1728 30617
rect 1768 30583 1820 30592
rect 1768 30549 1777 30583
rect 1777 30549 1811 30583
rect 1811 30549 1820 30583
rect 1768 30540 1820 30549
rect 30564 30676 30616 30728
rect 29276 30540 29328 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 1676 30379 1728 30388
rect 1676 30345 1685 30379
rect 1685 30345 1719 30379
rect 1719 30345 1728 30379
rect 1676 30336 1728 30345
rect 14740 30200 14792 30252
rect 38016 30243 38068 30252
rect 38016 30209 38025 30243
rect 38025 30209 38059 30243
rect 38059 30209 38068 30243
rect 38016 30200 38068 30209
rect 14740 30039 14792 30048
rect 14740 30005 14749 30039
rect 14749 30005 14783 30039
rect 14783 30005 14792 30039
rect 14740 29996 14792 30005
rect 36728 29996 36780 30048
rect 38200 30039 38252 30048
rect 38200 30005 38209 30039
rect 38209 30005 38243 30039
rect 38243 30005 38252 30039
rect 38200 29996 38252 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 38016 29835 38068 29844
rect 38016 29801 38025 29835
rect 38025 29801 38059 29835
rect 38059 29801 38068 29835
rect 38016 29792 38068 29801
rect 37832 29631 37884 29640
rect 37832 29597 37841 29631
rect 37841 29597 37875 29631
rect 37875 29597 37884 29631
rect 37832 29588 37884 29597
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 37832 29248 37884 29300
rect 38108 29291 38160 29300
rect 38108 29257 38117 29291
rect 38117 29257 38151 29291
rect 38151 29257 38160 29291
rect 38108 29248 38160 29257
rect 20536 29155 20588 29164
rect 20536 29121 20545 29155
rect 20545 29121 20579 29155
rect 20579 29121 20588 29155
rect 20536 29112 20588 29121
rect 1584 29087 1636 29096
rect 1584 29053 1593 29087
rect 1593 29053 1627 29087
rect 1627 29053 1636 29087
rect 1584 29044 1636 29053
rect 14740 29044 14792 29096
rect 20260 28976 20312 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 22284 28747 22336 28756
rect 22284 28713 22293 28747
rect 22293 28713 22327 28747
rect 22327 28713 22336 28747
rect 22284 28704 22336 28713
rect 1584 28679 1636 28688
rect 1584 28645 1593 28679
rect 1593 28645 1627 28679
rect 1627 28645 1636 28679
rect 1584 28636 1636 28645
rect 13360 28500 13412 28552
rect 22284 28500 22336 28552
rect 14280 28364 14332 28416
rect 22652 28364 22704 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 13176 28160 13228 28212
rect 16488 28024 16540 28076
rect 38200 27931 38252 27940
rect 38200 27897 38209 27931
rect 38209 27897 38243 27931
rect 38243 27897 38252 27931
rect 38200 27888 38252 27897
rect 17592 27820 17644 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 22100 27047 22152 27056
rect 22100 27013 22109 27047
rect 22109 27013 22143 27047
rect 22143 27013 22152 27047
rect 22100 27004 22152 27013
rect 6552 26936 6604 26988
rect 1676 26775 1728 26784
rect 1676 26741 1685 26775
rect 1685 26741 1719 26775
rect 1719 26741 1728 26775
rect 1676 26732 1728 26741
rect 37924 26936 37976 26988
rect 38016 26911 38068 26920
rect 38016 26877 38025 26911
rect 38025 26877 38059 26911
rect 38059 26877 38068 26911
rect 38016 26868 38068 26877
rect 38292 26911 38344 26920
rect 38292 26877 38301 26911
rect 38301 26877 38335 26911
rect 38335 26877 38344 26911
rect 38292 26868 38344 26877
rect 23388 26732 23440 26784
rect 26424 26732 26476 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 23388 26528 23440 26580
rect 38016 26528 38068 26580
rect 38292 26571 38344 26580
rect 38292 26537 38301 26571
rect 38301 26537 38335 26571
rect 38335 26537 38344 26571
rect 38292 26528 38344 26537
rect 16488 26503 16540 26512
rect 16488 26469 16497 26503
rect 16497 26469 16531 26503
rect 16531 26469 16540 26503
rect 16488 26460 16540 26469
rect 16304 26367 16356 26376
rect 16304 26333 16313 26367
rect 16313 26333 16347 26367
rect 16347 26333 16356 26367
rect 16304 26324 16356 26333
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 13268 25984 13320 26036
rect 18236 25848 18288 25900
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 12992 25483 13044 25492
rect 12992 25449 13001 25483
rect 13001 25449 13035 25483
rect 13035 25449 13044 25483
rect 12992 25440 13044 25449
rect 1584 25279 1636 25288
rect 1584 25245 1593 25279
rect 1593 25245 1627 25279
rect 1627 25245 1636 25279
rect 1584 25236 1636 25245
rect 2044 25236 2096 25288
rect 12992 25236 13044 25288
rect 16304 25236 16356 25288
rect 29644 25440 29696 25492
rect 16948 25168 17000 25220
rect 12900 25100 12952 25152
rect 25228 25100 25280 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 1584 24939 1636 24948
rect 1584 24905 1593 24939
rect 1593 24905 1627 24939
rect 1627 24905 1636 24939
rect 1584 24896 1636 24905
rect 38016 24803 38068 24812
rect 38016 24769 38025 24803
rect 38025 24769 38059 24803
rect 38059 24769 38068 24803
rect 38016 24760 38068 24769
rect 38200 24599 38252 24608
rect 38200 24565 38209 24599
rect 38209 24565 38243 24599
rect 38243 24565 38252 24599
rect 38200 24556 38252 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 38108 24352 38160 24404
rect 7104 24080 7156 24132
rect 17776 24080 17828 24132
rect 24124 24080 24176 24132
rect 30564 24080 30616 24132
rect 24860 24012 24912 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1860 23715 1912 23724
rect 1860 23681 1869 23715
rect 1869 23681 1903 23715
rect 1903 23681 1912 23715
rect 1860 23672 1912 23681
rect 1676 23511 1728 23520
rect 1676 23477 1685 23511
rect 1685 23477 1719 23511
rect 1719 23477 1728 23511
rect 1676 23468 1728 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 14832 22627 14884 22636
rect 14832 22593 14841 22627
rect 14841 22593 14875 22627
rect 14875 22593 14884 22627
rect 14832 22584 14884 22593
rect 38200 22627 38252 22636
rect 38200 22593 38209 22627
rect 38209 22593 38243 22627
rect 38243 22593 38252 22627
rect 38200 22584 38252 22593
rect 37924 22448 37976 22500
rect 14372 22380 14424 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 6552 21675 6604 21684
rect 6552 21641 6561 21675
rect 6561 21641 6595 21675
rect 6595 21641 6604 21675
rect 6552 21632 6604 21641
rect 19984 21675 20036 21684
rect 19984 21641 19993 21675
rect 19993 21641 20027 21675
rect 20027 21641 20036 21675
rect 19984 21632 20036 21641
rect 25872 21675 25924 21684
rect 25872 21641 25881 21675
rect 25881 21641 25915 21675
rect 25915 21641 25924 21675
rect 25872 21632 25924 21641
rect 1768 21496 1820 21548
rect 1676 21335 1728 21344
rect 1676 21301 1685 21335
rect 1685 21301 1719 21335
rect 1719 21301 1728 21335
rect 1676 21292 1728 21301
rect 17776 21496 17828 21548
rect 28632 21496 28684 21548
rect 37464 21496 37516 21548
rect 10048 21292 10100 21344
rect 37464 21335 37516 21344
rect 37464 21301 37473 21335
rect 37473 21301 37507 21335
rect 37507 21301 37516 21335
rect 37464 21292 37516 21301
rect 38200 21335 38252 21344
rect 38200 21301 38209 21335
rect 38209 21301 38243 21335
rect 38243 21301 38252 21335
rect 38200 21292 38252 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1768 21131 1820 21140
rect 1768 21097 1777 21131
rect 1777 21097 1811 21131
rect 1811 21097 1820 21131
rect 1768 21088 1820 21097
rect 2044 20884 2096 20936
rect 19432 20791 19484 20800
rect 19432 20757 19441 20791
rect 19441 20757 19475 20791
rect 19475 20757 19484 20791
rect 19432 20748 19484 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 19340 20519 19392 20528
rect 19340 20485 19349 20519
rect 19349 20485 19383 20519
rect 19383 20485 19392 20519
rect 19340 20476 19392 20485
rect 19432 20519 19484 20528
rect 19432 20485 19441 20519
rect 19441 20485 19475 20519
rect 19475 20485 19484 20519
rect 19432 20476 19484 20485
rect 19156 20383 19208 20392
rect 19156 20349 19165 20383
rect 19165 20349 19199 20383
rect 19199 20349 19208 20383
rect 19156 20340 19208 20349
rect 19616 20204 19668 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2320 20043 2372 20052
rect 2320 20009 2329 20043
rect 2329 20009 2363 20043
rect 2363 20009 2372 20043
rect 2320 20000 2372 20009
rect 19340 20000 19392 20052
rect 23388 20000 23440 20052
rect 1952 19864 2004 19916
rect 2596 19796 2648 19848
rect 4620 19728 4672 19780
rect 1676 19703 1728 19712
rect 1676 19669 1685 19703
rect 1685 19669 1719 19703
rect 1719 19669 1728 19703
rect 1676 19660 1728 19669
rect 16120 19660 16172 19712
rect 19616 19839 19668 19848
rect 19616 19805 19625 19839
rect 19625 19805 19659 19839
rect 19659 19805 19668 19839
rect 19616 19796 19668 19805
rect 22100 19796 22152 19848
rect 23388 19796 23440 19848
rect 19984 19728 20036 19780
rect 20076 19660 20128 19712
rect 23112 19703 23164 19712
rect 23112 19669 23121 19703
rect 23121 19669 23155 19703
rect 23155 19669 23164 19703
rect 23112 19660 23164 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 1860 19456 1912 19508
rect 2504 19456 2556 19508
rect 2044 19388 2096 19440
rect 12256 19456 12308 19508
rect 15476 19456 15528 19508
rect 2136 19363 2188 19372
rect 2136 19329 2145 19363
rect 2145 19329 2179 19363
rect 2179 19329 2188 19363
rect 2136 19320 2188 19329
rect 12256 19320 12308 19372
rect 9680 19116 9732 19168
rect 11520 19116 11572 19168
rect 20352 19363 20404 19372
rect 12716 19252 12768 19304
rect 20352 19329 20361 19363
rect 20361 19329 20395 19363
rect 20395 19329 20404 19363
rect 20352 19320 20404 19329
rect 36636 19320 36688 19372
rect 24492 19252 24544 19304
rect 19892 19184 19944 19236
rect 21088 19184 21140 19236
rect 24400 19184 24452 19236
rect 20168 19116 20220 19168
rect 23020 19159 23072 19168
rect 23020 19125 23029 19159
rect 23029 19125 23063 19159
rect 23063 19125 23072 19159
rect 23020 19116 23072 19125
rect 23756 19116 23808 19168
rect 38200 19159 38252 19168
rect 38200 19125 38209 19159
rect 38209 19125 38243 19159
rect 38243 19125 38252 19159
rect 38200 19116 38252 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 18236 18955 18288 18964
rect 18236 18921 18245 18955
rect 18245 18921 18279 18955
rect 18279 18921 18288 18955
rect 18236 18912 18288 18921
rect 18512 18912 18564 18964
rect 17132 18844 17184 18896
rect 26884 18844 26936 18896
rect 1768 18776 1820 18828
rect 19432 18776 19484 18828
rect 20444 18776 20496 18828
rect 18236 18708 18288 18760
rect 22100 18751 22152 18760
rect 22100 18717 22109 18751
rect 22109 18717 22143 18751
rect 22143 18717 22152 18751
rect 22100 18708 22152 18717
rect 24216 18708 24268 18760
rect 16212 18683 16264 18692
rect 16212 18649 16221 18683
rect 16221 18649 16255 18683
rect 16255 18649 16264 18683
rect 16212 18640 16264 18649
rect 20168 18640 20220 18692
rect 17132 18572 17184 18624
rect 18788 18615 18840 18624
rect 18788 18581 18797 18615
rect 18797 18581 18831 18615
rect 18831 18581 18840 18615
rect 18788 18572 18840 18581
rect 37464 18640 37516 18692
rect 23480 18572 23532 18624
rect 24584 18615 24636 18624
rect 24584 18581 24593 18615
rect 24593 18581 24627 18615
rect 24627 18581 24636 18615
rect 24584 18572 24636 18581
rect 25964 18572 26016 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 1768 18411 1820 18420
rect 1768 18377 1777 18411
rect 1777 18377 1811 18411
rect 1811 18377 1820 18411
rect 1768 18368 1820 18377
rect 4620 18411 4672 18420
rect 4620 18377 4629 18411
rect 4629 18377 4663 18411
rect 4663 18377 4672 18411
rect 4620 18368 4672 18377
rect 20996 18368 21048 18420
rect 20076 18343 20128 18352
rect 20076 18309 20085 18343
rect 20085 18309 20119 18343
rect 20119 18309 20128 18343
rect 20076 18300 20128 18309
rect 1584 18232 1636 18284
rect 16120 18275 16172 18284
rect 16120 18241 16129 18275
rect 16129 18241 16163 18275
rect 16163 18241 16172 18275
rect 16120 18232 16172 18241
rect 24216 18368 24268 18420
rect 26884 18368 26936 18420
rect 37740 18368 37792 18420
rect 22560 18343 22612 18352
rect 22560 18309 22569 18343
rect 22569 18309 22603 18343
rect 22603 18309 22612 18343
rect 22560 18300 22612 18309
rect 22652 18343 22704 18352
rect 22652 18309 22661 18343
rect 22661 18309 22695 18343
rect 22695 18309 22704 18343
rect 22652 18300 22704 18309
rect 23756 18275 23808 18284
rect 23756 18241 23765 18275
rect 23765 18241 23799 18275
rect 23799 18241 23808 18275
rect 23756 18232 23808 18241
rect 24584 18275 24636 18284
rect 24584 18241 24593 18275
rect 24593 18241 24627 18275
rect 24627 18241 24636 18275
rect 24584 18232 24636 18241
rect 16948 18207 17000 18216
rect 16948 18173 16957 18207
rect 16957 18173 16991 18207
rect 16991 18173 17000 18207
rect 16948 18164 17000 18173
rect 19984 18207 20036 18216
rect 19984 18173 19993 18207
rect 19993 18173 20027 18207
rect 20027 18173 20036 18207
rect 19984 18164 20036 18173
rect 23388 18164 23440 18216
rect 17408 18096 17460 18148
rect 19340 18139 19392 18148
rect 19340 18105 19349 18139
rect 19349 18105 19383 18139
rect 19383 18105 19392 18139
rect 19340 18096 19392 18105
rect 20536 18139 20588 18148
rect 20536 18105 20545 18139
rect 20545 18105 20579 18139
rect 20579 18105 20588 18139
rect 20536 18096 20588 18105
rect 8024 18028 8076 18080
rect 11152 18028 11204 18080
rect 18236 18071 18288 18080
rect 18236 18037 18245 18071
rect 18245 18037 18279 18071
rect 18279 18037 18288 18071
rect 18236 18028 18288 18037
rect 19156 18028 19208 18080
rect 25044 18096 25096 18148
rect 21180 18071 21232 18080
rect 21180 18037 21189 18071
rect 21189 18037 21223 18071
rect 21223 18037 21232 18071
rect 21180 18028 21232 18037
rect 22284 18028 22336 18080
rect 23296 18071 23348 18080
rect 23296 18037 23305 18071
rect 23305 18037 23339 18071
rect 23339 18037 23348 18071
rect 23296 18028 23348 18037
rect 24032 18028 24084 18080
rect 25136 18071 25188 18080
rect 25136 18037 25145 18071
rect 25145 18037 25179 18071
rect 25179 18037 25188 18071
rect 25136 18028 25188 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1584 17799 1636 17808
rect 1584 17765 1593 17799
rect 1593 17765 1627 17799
rect 1627 17765 1636 17799
rect 1584 17756 1636 17765
rect 14924 17620 14976 17672
rect 15936 17756 15988 17808
rect 18420 17688 18472 17740
rect 19892 17688 19944 17740
rect 20260 17731 20312 17740
rect 20260 17697 20269 17731
rect 20269 17697 20303 17731
rect 20303 17697 20312 17731
rect 20628 17731 20680 17740
rect 20260 17688 20312 17697
rect 20628 17697 20637 17731
rect 20637 17697 20671 17731
rect 20671 17697 20680 17731
rect 20628 17688 20680 17697
rect 17132 17620 17184 17672
rect 18236 17620 18288 17672
rect 18696 17620 18748 17672
rect 11244 17552 11296 17604
rect 16764 17552 16816 17604
rect 20076 17620 20128 17672
rect 22560 17824 22612 17876
rect 23296 17824 23348 17876
rect 27068 17824 27120 17876
rect 22376 17688 22428 17740
rect 21640 17620 21692 17672
rect 22284 17663 22336 17672
rect 22284 17629 22293 17663
rect 22293 17629 22327 17663
rect 22327 17629 22336 17663
rect 22284 17620 22336 17629
rect 25872 17756 25924 17808
rect 22652 17688 22704 17740
rect 23204 17688 23256 17740
rect 23756 17688 23808 17740
rect 26884 17688 26936 17740
rect 25964 17663 26016 17672
rect 25964 17629 25973 17663
rect 25973 17629 26007 17663
rect 26007 17629 26016 17663
rect 25964 17620 26016 17629
rect 15384 17484 15436 17536
rect 16672 17484 16724 17536
rect 17500 17484 17552 17536
rect 18604 17484 18656 17536
rect 23480 17552 23532 17604
rect 24308 17552 24360 17604
rect 25044 17552 25096 17604
rect 25228 17595 25280 17604
rect 25228 17561 25237 17595
rect 25237 17561 25271 17595
rect 25271 17561 25280 17595
rect 25228 17552 25280 17561
rect 20720 17484 20772 17536
rect 25412 17484 25464 17536
rect 27068 17527 27120 17536
rect 27068 17493 27077 17527
rect 27077 17493 27111 17527
rect 27111 17493 27120 17527
rect 27068 17484 27120 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 12808 17212 12860 17264
rect 16028 17212 16080 17264
rect 16580 17212 16632 17264
rect 14924 17187 14976 17196
rect 14924 17153 14933 17187
rect 14933 17153 14967 17187
rect 14967 17153 14976 17187
rect 14924 17144 14976 17153
rect 15844 17076 15896 17128
rect 15936 17119 15988 17128
rect 15936 17085 15945 17119
rect 15945 17085 15979 17119
rect 15979 17085 15988 17119
rect 15936 17076 15988 17085
rect 19892 17280 19944 17332
rect 20352 17280 20404 17332
rect 20996 17323 21048 17332
rect 20996 17289 21005 17323
rect 21005 17289 21039 17323
rect 21039 17289 21048 17323
rect 20996 17280 21048 17289
rect 18328 17212 18380 17264
rect 16764 17076 16816 17128
rect 18420 17144 18472 17196
rect 18788 17212 18840 17264
rect 19708 17212 19760 17264
rect 21180 17212 21232 17264
rect 21088 17187 21140 17196
rect 21088 17153 21097 17187
rect 21097 17153 21131 17187
rect 21131 17153 21140 17187
rect 21088 17144 21140 17153
rect 27344 17280 27396 17332
rect 25412 17255 25464 17264
rect 25412 17221 25421 17255
rect 25421 17221 25455 17255
rect 25455 17221 25464 17255
rect 25412 17212 25464 17221
rect 15660 17008 15712 17060
rect 16028 17008 16080 17060
rect 19616 17076 19668 17128
rect 19892 17119 19944 17128
rect 19892 17085 19901 17119
rect 19901 17085 19935 17119
rect 19935 17085 19944 17119
rect 19892 17076 19944 17085
rect 17868 17008 17920 17060
rect 19340 17051 19392 17060
rect 19340 17017 19349 17051
rect 19349 17017 19383 17051
rect 19383 17017 19392 17051
rect 19340 17008 19392 17017
rect 21456 17008 21508 17060
rect 24400 17144 24452 17196
rect 22376 17076 22428 17128
rect 22836 17119 22888 17128
rect 22836 17085 22845 17119
rect 22845 17085 22879 17119
rect 22879 17085 22888 17119
rect 22836 17076 22888 17085
rect 23388 17119 23440 17128
rect 23388 17085 23397 17119
rect 23397 17085 23431 17119
rect 23431 17085 23440 17119
rect 23388 17076 23440 17085
rect 24308 17076 24360 17128
rect 25320 17119 25372 17128
rect 25320 17085 25329 17119
rect 25329 17085 25363 17119
rect 25363 17085 25372 17119
rect 25320 17076 25372 17085
rect 27160 17212 27212 17264
rect 27068 17144 27120 17196
rect 38200 17187 38252 17196
rect 38200 17153 38209 17187
rect 38209 17153 38243 17187
rect 38243 17153 38252 17187
rect 38200 17144 38252 17153
rect 13176 16983 13228 16992
rect 13176 16949 13185 16983
rect 13185 16949 13219 16983
rect 13219 16949 13228 16983
rect 13176 16940 13228 16949
rect 13820 16983 13872 16992
rect 13820 16949 13829 16983
rect 13829 16949 13863 16983
rect 13863 16949 13872 16983
rect 13820 16940 13872 16949
rect 14188 16940 14240 16992
rect 16396 16940 16448 16992
rect 20996 16940 21048 16992
rect 22192 16983 22244 16992
rect 22192 16949 22201 16983
rect 22201 16949 22235 16983
rect 22235 16949 22244 16983
rect 22192 16940 22244 16949
rect 22652 16940 22704 16992
rect 26240 17076 26292 17128
rect 26056 17008 26108 17060
rect 27804 17008 27856 17060
rect 35900 17008 35952 17060
rect 26148 16940 26200 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2228 16736 2280 16788
rect 20168 16736 20220 16788
rect 23204 16736 23256 16788
rect 15844 16668 15896 16720
rect 14372 16643 14424 16652
rect 8208 16464 8260 16516
rect 12624 16464 12676 16516
rect 13176 16532 13228 16584
rect 14372 16609 14381 16643
rect 14381 16609 14415 16643
rect 14415 16609 14424 16643
rect 14372 16600 14424 16609
rect 15292 16600 15344 16652
rect 14464 16507 14516 16516
rect 14464 16473 14473 16507
rect 14473 16473 14507 16507
rect 14507 16473 14516 16507
rect 15016 16507 15068 16516
rect 14464 16464 14516 16473
rect 15016 16473 15025 16507
rect 15025 16473 15059 16507
rect 15059 16473 15068 16507
rect 15016 16464 15068 16473
rect 16212 16600 16264 16652
rect 16580 16575 16632 16584
rect 16580 16541 16589 16575
rect 16589 16541 16623 16575
rect 16623 16541 16632 16575
rect 16580 16532 16632 16541
rect 17592 16668 17644 16720
rect 18052 16668 18104 16720
rect 19708 16668 19760 16720
rect 17868 16643 17920 16652
rect 17868 16609 17877 16643
rect 17877 16609 17911 16643
rect 17911 16609 17920 16643
rect 17868 16600 17920 16609
rect 20444 16600 20496 16652
rect 20904 16668 20956 16720
rect 22560 16600 22612 16652
rect 21548 16575 21600 16584
rect 21548 16541 21557 16575
rect 21557 16541 21591 16575
rect 21591 16541 21600 16575
rect 21548 16532 21600 16541
rect 11244 16396 11296 16448
rect 12716 16396 12768 16448
rect 12992 16439 13044 16448
rect 12992 16405 13001 16439
rect 13001 16405 13035 16439
rect 13035 16405 13044 16439
rect 12992 16396 13044 16405
rect 14556 16396 14608 16448
rect 15752 16396 15804 16448
rect 17224 16439 17276 16448
rect 17224 16405 17233 16439
rect 17233 16405 17267 16439
rect 17267 16405 17276 16439
rect 17224 16396 17276 16405
rect 17684 16396 17736 16448
rect 18052 16464 18104 16516
rect 19616 16507 19668 16516
rect 19616 16473 19625 16507
rect 19625 16473 19659 16507
rect 19659 16473 19668 16507
rect 19616 16464 19668 16473
rect 20076 16464 20128 16516
rect 20260 16507 20312 16516
rect 20260 16473 20269 16507
rect 20269 16473 20303 16507
rect 20303 16473 20312 16507
rect 20260 16464 20312 16473
rect 20720 16464 20772 16516
rect 21364 16464 21416 16516
rect 20628 16396 20680 16448
rect 20812 16396 20864 16448
rect 22652 16464 22704 16516
rect 23020 16464 23072 16516
rect 24860 16600 24912 16652
rect 25044 16600 25096 16652
rect 25780 16668 25832 16720
rect 26056 16643 26108 16652
rect 26056 16609 26065 16643
rect 26065 16609 26099 16643
rect 26099 16609 26108 16643
rect 26056 16600 26108 16609
rect 26424 16643 26476 16652
rect 26424 16609 26433 16643
rect 26433 16609 26467 16643
rect 26467 16609 26476 16643
rect 26424 16600 26476 16609
rect 26792 16532 26844 16584
rect 27344 16600 27396 16652
rect 24584 16507 24636 16516
rect 24584 16473 24593 16507
rect 24593 16473 24627 16507
rect 24627 16473 24636 16507
rect 24584 16464 24636 16473
rect 26332 16507 26384 16516
rect 23388 16439 23440 16448
rect 23388 16405 23397 16439
rect 23397 16405 23431 16439
rect 23431 16405 23440 16439
rect 23388 16396 23440 16405
rect 26332 16473 26341 16507
rect 26341 16473 26375 16507
rect 26375 16473 26384 16507
rect 26332 16464 26384 16473
rect 26424 16464 26476 16516
rect 30288 16464 30340 16516
rect 26148 16396 26200 16448
rect 26608 16396 26660 16448
rect 28448 16396 28500 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 11060 16192 11112 16244
rect 12992 16167 13044 16176
rect 12992 16133 13001 16167
rect 13001 16133 13035 16167
rect 13035 16133 13044 16167
rect 12992 16124 13044 16133
rect 17316 16192 17368 16244
rect 18328 16235 18380 16244
rect 18328 16201 18337 16235
rect 18337 16201 18371 16235
rect 18371 16201 18380 16235
rect 18328 16192 18380 16201
rect 15752 16167 15804 16176
rect 15752 16133 15761 16167
rect 15761 16133 15795 16167
rect 15795 16133 15804 16167
rect 15752 16124 15804 16133
rect 16396 16124 16448 16176
rect 8116 16056 8168 16108
rect 11152 16099 11204 16108
rect 11152 16065 11161 16099
rect 11161 16065 11195 16099
rect 11195 16065 11204 16099
rect 21548 16192 21600 16244
rect 20352 16124 20404 16176
rect 22192 16192 22244 16244
rect 26240 16192 26292 16244
rect 26332 16192 26384 16244
rect 11152 16056 11204 16065
rect 19064 16099 19116 16108
rect 12900 16031 12952 16040
rect 12900 15997 12909 16031
rect 12909 15997 12943 16031
rect 12943 15997 12952 16031
rect 12900 15988 12952 15997
rect 9772 15920 9824 15972
rect 12532 15920 12584 15972
rect 12624 15920 12676 15972
rect 13544 15920 13596 15972
rect 14372 15988 14424 16040
rect 15108 15988 15160 16040
rect 16764 15988 16816 16040
rect 16948 16031 17000 16040
rect 16948 15997 16957 16031
rect 16957 15997 16991 16031
rect 16991 15997 17000 16031
rect 16948 15988 17000 15997
rect 19064 16065 19073 16099
rect 19073 16065 19107 16099
rect 19107 16065 19116 16099
rect 19064 16056 19116 16065
rect 22008 16099 22060 16108
rect 22008 16065 22017 16099
rect 22017 16065 22051 16099
rect 22051 16065 22060 16099
rect 22008 16056 22060 16065
rect 23572 16124 23624 16176
rect 24032 16124 24084 16176
rect 24492 16167 24544 16176
rect 24492 16133 24501 16167
rect 24501 16133 24535 16167
rect 24535 16133 24544 16167
rect 24492 16124 24544 16133
rect 38016 16124 38068 16176
rect 15568 15920 15620 15972
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 18788 15988 18840 16040
rect 23204 16031 23256 16040
rect 23204 15997 23213 16031
rect 23213 15997 23247 16031
rect 23247 15997 23256 16031
rect 23204 15988 23256 15997
rect 17960 15920 18012 15972
rect 19156 15920 19208 15972
rect 20444 15963 20496 15972
rect 20444 15929 20453 15963
rect 20453 15929 20487 15963
rect 20487 15929 20496 15963
rect 20444 15920 20496 15929
rect 20628 15920 20680 15972
rect 22100 15920 22152 15972
rect 23756 15988 23808 16040
rect 24768 15988 24820 16040
rect 26516 16056 26568 16108
rect 25780 16031 25832 16040
rect 15752 15852 15804 15904
rect 18144 15852 18196 15904
rect 20076 15852 20128 15904
rect 23480 15920 23532 15972
rect 25504 15920 25556 15972
rect 25780 15997 25789 16031
rect 25789 15997 25823 16031
rect 25823 15997 25832 16031
rect 25780 15988 25832 15997
rect 25964 15988 26016 16040
rect 26792 16056 26844 16108
rect 27160 16099 27212 16108
rect 27160 16065 27169 16099
rect 27169 16065 27203 16099
rect 27203 16065 27212 16099
rect 27160 16056 27212 16065
rect 27988 16099 28040 16108
rect 27988 16065 27997 16099
rect 27997 16065 28031 16099
rect 28031 16065 28040 16099
rect 27988 16056 28040 16065
rect 28448 16099 28500 16108
rect 28448 16065 28457 16099
rect 28457 16065 28491 16099
rect 28491 16065 28500 16099
rect 28448 16056 28500 16065
rect 38200 16099 38252 16108
rect 38200 16065 38209 16099
rect 38209 16065 38243 16099
rect 38243 16065 38252 16099
rect 38200 16056 38252 16065
rect 30196 15920 30248 15972
rect 38016 15963 38068 15972
rect 38016 15929 38025 15963
rect 38025 15929 38059 15963
rect 38059 15929 38068 15963
rect 38016 15920 38068 15929
rect 23204 15852 23256 15904
rect 23664 15852 23716 15904
rect 26332 15852 26384 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 8116 15691 8168 15700
rect 8116 15657 8125 15691
rect 8125 15657 8159 15691
rect 8159 15657 8168 15691
rect 8116 15648 8168 15657
rect 9680 15691 9732 15700
rect 9680 15657 9689 15691
rect 9689 15657 9723 15691
rect 9723 15657 9732 15691
rect 9680 15648 9732 15657
rect 14464 15648 14516 15700
rect 15108 15648 15160 15700
rect 17868 15648 17920 15700
rect 18788 15691 18840 15700
rect 18788 15657 18797 15691
rect 18797 15657 18831 15691
rect 18831 15657 18840 15691
rect 18788 15648 18840 15657
rect 14280 15580 14332 15632
rect 15568 15580 15620 15632
rect 16948 15580 17000 15632
rect 17224 15580 17276 15632
rect 19524 15580 19576 15632
rect 10968 15512 11020 15564
rect 8208 15487 8260 15496
rect 8208 15453 8217 15487
rect 8217 15453 8251 15487
rect 8251 15453 8260 15487
rect 8208 15444 8260 15453
rect 9680 15444 9732 15496
rect 11152 15487 11204 15496
rect 11152 15453 11161 15487
rect 11161 15453 11195 15487
rect 11195 15453 11204 15487
rect 11152 15444 11204 15453
rect 20536 15648 20588 15700
rect 23940 15648 23992 15700
rect 27436 15648 27488 15700
rect 36636 15648 36688 15700
rect 19984 15580 20036 15632
rect 20444 15580 20496 15632
rect 24584 15580 24636 15632
rect 12716 15444 12768 15496
rect 12900 15444 12952 15496
rect 11796 15308 11848 15360
rect 12440 15308 12492 15360
rect 13636 15308 13688 15360
rect 14556 15376 14608 15428
rect 15108 15376 15160 15428
rect 16304 15419 16356 15428
rect 16304 15385 16313 15419
rect 16313 15385 16347 15419
rect 16347 15385 16356 15419
rect 16304 15376 16356 15385
rect 20260 15512 20312 15564
rect 23112 15555 23164 15564
rect 23112 15521 23121 15555
rect 23121 15521 23155 15555
rect 23155 15521 23164 15555
rect 23112 15512 23164 15521
rect 23388 15555 23440 15564
rect 23388 15521 23397 15555
rect 23397 15521 23431 15555
rect 23431 15521 23440 15555
rect 23388 15512 23440 15521
rect 23572 15512 23624 15564
rect 26976 15512 27028 15564
rect 18512 15444 18564 15496
rect 19892 15444 19944 15496
rect 20536 15444 20588 15496
rect 21916 15444 21968 15496
rect 22928 15444 22980 15496
rect 25504 15444 25556 15496
rect 28540 15512 28592 15564
rect 27252 15444 27304 15496
rect 29000 15444 29052 15496
rect 17500 15419 17552 15428
rect 17500 15385 17509 15419
rect 17509 15385 17543 15419
rect 17543 15385 17552 15419
rect 17500 15376 17552 15385
rect 17960 15376 18012 15428
rect 16856 15308 16908 15360
rect 17408 15308 17460 15360
rect 20076 15376 20128 15428
rect 20444 15376 20496 15428
rect 20996 15419 21048 15428
rect 20996 15385 21005 15419
rect 21005 15385 21039 15419
rect 21039 15385 21048 15419
rect 21548 15419 21600 15428
rect 20996 15376 21048 15385
rect 21548 15385 21557 15419
rect 21557 15385 21591 15419
rect 21591 15385 21600 15419
rect 21548 15376 21600 15385
rect 18144 15351 18196 15360
rect 18144 15317 18153 15351
rect 18153 15317 18187 15351
rect 18187 15317 18196 15351
rect 20260 15351 20312 15360
rect 18144 15308 18196 15317
rect 20260 15317 20269 15351
rect 20269 15317 20303 15351
rect 20303 15317 20312 15351
rect 20260 15308 20312 15317
rect 22928 15308 22980 15360
rect 24952 15376 25004 15428
rect 25136 15419 25188 15428
rect 25136 15385 25145 15419
rect 25145 15385 25179 15419
rect 25179 15385 25188 15419
rect 25136 15376 25188 15385
rect 26332 15419 26384 15428
rect 26332 15385 26341 15419
rect 26341 15385 26375 15419
rect 26375 15385 26384 15419
rect 26332 15376 26384 15385
rect 26424 15419 26476 15428
rect 26424 15385 26433 15419
rect 26433 15385 26467 15419
rect 26467 15385 26476 15419
rect 26424 15376 26476 15385
rect 26792 15376 26844 15428
rect 24768 15308 24820 15360
rect 27712 15351 27764 15360
rect 27712 15317 27721 15351
rect 27721 15317 27755 15351
rect 27755 15317 27764 15351
rect 27712 15308 27764 15317
rect 28172 15308 28224 15360
rect 28540 15308 28592 15360
rect 30932 15308 30984 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 11060 15147 11112 15156
rect 11060 15113 11069 15147
rect 11069 15113 11103 15147
rect 11103 15113 11112 15147
rect 11060 15104 11112 15113
rect 15016 15104 15068 15156
rect 17960 15104 18012 15156
rect 20352 15147 20404 15156
rect 10232 14968 10284 15020
rect 10416 14968 10468 15020
rect 10968 15011 11020 15020
rect 10968 14977 10977 15011
rect 10977 14977 11011 15011
rect 11011 14977 11020 15011
rect 10968 14968 11020 14977
rect 12164 15011 12216 15020
rect 12164 14977 12173 15011
rect 12173 14977 12207 15011
rect 12207 14977 12216 15011
rect 12164 14968 12216 14977
rect 13084 15036 13136 15088
rect 13544 15079 13596 15088
rect 13544 15045 13553 15079
rect 13553 15045 13587 15079
rect 13587 15045 13596 15079
rect 13544 15036 13596 15045
rect 14188 15079 14240 15088
rect 14188 15045 14197 15079
rect 14197 15045 14231 15079
rect 14231 15045 14240 15079
rect 14188 15036 14240 15045
rect 15384 15079 15436 15088
rect 15384 15045 15393 15079
rect 15393 15045 15427 15079
rect 15427 15045 15436 15079
rect 15384 15036 15436 15045
rect 16028 15036 16080 15088
rect 18144 15036 18196 15088
rect 18604 15079 18656 15088
rect 18604 15045 18613 15079
rect 18613 15045 18647 15079
rect 18647 15045 18656 15079
rect 18604 15036 18656 15045
rect 18880 15036 18932 15088
rect 19340 15036 19392 15088
rect 19892 15036 19944 15088
rect 17868 14968 17920 15020
rect 12440 14900 12492 14952
rect 13084 14900 13136 14952
rect 9312 14832 9364 14884
rect 10324 14832 10376 14884
rect 12072 14832 12124 14884
rect 14832 14900 14884 14952
rect 11428 14764 11480 14816
rect 14648 14875 14700 14884
rect 14648 14841 14657 14875
rect 14657 14841 14691 14875
rect 14691 14841 14700 14875
rect 15476 14900 15528 14952
rect 17592 14943 17644 14952
rect 14648 14832 14700 14841
rect 16304 14832 16356 14884
rect 17592 14909 17601 14943
rect 17601 14909 17635 14943
rect 17635 14909 17644 14943
rect 17592 14900 17644 14909
rect 19432 14968 19484 15020
rect 19800 15011 19852 15020
rect 19800 14977 19809 15011
rect 19809 14977 19843 15011
rect 19843 14977 19852 15011
rect 19800 14968 19852 14977
rect 20352 15113 20361 15147
rect 20361 15113 20395 15147
rect 20395 15113 20404 15147
rect 20352 15104 20404 15113
rect 21364 15147 21416 15156
rect 21364 15113 21373 15147
rect 21373 15113 21407 15147
rect 21407 15113 21416 15147
rect 21364 15104 21416 15113
rect 20076 15036 20128 15088
rect 24400 15104 24452 15156
rect 24952 15104 25004 15156
rect 20536 14968 20588 15020
rect 21272 15011 21324 15020
rect 21272 14977 21281 15011
rect 21281 14977 21315 15011
rect 21315 14977 21324 15011
rect 21272 14968 21324 14977
rect 21364 14968 21416 15020
rect 22376 15036 22428 15088
rect 22468 15036 22520 15088
rect 23572 15079 23624 15088
rect 23572 15045 23581 15079
rect 23581 15045 23615 15079
rect 23615 15045 23624 15079
rect 23572 15036 23624 15045
rect 24676 15079 24728 15088
rect 24676 15045 24685 15079
rect 24685 15045 24719 15079
rect 24719 15045 24728 15079
rect 24676 15036 24728 15045
rect 24768 15079 24820 15088
rect 24768 15045 24777 15079
rect 24777 15045 24811 15079
rect 24811 15045 24820 15079
rect 24768 15036 24820 15045
rect 25964 15036 26016 15088
rect 26424 15104 26476 15156
rect 27344 15011 27396 15020
rect 27344 14977 27353 15011
rect 27353 14977 27387 15011
rect 27387 14977 27396 15011
rect 27344 14968 27396 14977
rect 27528 14968 27580 15020
rect 28632 15011 28684 15020
rect 28632 14977 28641 15011
rect 28641 14977 28675 15011
rect 28675 14977 28684 15011
rect 29644 15011 29696 15020
rect 28632 14968 28684 14977
rect 29644 14977 29653 15011
rect 29653 14977 29687 15011
rect 29687 14977 29696 15011
rect 29644 14968 29696 14977
rect 19248 14900 19300 14952
rect 21916 14900 21968 14952
rect 22192 14943 22244 14952
rect 22192 14909 22201 14943
rect 22201 14909 22235 14943
rect 22235 14909 22244 14943
rect 22192 14900 22244 14909
rect 22376 14900 22428 14952
rect 22836 14900 22888 14952
rect 20720 14832 20772 14884
rect 22008 14832 22060 14884
rect 24952 14900 25004 14952
rect 25504 14900 25556 14952
rect 26424 14900 26476 14952
rect 17040 14764 17092 14816
rect 19432 14764 19484 14816
rect 23020 14764 23072 14816
rect 23848 14764 23900 14816
rect 24400 14832 24452 14884
rect 28448 14832 28500 14884
rect 25412 14764 25464 14816
rect 26516 14807 26568 14816
rect 26516 14773 26525 14807
rect 26525 14773 26559 14807
rect 26559 14773 26568 14807
rect 26516 14764 26568 14773
rect 26700 14764 26752 14816
rect 29000 14764 29052 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 3424 14560 3476 14612
rect 11980 14560 12032 14612
rect 12164 14560 12216 14612
rect 21364 14560 21416 14612
rect 21916 14560 21968 14612
rect 23940 14560 23992 14612
rect 24676 14560 24728 14612
rect 12256 14492 12308 14544
rect 17500 14492 17552 14544
rect 18696 14492 18748 14544
rect 20720 14492 20772 14544
rect 9404 14424 9456 14476
rect 9312 14399 9364 14408
rect 9312 14365 9321 14399
rect 9321 14365 9355 14399
rect 9355 14365 9364 14399
rect 9312 14356 9364 14365
rect 9772 14399 9824 14408
rect 9772 14365 9781 14399
rect 9781 14365 9815 14399
rect 9815 14365 9824 14399
rect 9772 14356 9824 14365
rect 16764 14424 16816 14476
rect 16948 14467 17000 14476
rect 16948 14433 16957 14467
rect 16957 14433 16991 14467
rect 16991 14433 17000 14467
rect 16948 14424 17000 14433
rect 17408 14424 17460 14476
rect 19432 14424 19484 14476
rect 20352 14467 20404 14476
rect 20352 14433 20361 14467
rect 20361 14433 20395 14467
rect 20395 14433 20404 14467
rect 20352 14424 20404 14433
rect 22008 14492 22060 14544
rect 24952 14492 25004 14544
rect 25044 14492 25096 14544
rect 10508 14399 10560 14408
rect 10508 14365 10517 14399
rect 10517 14365 10551 14399
rect 10551 14365 10560 14399
rect 10508 14356 10560 14365
rect 11980 14356 12032 14408
rect 12532 14399 12584 14408
rect 12532 14365 12541 14399
rect 12541 14365 12575 14399
rect 12575 14365 12584 14399
rect 12532 14356 12584 14365
rect 13820 14356 13872 14408
rect 14372 14356 14424 14408
rect 14924 14356 14976 14408
rect 16304 14399 16356 14408
rect 16304 14365 16313 14399
rect 16313 14365 16347 14399
rect 16347 14365 16356 14399
rect 16304 14356 16356 14365
rect 16396 14356 16448 14408
rect 17960 14356 18012 14408
rect 19340 14356 19392 14408
rect 13084 14331 13136 14340
rect 13084 14297 13093 14331
rect 13093 14297 13127 14331
rect 13127 14297 13136 14331
rect 13084 14288 13136 14297
rect 13176 14331 13228 14340
rect 13176 14297 13185 14331
rect 13185 14297 13219 14331
rect 13219 14297 13228 14331
rect 13728 14331 13780 14340
rect 13176 14288 13228 14297
rect 13728 14297 13737 14331
rect 13737 14297 13771 14331
rect 13771 14297 13780 14331
rect 13728 14288 13780 14297
rect 14740 14288 14792 14340
rect 17500 14331 17552 14340
rect 1676 14263 1728 14272
rect 1676 14229 1685 14263
rect 1685 14229 1719 14263
rect 1719 14229 1728 14263
rect 1676 14220 1728 14229
rect 11888 14263 11940 14272
rect 11888 14229 11897 14263
rect 11897 14229 11931 14263
rect 11931 14229 11940 14263
rect 11888 14220 11940 14229
rect 14188 14220 14240 14272
rect 17500 14297 17509 14331
rect 17509 14297 17543 14331
rect 17543 14297 17552 14331
rect 17500 14288 17552 14297
rect 18972 14288 19024 14340
rect 20168 14220 20220 14272
rect 20812 14288 20864 14340
rect 20996 14288 21048 14340
rect 21364 14220 21416 14272
rect 23112 14467 23164 14476
rect 23112 14433 23121 14467
rect 23121 14433 23155 14467
rect 23155 14433 23164 14467
rect 23112 14424 23164 14433
rect 23388 14424 23440 14476
rect 25136 14424 25188 14476
rect 22376 14331 22428 14340
rect 22376 14297 22385 14331
rect 22385 14297 22419 14331
rect 22419 14297 22428 14331
rect 22376 14288 22428 14297
rect 22928 14288 22980 14340
rect 24032 14220 24084 14272
rect 25504 14331 25556 14340
rect 25504 14297 25513 14331
rect 25513 14297 25547 14331
rect 25547 14297 25556 14331
rect 25504 14288 25556 14297
rect 25964 14288 26016 14340
rect 26608 14331 26660 14340
rect 26608 14297 26617 14331
rect 26617 14297 26651 14331
rect 26651 14297 26660 14331
rect 26608 14288 26660 14297
rect 26976 14356 27028 14408
rect 27528 14356 27580 14408
rect 29000 14424 29052 14476
rect 28540 14399 28592 14408
rect 28540 14365 28549 14399
rect 28549 14365 28583 14399
rect 28583 14365 28592 14399
rect 28540 14356 28592 14365
rect 27068 14220 27120 14272
rect 27528 14220 27580 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 11612 14016 11664 14068
rect 11888 14016 11940 14068
rect 12440 14016 12492 14068
rect 9772 13948 9824 14000
rect 10324 13948 10376 14000
rect 11244 13948 11296 14000
rect 18420 14016 18472 14068
rect 7840 13812 7892 13864
rect 10876 13812 10928 13864
rect 11152 13880 11204 13932
rect 13912 13948 13964 14000
rect 11428 13880 11480 13932
rect 11244 13744 11296 13796
rect 12348 13787 12400 13796
rect 7932 13676 7984 13728
rect 11704 13676 11756 13728
rect 12348 13753 12357 13787
rect 12357 13753 12391 13787
rect 12391 13753 12400 13787
rect 12348 13744 12400 13753
rect 12440 13744 12492 13796
rect 12808 13744 12860 13796
rect 12532 13676 12584 13728
rect 13360 13812 13412 13864
rect 13636 13812 13688 13864
rect 13820 13812 13872 13864
rect 16672 13948 16724 14000
rect 17040 13991 17092 14000
rect 17040 13957 17049 13991
rect 17049 13957 17083 13991
rect 17083 13957 17092 13991
rect 17040 13948 17092 13957
rect 19064 13948 19116 14000
rect 20260 13948 20312 14000
rect 14464 13855 14516 13864
rect 14464 13821 14473 13855
rect 14473 13821 14507 13855
rect 14507 13821 14516 13855
rect 14464 13812 14516 13821
rect 14648 13812 14700 13864
rect 14924 13812 14976 13864
rect 16304 13880 16356 13932
rect 18696 13923 18748 13932
rect 18696 13889 18705 13923
rect 18705 13889 18739 13923
rect 18739 13889 18748 13923
rect 18696 13880 18748 13889
rect 16948 13855 17000 13864
rect 16948 13821 16957 13855
rect 16957 13821 16991 13855
rect 16991 13821 17000 13855
rect 16948 13812 17000 13821
rect 19156 13812 19208 13864
rect 19432 13812 19484 13864
rect 20444 14016 20496 14068
rect 28264 14016 28316 14068
rect 20812 13880 20864 13932
rect 21180 13880 21232 13932
rect 23112 13948 23164 14000
rect 23388 13991 23440 14000
rect 23388 13957 23397 13991
rect 23397 13957 23431 13991
rect 23431 13957 23440 13991
rect 23940 13991 23992 14000
rect 23388 13948 23440 13957
rect 23940 13957 23949 13991
rect 23949 13957 23983 13991
rect 23983 13957 23992 13991
rect 23940 13948 23992 13957
rect 25320 13948 25372 14000
rect 25412 13948 25464 14000
rect 25964 13948 26016 14000
rect 24032 13880 24084 13932
rect 21272 13855 21324 13864
rect 13912 13744 13964 13796
rect 14740 13744 14792 13796
rect 14556 13676 14608 13728
rect 14648 13676 14700 13728
rect 18144 13744 18196 13796
rect 18236 13744 18288 13796
rect 21272 13821 21281 13855
rect 21281 13821 21315 13855
rect 21315 13821 21324 13855
rect 21272 13812 21324 13821
rect 21824 13812 21876 13864
rect 23388 13812 23440 13864
rect 25044 13812 25096 13864
rect 16212 13676 16264 13728
rect 20628 13676 20680 13728
rect 21732 13744 21784 13796
rect 22008 13676 22060 13728
rect 24032 13744 24084 13796
rect 26884 13880 26936 13932
rect 27344 13923 27396 13932
rect 27344 13889 27353 13923
rect 27353 13889 27387 13923
rect 27387 13889 27396 13923
rect 27344 13880 27396 13889
rect 27528 13880 27580 13932
rect 25780 13812 25832 13864
rect 27252 13812 27304 13864
rect 27896 13855 27948 13864
rect 27896 13821 27905 13855
rect 27905 13821 27939 13855
rect 27939 13821 27948 13855
rect 27896 13812 27948 13821
rect 28080 13880 28132 13932
rect 28724 13880 28776 13932
rect 29276 13923 29328 13932
rect 29276 13889 29285 13923
rect 29285 13889 29319 13923
rect 29319 13889 29328 13923
rect 29276 13880 29328 13889
rect 29460 13880 29512 13932
rect 38200 13923 38252 13932
rect 38200 13889 38209 13923
rect 38209 13889 38243 13923
rect 38243 13889 38252 13923
rect 38200 13880 38252 13889
rect 29828 13812 29880 13864
rect 24676 13676 24728 13728
rect 27620 13744 27672 13796
rect 27252 13719 27304 13728
rect 27252 13685 27261 13719
rect 27261 13685 27295 13719
rect 27295 13685 27304 13719
rect 27252 13676 27304 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 10968 13472 11020 13524
rect 9128 13404 9180 13456
rect 13544 13472 13596 13524
rect 11704 13404 11756 13456
rect 12164 13404 12216 13456
rect 13360 13404 13412 13456
rect 13728 13472 13780 13524
rect 14464 13404 14516 13456
rect 16212 13472 16264 13524
rect 16304 13472 16356 13524
rect 18236 13472 18288 13524
rect 18604 13472 18656 13524
rect 21732 13472 21784 13524
rect 22008 13472 22060 13524
rect 27068 13515 27120 13524
rect 11060 13336 11112 13388
rect 8852 13268 8904 13320
rect 18512 13379 18564 13388
rect 18512 13345 18521 13379
rect 18521 13345 18555 13379
rect 18555 13345 18564 13379
rect 18512 13336 18564 13345
rect 19064 13336 19116 13388
rect 19524 13379 19576 13388
rect 19524 13345 19533 13379
rect 19533 13345 19567 13379
rect 19567 13345 19576 13379
rect 19524 13336 19576 13345
rect 19892 13336 19944 13388
rect 21916 13336 21968 13388
rect 23020 13379 23072 13388
rect 23020 13345 23029 13379
rect 23029 13345 23063 13379
rect 23063 13345 23072 13379
rect 23020 13336 23072 13345
rect 23388 13404 23440 13456
rect 23940 13336 23992 13388
rect 24124 13336 24176 13388
rect 24952 13379 25004 13388
rect 24952 13345 24961 13379
rect 24961 13345 24995 13379
rect 24995 13345 25004 13379
rect 24952 13336 25004 13345
rect 25780 13404 25832 13456
rect 27068 13481 27077 13515
rect 27077 13481 27111 13515
rect 27111 13481 27120 13515
rect 27068 13472 27120 13481
rect 27344 13472 27396 13524
rect 25964 13404 26016 13456
rect 28632 13404 28684 13456
rect 26056 13336 26108 13388
rect 28540 13336 28592 13388
rect 28724 13336 28776 13388
rect 11244 13311 11296 13320
rect 11244 13277 11253 13311
rect 11253 13277 11287 13311
rect 11287 13277 11296 13311
rect 11244 13268 11296 13277
rect 11796 13268 11848 13320
rect 12072 13311 12124 13320
rect 12072 13277 12081 13311
rect 12081 13277 12115 13311
rect 12115 13277 12124 13311
rect 12072 13268 12124 13277
rect 12164 13268 12216 13320
rect 14464 13311 14516 13320
rect 9864 13200 9916 13252
rect 12348 13200 12400 13252
rect 14464 13277 14473 13311
rect 14473 13277 14507 13311
rect 14507 13277 14516 13311
rect 14464 13268 14516 13277
rect 20260 13268 20312 13320
rect 20904 13268 20956 13320
rect 13084 13243 13136 13252
rect 13084 13209 13093 13243
rect 13093 13209 13127 13243
rect 13127 13209 13136 13243
rect 13084 13200 13136 13209
rect 10600 13132 10652 13184
rect 10968 13132 11020 13184
rect 11796 13132 11848 13184
rect 12256 13132 12308 13184
rect 13360 13200 13412 13252
rect 13820 13132 13872 13184
rect 14556 13200 14608 13252
rect 15476 13132 15528 13184
rect 16764 13243 16816 13252
rect 16764 13209 16773 13243
rect 16773 13209 16807 13243
rect 16807 13209 16816 13243
rect 16764 13200 16816 13209
rect 18236 13200 18288 13252
rect 19616 13243 19668 13252
rect 19616 13209 19625 13243
rect 19625 13209 19659 13243
rect 19659 13209 19668 13243
rect 19616 13200 19668 13209
rect 20352 13200 20404 13252
rect 21088 13200 21140 13252
rect 20536 13132 20588 13184
rect 24032 13200 24084 13252
rect 26792 13268 26844 13320
rect 26976 13311 27028 13320
rect 26976 13277 26985 13311
rect 26985 13277 27019 13311
rect 27019 13277 27028 13311
rect 26976 13268 27028 13277
rect 24952 13200 25004 13252
rect 25136 13243 25188 13252
rect 25136 13209 25145 13243
rect 25145 13209 25179 13243
rect 25179 13209 25188 13243
rect 25136 13200 25188 13209
rect 25228 13200 25280 13252
rect 25688 13200 25740 13252
rect 27528 13200 27580 13252
rect 27804 13200 27856 13252
rect 28172 13243 28224 13252
rect 28172 13209 28181 13243
rect 28181 13209 28215 13243
rect 28215 13209 28224 13243
rect 28172 13200 28224 13209
rect 28264 13243 28316 13252
rect 28264 13209 28273 13243
rect 28273 13209 28307 13243
rect 28307 13209 28316 13243
rect 28264 13200 28316 13209
rect 23480 13132 23532 13184
rect 24124 13132 24176 13184
rect 26700 13132 26752 13184
rect 27068 13132 27120 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 7932 12928 7984 12980
rect 9128 12971 9180 12980
rect 9128 12937 9137 12971
rect 9137 12937 9171 12971
rect 9171 12937 9180 12971
rect 9128 12928 9180 12937
rect 11980 12928 12032 12980
rect 13452 12928 13504 12980
rect 18236 12928 18288 12980
rect 18696 12928 18748 12980
rect 19432 12928 19484 12980
rect 5540 12792 5592 12844
rect 7748 12835 7800 12844
rect 7748 12801 7757 12835
rect 7757 12801 7791 12835
rect 7791 12801 7800 12835
rect 7748 12792 7800 12801
rect 9680 12860 9732 12912
rect 9036 12835 9088 12844
rect 9036 12801 9045 12835
rect 9045 12801 9079 12835
rect 9079 12801 9088 12835
rect 9036 12792 9088 12801
rect 9864 12835 9916 12844
rect 9864 12801 9873 12835
rect 9873 12801 9907 12835
rect 9907 12801 9916 12835
rect 9864 12792 9916 12801
rect 10692 12792 10744 12844
rect 10968 12835 11020 12844
rect 10968 12801 10977 12835
rect 10977 12801 11011 12835
rect 11011 12801 11020 12835
rect 10968 12792 11020 12801
rect 11152 12860 11204 12912
rect 11520 12860 11572 12912
rect 11612 12860 11664 12912
rect 12072 12860 12124 12912
rect 15384 12860 15436 12912
rect 17224 12860 17276 12912
rect 16396 12792 16448 12844
rect 13084 12724 13136 12776
rect 14188 12724 14240 12776
rect 14740 12767 14792 12776
rect 14740 12733 14749 12767
rect 14749 12733 14783 12767
rect 14783 12733 14792 12767
rect 14740 12724 14792 12733
rect 15016 12767 15068 12776
rect 15016 12733 15025 12767
rect 15025 12733 15059 12767
rect 15059 12733 15068 12767
rect 15016 12724 15068 12733
rect 15476 12724 15528 12776
rect 18328 12860 18380 12912
rect 20444 12903 20496 12912
rect 20444 12869 20453 12903
rect 20453 12869 20487 12903
rect 20487 12869 20496 12903
rect 20444 12860 20496 12869
rect 20812 12928 20864 12980
rect 22744 12928 22796 12980
rect 21364 12860 21416 12912
rect 21732 12860 21784 12912
rect 22928 12860 22980 12912
rect 23480 12903 23532 12912
rect 23480 12869 23489 12903
rect 23489 12869 23523 12903
rect 23523 12869 23532 12903
rect 23480 12860 23532 12869
rect 24124 12860 24176 12912
rect 17408 12835 17460 12844
rect 17408 12801 17417 12835
rect 17417 12801 17451 12835
rect 17451 12801 17460 12835
rect 17408 12792 17460 12801
rect 17776 12792 17828 12844
rect 12072 12656 12124 12708
rect 12348 12699 12400 12708
rect 12348 12665 12357 12699
rect 12357 12665 12391 12699
rect 12391 12665 12400 12699
rect 12348 12656 12400 12665
rect 14924 12656 14976 12708
rect 1676 12631 1728 12640
rect 1676 12597 1685 12631
rect 1685 12597 1719 12631
rect 1719 12597 1728 12631
rect 1676 12588 1728 12597
rect 10784 12588 10836 12640
rect 18236 12724 18288 12776
rect 18512 12767 18564 12776
rect 18512 12733 18521 12767
rect 18521 12733 18555 12767
rect 18555 12733 18564 12767
rect 18512 12724 18564 12733
rect 19340 12724 19392 12776
rect 19524 12724 19576 12776
rect 23388 12792 23440 12844
rect 20996 12724 21048 12776
rect 22284 12767 22336 12776
rect 22284 12733 22293 12767
rect 22293 12733 22327 12767
rect 22327 12733 22336 12767
rect 22284 12724 22336 12733
rect 25872 12928 25924 12980
rect 27528 12928 27580 12980
rect 24676 12903 24728 12912
rect 24676 12869 24685 12903
rect 24685 12869 24719 12903
rect 24719 12869 24728 12903
rect 24676 12860 24728 12869
rect 25044 12860 25096 12912
rect 25780 12860 25832 12912
rect 35900 12928 35952 12980
rect 23388 12656 23440 12708
rect 25688 12792 25740 12844
rect 26056 12835 26108 12844
rect 26056 12801 26065 12835
rect 26065 12801 26099 12835
rect 26099 12801 26108 12835
rect 26056 12792 26108 12801
rect 15936 12588 15988 12640
rect 18512 12588 18564 12640
rect 18696 12588 18748 12640
rect 21548 12588 21600 12640
rect 22928 12588 22980 12640
rect 23940 12588 23992 12640
rect 28632 12835 28684 12844
rect 28632 12801 28641 12835
rect 28641 12801 28675 12835
rect 28675 12801 28684 12835
rect 28632 12792 28684 12801
rect 28724 12724 28776 12776
rect 27712 12656 27764 12708
rect 27528 12588 27580 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 5540 12384 5592 12436
rect 10140 12384 10192 12436
rect 10784 12384 10836 12436
rect 11244 12427 11296 12436
rect 11244 12393 11253 12427
rect 11253 12393 11287 12427
rect 11287 12393 11296 12427
rect 11244 12384 11296 12393
rect 9772 12316 9824 12368
rect 11152 12316 11204 12368
rect 19708 12384 19760 12436
rect 13176 12316 13228 12368
rect 13452 12316 13504 12368
rect 14556 12316 14608 12368
rect 16396 12316 16448 12368
rect 17040 12316 17092 12368
rect 12900 12248 12952 12300
rect 13360 12248 13412 12300
rect 13728 12291 13780 12300
rect 13728 12257 13737 12291
rect 13737 12257 13771 12291
rect 13771 12257 13780 12291
rect 13728 12248 13780 12257
rect 14004 12248 14056 12300
rect 14924 12248 14976 12300
rect 1860 12044 1912 12096
rect 2596 12044 2648 12096
rect 7748 12112 7800 12164
rect 9036 12180 9088 12232
rect 9496 12180 9548 12232
rect 10692 12223 10744 12232
rect 10692 12189 10701 12223
rect 10701 12189 10735 12223
rect 10735 12189 10744 12223
rect 10692 12180 10744 12189
rect 11704 12180 11756 12232
rect 18880 12316 18932 12368
rect 20352 12384 20404 12436
rect 20444 12384 20496 12436
rect 20720 12316 20772 12368
rect 25780 12384 25832 12436
rect 27620 12384 27672 12436
rect 29828 12427 29880 12436
rect 29828 12393 29837 12427
rect 29837 12393 29871 12427
rect 29871 12393 29880 12427
rect 29828 12384 29880 12393
rect 30288 12384 30340 12436
rect 38016 12384 38068 12436
rect 23296 12316 23348 12368
rect 23664 12316 23716 12368
rect 18972 12248 19024 12300
rect 19248 12248 19300 12300
rect 20260 12248 20312 12300
rect 20352 12248 20404 12300
rect 23388 12291 23440 12300
rect 19432 12223 19484 12232
rect 19432 12189 19441 12223
rect 19441 12189 19475 12223
rect 19475 12189 19484 12223
rect 19432 12180 19484 12189
rect 21364 12180 21416 12232
rect 22284 12223 22336 12232
rect 22284 12189 22293 12223
rect 22293 12189 22327 12223
rect 22327 12189 22336 12223
rect 22284 12180 22336 12189
rect 8760 12112 8812 12164
rect 9588 12112 9640 12164
rect 10416 12044 10468 12096
rect 11428 12112 11480 12164
rect 11980 12155 12032 12164
rect 11980 12121 11989 12155
rect 11989 12121 12023 12155
rect 12023 12121 12032 12155
rect 11980 12112 12032 12121
rect 12532 12112 12584 12164
rect 12716 12112 12768 12164
rect 13728 12112 13780 12164
rect 13452 12044 13504 12096
rect 15568 12112 15620 12164
rect 16672 12155 16724 12164
rect 16672 12121 16681 12155
rect 16681 12121 16715 12155
rect 16715 12121 16724 12155
rect 16672 12112 16724 12121
rect 17316 12112 17368 12164
rect 19340 12112 19392 12164
rect 19708 12112 19760 12164
rect 21732 12112 21784 12164
rect 19064 12044 19116 12096
rect 20812 12044 20864 12096
rect 23388 12257 23397 12291
rect 23397 12257 23431 12291
rect 23431 12257 23440 12291
rect 23388 12248 23440 12257
rect 23572 12248 23624 12300
rect 27436 12316 27488 12368
rect 25136 12248 25188 12300
rect 27896 12248 27948 12300
rect 26608 12180 26660 12232
rect 27436 12180 27488 12232
rect 27620 12223 27672 12232
rect 27620 12189 27629 12223
rect 27629 12189 27663 12223
rect 27663 12189 27672 12223
rect 27620 12180 27672 12189
rect 27988 12180 28040 12232
rect 28908 12180 28960 12232
rect 22928 12112 22980 12164
rect 23204 12112 23256 12164
rect 23480 12155 23532 12164
rect 23480 12121 23489 12155
rect 23489 12121 23523 12155
rect 23523 12121 23532 12155
rect 23480 12112 23532 12121
rect 23664 12112 23716 12164
rect 24860 12112 24912 12164
rect 25136 12155 25188 12164
rect 25136 12121 25145 12155
rect 25145 12121 25179 12155
rect 25179 12121 25188 12155
rect 25136 12112 25188 12121
rect 25228 12155 25280 12164
rect 25228 12121 25237 12155
rect 25237 12121 25271 12155
rect 25271 12121 25280 12155
rect 25228 12112 25280 12121
rect 25504 12112 25556 12164
rect 28356 12087 28408 12096
rect 28356 12053 28365 12087
rect 28365 12053 28399 12087
rect 28399 12053 28408 12087
rect 28356 12044 28408 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 9036 11840 9088 11892
rect 10324 11840 10376 11892
rect 11152 11840 11204 11892
rect 12256 11772 12308 11824
rect 12532 11772 12584 11824
rect 12900 11772 12952 11824
rect 13728 11772 13780 11824
rect 13912 11772 13964 11824
rect 14924 11815 14976 11824
rect 14924 11781 14933 11815
rect 14933 11781 14967 11815
rect 14967 11781 14976 11815
rect 14924 11772 14976 11781
rect 17316 11840 17368 11892
rect 23664 11840 23716 11892
rect 18236 11815 18288 11824
rect 8116 11704 8168 11756
rect 10508 11747 10560 11756
rect 10508 11713 10517 11747
rect 10517 11713 10551 11747
rect 10551 11713 10560 11747
rect 10508 11704 10560 11713
rect 10968 11704 11020 11756
rect 11152 11747 11204 11756
rect 11152 11713 11161 11747
rect 11161 11713 11195 11747
rect 11195 11713 11204 11747
rect 11152 11704 11204 11713
rect 16304 11747 16356 11756
rect 16304 11713 16313 11747
rect 16313 11713 16347 11747
rect 16347 11713 16356 11747
rect 17040 11747 17092 11756
rect 16304 11704 16356 11713
rect 17040 11713 17049 11747
rect 17049 11713 17083 11747
rect 17083 11713 17092 11747
rect 17040 11704 17092 11713
rect 11060 11568 11112 11620
rect 11244 11568 11296 11620
rect 11336 11568 11388 11620
rect 12440 11568 12492 11620
rect 13176 11636 13228 11688
rect 14004 11636 14056 11688
rect 17592 11636 17644 11688
rect 15476 11568 15528 11620
rect 18236 11781 18245 11815
rect 18245 11781 18279 11815
rect 18279 11781 18288 11815
rect 18236 11772 18288 11781
rect 19064 11815 19116 11824
rect 19064 11781 19073 11815
rect 19073 11781 19107 11815
rect 19107 11781 19116 11815
rect 19064 11772 19116 11781
rect 20168 11772 20220 11824
rect 20812 11772 20864 11824
rect 22376 11772 22428 11824
rect 21364 11747 21416 11756
rect 21364 11713 21373 11747
rect 21373 11713 21407 11747
rect 21407 11713 21416 11747
rect 21364 11704 21416 11713
rect 21548 11704 21600 11756
rect 21824 11704 21876 11756
rect 23020 11772 23072 11824
rect 23940 11772 23992 11824
rect 24584 11772 24636 11824
rect 24860 11815 24912 11824
rect 24860 11781 24869 11815
rect 24869 11781 24903 11815
rect 24903 11781 24912 11815
rect 24860 11772 24912 11781
rect 26332 11772 26384 11824
rect 27896 11772 27948 11824
rect 23204 11704 23256 11756
rect 27344 11747 27396 11756
rect 17868 11679 17920 11688
rect 17868 11645 17877 11679
rect 17877 11645 17911 11679
rect 17911 11645 17920 11679
rect 17868 11636 17920 11645
rect 18696 11636 18748 11688
rect 18972 11679 19024 11688
rect 18972 11645 18981 11679
rect 18981 11645 19015 11679
rect 19015 11645 19024 11679
rect 18972 11636 19024 11645
rect 19984 11636 20036 11688
rect 19156 11568 19208 11620
rect 22100 11679 22152 11688
rect 22100 11645 22109 11679
rect 22109 11645 22143 11679
rect 22143 11645 22152 11679
rect 22100 11636 22152 11645
rect 23572 11636 23624 11688
rect 25228 11636 25280 11688
rect 25504 11679 25556 11688
rect 25504 11645 25513 11679
rect 25513 11645 25547 11679
rect 25547 11645 25556 11679
rect 25504 11636 25556 11645
rect 27344 11713 27353 11747
rect 27353 11713 27387 11747
rect 27387 11713 27396 11747
rect 27344 11704 27396 11713
rect 27436 11704 27488 11756
rect 28448 11747 28500 11756
rect 28448 11713 28457 11747
rect 28457 11713 28491 11747
rect 28491 11713 28500 11747
rect 28448 11704 28500 11713
rect 38200 11747 38252 11756
rect 38200 11713 38209 11747
rect 38209 11713 38243 11747
rect 38243 11713 38252 11747
rect 38200 11704 38252 11713
rect 22560 11568 22612 11620
rect 23388 11568 23440 11620
rect 7288 11543 7340 11552
rect 7288 11509 7297 11543
rect 7297 11509 7331 11543
rect 7331 11509 7340 11543
rect 7288 11500 7340 11509
rect 9128 11543 9180 11552
rect 9128 11509 9137 11543
rect 9137 11509 9171 11543
rect 9171 11509 9180 11543
rect 9128 11500 9180 11509
rect 10416 11500 10468 11552
rect 13360 11500 13412 11552
rect 20720 11500 20772 11552
rect 23480 11500 23532 11552
rect 30748 11568 30800 11620
rect 25872 11500 25924 11552
rect 27068 11500 27120 11552
rect 27252 11543 27304 11552
rect 27252 11509 27261 11543
rect 27261 11509 27295 11543
rect 27295 11509 27304 11543
rect 27252 11500 27304 11509
rect 27528 11500 27580 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 13452 11296 13504 11348
rect 13636 11296 13688 11348
rect 15568 11296 15620 11348
rect 11612 11228 11664 11280
rect 15016 11228 15068 11280
rect 12256 11160 12308 11212
rect 13544 11160 13596 11212
rect 11336 11135 11388 11144
rect 11336 11101 11345 11135
rect 11345 11101 11379 11135
rect 11379 11101 11388 11135
rect 11336 11092 11388 11101
rect 14004 11092 14056 11144
rect 14924 11135 14976 11144
rect 14924 11101 14933 11135
rect 14933 11101 14967 11135
rect 14967 11101 14976 11135
rect 14924 11092 14976 11101
rect 2872 11024 2924 11076
rect 7840 11024 7892 11076
rect 8576 11067 8628 11076
rect 8576 11033 8585 11067
rect 8585 11033 8619 11067
rect 8619 11033 8628 11067
rect 8576 11024 8628 11033
rect 9496 11024 9548 11076
rect 9772 11067 9824 11076
rect 9772 11033 9781 11067
rect 9781 11033 9815 11067
rect 9815 11033 9824 11067
rect 9772 11024 9824 11033
rect 10324 11067 10376 11076
rect 10324 11033 10333 11067
rect 10333 11033 10367 11067
rect 10367 11033 10376 11067
rect 10324 11024 10376 11033
rect 10416 11024 10468 11076
rect 11428 11024 11480 11076
rect 11520 11024 11572 11076
rect 9220 10999 9272 11008
rect 9220 10965 9229 10999
rect 9229 10965 9263 10999
rect 9263 10965 9272 10999
rect 9220 10956 9272 10965
rect 9864 10956 9916 11008
rect 13176 11067 13228 11076
rect 13176 11033 13185 11067
rect 13185 11033 13219 11067
rect 13219 11033 13228 11067
rect 13176 11024 13228 11033
rect 13452 11024 13504 11076
rect 16212 11228 16264 11280
rect 19156 11228 19208 11280
rect 19432 11228 19484 11280
rect 19892 11296 19944 11348
rect 21272 11296 21324 11348
rect 21364 11296 21416 11348
rect 27252 11296 27304 11348
rect 20628 11228 20680 11280
rect 22376 11228 22428 11280
rect 22560 11228 22612 11280
rect 24676 11271 24728 11280
rect 24676 11237 24685 11271
rect 24685 11237 24719 11271
rect 24719 11237 24728 11271
rect 24676 11228 24728 11237
rect 15476 11203 15528 11212
rect 15476 11169 15485 11203
rect 15485 11169 15519 11203
rect 15519 11169 15528 11203
rect 15476 11160 15528 11169
rect 19248 11160 19300 11212
rect 19892 11203 19944 11212
rect 19892 11169 19901 11203
rect 19901 11169 19935 11203
rect 19935 11169 19944 11203
rect 19892 11160 19944 11169
rect 22100 11160 22152 11212
rect 22284 11160 22336 11212
rect 24584 11160 24636 11212
rect 18512 11092 18564 11144
rect 20444 11092 20496 11144
rect 15568 11067 15620 11076
rect 15568 11033 15577 11067
rect 15577 11033 15611 11067
rect 15611 11033 15620 11067
rect 15568 11024 15620 11033
rect 18144 11067 18196 11076
rect 12716 10956 12768 11008
rect 13820 10956 13872 11008
rect 18144 11033 18153 11067
rect 18153 11033 18187 11067
rect 18187 11033 18196 11067
rect 18144 11024 18196 11033
rect 18696 11024 18748 11076
rect 18052 10956 18104 11008
rect 19064 10956 19116 11008
rect 19524 10956 19576 11008
rect 20076 10956 20128 11008
rect 20720 11067 20772 11076
rect 20720 11033 20729 11067
rect 20729 11033 20763 11067
rect 20763 11033 20772 11067
rect 20720 11024 20772 11033
rect 21272 11024 21324 11076
rect 20904 10956 20956 11008
rect 21364 10956 21416 11008
rect 21916 11067 21968 11076
rect 21916 11033 21925 11067
rect 21925 11033 21959 11067
rect 21959 11033 21968 11067
rect 21916 11024 21968 11033
rect 22284 11024 22336 11076
rect 23480 11067 23532 11076
rect 23480 11033 23489 11067
rect 23489 11033 23523 11067
rect 23523 11033 23532 11067
rect 23480 11024 23532 11033
rect 28356 11228 28408 11280
rect 25780 11203 25832 11212
rect 25780 11169 25789 11203
rect 25789 11169 25823 11203
rect 25823 11169 25832 11203
rect 26424 11203 26476 11212
rect 25780 11160 25832 11169
rect 26424 11169 26433 11203
rect 26433 11169 26467 11203
rect 26467 11169 26476 11203
rect 26424 11160 26476 11169
rect 26608 11160 26660 11212
rect 27988 11092 28040 11144
rect 23388 10956 23440 11008
rect 26148 11024 26200 11076
rect 26332 11067 26384 11076
rect 26332 11033 26341 11067
rect 26341 11033 26375 11067
rect 26375 11033 26384 11067
rect 26332 11024 26384 11033
rect 27620 10956 27672 11008
rect 28264 10999 28316 11008
rect 28264 10965 28273 10999
rect 28273 10965 28307 10999
rect 28307 10965 28316 10999
rect 28264 10956 28316 10965
rect 30196 10956 30248 11008
rect 34796 10956 34848 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 8760 10795 8812 10804
rect 8760 10761 8769 10795
rect 8769 10761 8803 10795
rect 8803 10761 8812 10795
rect 8760 10752 8812 10761
rect 9220 10752 9272 10804
rect 12256 10684 12308 10736
rect 13084 10684 13136 10736
rect 13268 10684 13320 10736
rect 14004 10684 14056 10736
rect 14740 10752 14792 10804
rect 14648 10684 14700 10736
rect 16580 10684 16632 10736
rect 1584 10616 1636 10668
rect 8852 10616 8904 10668
rect 11244 10616 11296 10668
rect 11336 10616 11388 10668
rect 8852 10480 8904 10532
rect 10968 10480 11020 10532
rect 12256 10548 12308 10600
rect 12532 10548 12584 10600
rect 13268 10591 13320 10600
rect 11612 10480 11664 10532
rect 13268 10557 13277 10591
rect 13277 10557 13311 10591
rect 13311 10557 13320 10591
rect 13268 10548 13320 10557
rect 14004 10548 14056 10600
rect 14924 10548 14976 10600
rect 17040 10616 17092 10668
rect 18512 10752 18564 10804
rect 19156 10752 19208 10804
rect 21272 10752 21324 10804
rect 21640 10752 21692 10804
rect 19524 10616 19576 10668
rect 20168 10684 20220 10736
rect 20996 10616 21048 10668
rect 18880 10548 18932 10600
rect 19064 10548 19116 10600
rect 21272 10548 21324 10600
rect 14832 10480 14884 10532
rect 15016 10523 15068 10532
rect 15016 10489 15025 10523
rect 15025 10489 15059 10523
rect 15059 10489 15068 10523
rect 15016 10480 15068 10489
rect 8116 10455 8168 10464
rect 8116 10421 8125 10455
rect 8125 10421 8159 10455
rect 8159 10421 8168 10455
rect 8116 10412 8168 10421
rect 11060 10455 11112 10464
rect 11060 10421 11069 10455
rect 11069 10421 11103 10455
rect 11103 10421 11112 10455
rect 11060 10412 11112 10421
rect 12532 10412 12584 10464
rect 12808 10412 12860 10464
rect 24860 10727 24912 10736
rect 24860 10693 24869 10727
rect 24869 10693 24903 10727
rect 24903 10693 24912 10727
rect 24860 10684 24912 10693
rect 25780 10684 25832 10736
rect 28264 10684 28316 10736
rect 21640 10548 21692 10600
rect 23756 10548 23808 10600
rect 29000 10616 29052 10668
rect 38200 10659 38252 10668
rect 38200 10625 38209 10659
rect 38209 10625 38243 10659
rect 38243 10625 38252 10659
rect 38200 10616 38252 10625
rect 25136 10548 25188 10600
rect 25596 10591 25648 10600
rect 25596 10557 25605 10591
rect 25605 10557 25639 10591
rect 25639 10557 25648 10591
rect 25596 10548 25648 10557
rect 25688 10548 25740 10600
rect 27068 10548 27120 10600
rect 27896 10591 27948 10600
rect 27896 10557 27905 10591
rect 27905 10557 27939 10591
rect 27939 10557 27948 10591
rect 27896 10548 27948 10557
rect 28816 10548 28868 10600
rect 27712 10480 27764 10532
rect 28356 10480 28408 10532
rect 37004 10480 37056 10532
rect 22836 10412 22888 10464
rect 25136 10412 25188 10464
rect 28908 10412 28960 10464
rect 29368 10455 29420 10464
rect 29368 10421 29377 10455
rect 29377 10421 29411 10455
rect 29411 10421 29420 10455
rect 29368 10412 29420 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 1584 10251 1636 10260
rect 1584 10217 1593 10251
rect 1593 10217 1627 10251
rect 1627 10217 1636 10251
rect 1584 10208 1636 10217
rect 8760 10208 8812 10260
rect 9680 10208 9732 10260
rect 10968 10208 11020 10260
rect 11060 10208 11112 10260
rect 16672 10208 16724 10260
rect 9036 10140 9088 10192
rect 10508 10140 10560 10192
rect 10600 10140 10652 10192
rect 9864 10115 9916 10124
rect 9864 10081 9873 10115
rect 9873 10081 9907 10115
rect 9907 10081 9916 10115
rect 9864 10072 9916 10081
rect 8760 10004 8812 10056
rect 12164 10140 12216 10192
rect 12992 10140 13044 10192
rect 16396 10140 16448 10192
rect 10968 10004 11020 10056
rect 11336 10004 11388 10056
rect 14924 10072 14976 10124
rect 15200 10072 15252 10124
rect 17500 10208 17552 10260
rect 19156 10208 19208 10260
rect 21364 10208 21416 10260
rect 18420 10140 18472 10192
rect 19248 10140 19300 10192
rect 19616 10140 19668 10192
rect 23296 10208 23348 10260
rect 25044 10208 25096 10260
rect 25964 10208 26016 10260
rect 29092 10208 29144 10260
rect 17040 10115 17092 10124
rect 17040 10081 17049 10115
rect 17049 10081 17083 10115
rect 17083 10081 17092 10115
rect 17040 10072 17092 10081
rect 17316 10115 17368 10124
rect 17316 10081 17325 10115
rect 17325 10081 17359 10115
rect 17359 10081 17368 10115
rect 17316 10072 17368 10081
rect 17868 10072 17920 10124
rect 14464 10004 14516 10056
rect 20904 10072 20956 10124
rect 21640 10115 21692 10124
rect 21640 10081 21649 10115
rect 21649 10081 21683 10115
rect 21683 10081 21692 10115
rect 21640 10072 21692 10081
rect 25136 10140 25188 10192
rect 25320 10140 25372 10192
rect 26608 10140 26660 10192
rect 28264 10140 28316 10192
rect 22284 10072 22336 10124
rect 12256 9979 12308 9988
rect 9404 9868 9456 9920
rect 11244 9868 11296 9920
rect 12256 9945 12265 9979
rect 12265 9945 12299 9979
rect 12299 9945 12308 9979
rect 12256 9936 12308 9945
rect 12808 9936 12860 9988
rect 13360 9936 13412 9988
rect 14924 9936 14976 9988
rect 16488 9936 16540 9988
rect 16764 9936 16816 9988
rect 17316 9936 17368 9988
rect 18328 9936 18380 9988
rect 20352 10004 20404 10056
rect 24768 10004 24820 10056
rect 27528 10004 27580 10056
rect 29368 10072 29420 10124
rect 29000 10047 29052 10056
rect 29000 10013 29009 10047
rect 29009 10013 29043 10047
rect 29043 10013 29052 10047
rect 30196 10047 30248 10056
rect 29000 10004 29052 10013
rect 30196 10013 30205 10047
rect 30205 10013 30239 10047
rect 30239 10013 30248 10047
rect 30196 10004 30248 10013
rect 19616 9936 19668 9988
rect 20904 9979 20956 9988
rect 20904 9945 20913 9979
rect 20913 9945 20947 9979
rect 20947 9945 20956 9979
rect 20904 9936 20956 9945
rect 21456 9936 21508 9988
rect 21916 9979 21968 9988
rect 21916 9945 21925 9979
rect 21925 9945 21959 9979
rect 21959 9945 21968 9979
rect 21916 9936 21968 9945
rect 24676 9936 24728 9988
rect 25044 9979 25096 9988
rect 25044 9945 25053 9979
rect 25053 9945 25087 9979
rect 25087 9945 25096 9979
rect 25964 9979 26016 9988
rect 25044 9936 25096 9945
rect 25964 9945 25973 9979
rect 25973 9945 26007 9979
rect 26007 9945 26016 9979
rect 25964 9936 26016 9945
rect 26148 9936 26200 9988
rect 27068 9979 27120 9988
rect 27068 9945 27077 9979
rect 27077 9945 27111 9979
rect 27111 9945 27120 9979
rect 27068 9936 27120 9945
rect 28632 9936 28684 9988
rect 29920 9979 29972 9988
rect 29920 9945 29929 9979
rect 29929 9945 29963 9979
rect 29963 9945 29972 9979
rect 29920 9936 29972 9945
rect 13176 9868 13228 9920
rect 18788 9911 18840 9920
rect 18788 9877 18797 9911
rect 18797 9877 18831 9911
rect 18831 9877 18840 9911
rect 18788 9868 18840 9877
rect 19156 9868 19208 9920
rect 19708 9868 19760 9920
rect 20628 9868 20680 9920
rect 23296 9868 23348 9920
rect 23388 9911 23440 9920
rect 23388 9877 23397 9911
rect 23397 9877 23431 9911
rect 23431 9877 23440 9911
rect 23388 9868 23440 9877
rect 26240 9868 26292 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 9128 9664 9180 9716
rect 12808 9664 12860 9716
rect 14004 9707 14056 9716
rect 9680 9596 9732 9648
rect 10324 9596 10376 9648
rect 11244 9596 11296 9648
rect 14004 9673 14013 9707
rect 14013 9673 14047 9707
rect 14047 9673 14056 9707
rect 14004 9664 14056 9673
rect 14832 9664 14884 9716
rect 14740 9596 14792 9648
rect 13268 9528 13320 9580
rect 17960 9664 18012 9716
rect 19064 9664 19116 9716
rect 16488 9596 16540 9648
rect 18144 9596 18196 9648
rect 20996 9664 21048 9716
rect 12348 9460 12400 9512
rect 12624 9460 12676 9512
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 7196 9392 7248 9444
rect 12900 9392 12952 9444
rect 8760 9367 8812 9376
rect 8760 9333 8769 9367
rect 8769 9333 8803 9367
rect 8803 9333 8812 9367
rect 8760 9324 8812 9333
rect 10416 9324 10468 9376
rect 10784 9324 10836 9376
rect 13912 9324 13964 9376
rect 14004 9324 14056 9376
rect 15752 9324 15804 9376
rect 20168 9571 20220 9580
rect 20168 9537 20177 9571
rect 20177 9537 20211 9571
rect 20211 9537 20220 9571
rect 20168 9528 20220 9537
rect 20352 9528 20404 9580
rect 16764 9460 16816 9512
rect 16856 9460 16908 9512
rect 17776 9460 17828 9512
rect 16396 9392 16448 9444
rect 19340 9460 19392 9512
rect 22192 9596 22244 9648
rect 24216 9596 24268 9648
rect 24400 9639 24452 9648
rect 24400 9605 24409 9639
rect 24409 9605 24443 9639
rect 24443 9605 24452 9639
rect 24400 9596 24452 9605
rect 21640 9528 21692 9580
rect 24124 9528 24176 9580
rect 24768 9664 24820 9716
rect 27436 9664 27488 9716
rect 24952 9639 25004 9648
rect 24952 9605 24961 9639
rect 24961 9605 24995 9639
rect 24995 9605 25004 9639
rect 24952 9596 25004 9605
rect 26240 9596 26292 9648
rect 26424 9596 26476 9648
rect 26332 9571 26384 9580
rect 26332 9537 26341 9571
rect 26341 9537 26375 9571
rect 26375 9537 26384 9571
rect 26332 9528 26384 9537
rect 27528 9596 27580 9648
rect 27620 9596 27672 9648
rect 28356 9664 28408 9716
rect 28540 9664 28592 9716
rect 28172 9596 28224 9648
rect 37004 9596 37056 9648
rect 29920 9528 29972 9580
rect 22054 9448 22106 9500
rect 22376 9460 22428 9512
rect 22652 9460 22704 9512
rect 24860 9460 24912 9512
rect 24952 9460 25004 9512
rect 27068 9460 27120 9512
rect 27160 9460 27212 9512
rect 27804 9460 27856 9512
rect 27896 9460 27948 9512
rect 29092 9503 29144 9512
rect 29092 9469 29101 9503
rect 29101 9469 29135 9503
rect 29135 9469 29144 9503
rect 29092 9460 29144 9469
rect 29368 9460 29420 9512
rect 21180 9392 21232 9444
rect 21548 9392 21600 9444
rect 23296 9392 23348 9444
rect 27528 9392 27580 9444
rect 27620 9392 27672 9444
rect 29000 9392 29052 9444
rect 20076 9324 20128 9376
rect 20720 9367 20772 9376
rect 20720 9333 20729 9367
rect 20729 9333 20763 9367
rect 20763 9333 20772 9367
rect 20720 9324 20772 9333
rect 20812 9324 20864 9376
rect 21272 9324 21324 9376
rect 22008 9324 22060 9376
rect 22744 9324 22796 9376
rect 23388 9324 23440 9376
rect 23756 9367 23808 9376
rect 23756 9333 23765 9367
rect 23765 9333 23799 9367
rect 23799 9333 23808 9367
rect 23756 9324 23808 9333
rect 24124 9324 24176 9376
rect 33692 9324 33744 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 9772 9120 9824 9172
rect 11336 9120 11388 9172
rect 11520 9163 11572 9172
rect 11520 9129 11529 9163
rect 11529 9129 11563 9163
rect 11563 9129 11572 9163
rect 11520 9120 11572 9129
rect 11796 9120 11848 9172
rect 13820 9052 13872 9104
rect 14372 9052 14424 9104
rect 16488 9052 16540 9104
rect 7288 8984 7340 9036
rect 10048 8984 10100 9036
rect 10784 8984 10836 9036
rect 12624 9027 12676 9036
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 10968 8959 11020 8968
rect 10968 8925 10977 8959
rect 10977 8925 11011 8959
rect 11011 8925 11020 8959
rect 10968 8916 11020 8925
rect 12624 8993 12633 9027
rect 12633 8993 12667 9027
rect 12667 8993 12676 9027
rect 12624 8984 12676 8993
rect 14648 8984 14700 9036
rect 16396 9027 16448 9036
rect 16396 8993 16405 9027
rect 16405 8993 16439 9027
rect 16439 8993 16448 9027
rect 16396 8984 16448 8993
rect 14004 8916 14056 8968
rect 14372 8959 14424 8968
rect 14372 8925 14381 8959
rect 14381 8925 14415 8959
rect 14415 8925 14424 8959
rect 14372 8916 14424 8925
rect 18144 9052 18196 9104
rect 18972 9052 19024 9104
rect 20720 9052 20772 9104
rect 22284 9052 22336 9104
rect 24584 9120 24636 9172
rect 24768 9120 24820 9172
rect 30748 9163 30800 9172
rect 30748 9129 30757 9163
rect 30757 9129 30791 9163
rect 30791 9129 30800 9163
rect 30748 9120 30800 9129
rect 26792 9052 26844 9104
rect 16856 9027 16908 9036
rect 16856 8993 16865 9027
rect 16865 8993 16899 9027
rect 16899 8993 16908 9027
rect 16856 8984 16908 8993
rect 17132 8984 17184 9036
rect 11060 8848 11112 8900
rect 12164 8891 12216 8900
rect 12164 8857 12173 8891
rect 12173 8857 12207 8891
rect 12207 8857 12216 8891
rect 12164 8848 12216 8857
rect 14556 8848 14608 8900
rect 17408 8848 17460 8900
rect 18788 8848 18840 8900
rect 12348 8780 12400 8832
rect 18144 8780 18196 8832
rect 21088 8984 21140 9036
rect 21640 8984 21692 9036
rect 24308 8984 24360 9036
rect 24400 8984 24452 9036
rect 25872 8984 25924 9036
rect 27160 8984 27212 9036
rect 27712 9052 27764 9104
rect 30564 8984 30616 9036
rect 19616 8959 19668 8968
rect 19616 8925 19625 8959
rect 19625 8925 19659 8959
rect 19659 8925 19668 8959
rect 19616 8916 19668 8925
rect 20168 8959 20220 8968
rect 20168 8925 20177 8959
rect 20177 8925 20211 8959
rect 20211 8925 20220 8959
rect 20168 8916 20220 8925
rect 20996 8916 21048 8968
rect 24768 8959 24820 8968
rect 24768 8925 24777 8959
rect 24777 8925 24811 8959
rect 24811 8925 24820 8959
rect 24768 8916 24820 8925
rect 20536 8848 20588 8900
rect 20720 8848 20772 8900
rect 20904 8891 20956 8900
rect 20904 8857 20913 8891
rect 20913 8857 20947 8891
rect 20947 8857 20956 8891
rect 20904 8848 20956 8857
rect 23204 8848 23256 8900
rect 21732 8780 21784 8832
rect 22284 8780 22336 8832
rect 25136 8848 25188 8900
rect 26516 8848 26568 8900
rect 26608 8780 26660 8832
rect 28172 8959 28224 8968
rect 28172 8925 28181 8959
rect 28181 8925 28215 8959
rect 28215 8925 28224 8959
rect 28172 8916 28224 8925
rect 30196 8959 30248 8968
rect 28816 8848 28868 8900
rect 30196 8925 30205 8959
rect 30205 8925 30239 8959
rect 30239 8925 30248 8959
rect 30196 8916 30248 8925
rect 33048 8916 33100 8968
rect 37924 9120 37976 9172
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 10968 8576 11020 8628
rect 13912 8576 13964 8628
rect 14188 8576 14240 8628
rect 18144 8576 18196 8628
rect 22560 8576 22612 8628
rect 11244 8508 11296 8560
rect 12072 8508 12124 8560
rect 14740 8551 14792 8560
rect 9772 8440 9824 8492
rect 14740 8517 14749 8551
rect 14749 8517 14783 8551
rect 14783 8517 14792 8551
rect 14740 8508 14792 8517
rect 18512 8508 18564 8560
rect 24124 8576 24176 8628
rect 24308 8619 24360 8628
rect 24308 8585 24317 8619
rect 24317 8585 24351 8619
rect 24351 8585 24360 8619
rect 24308 8576 24360 8585
rect 24676 8508 24728 8560
rect 25872 8508 25924 8560
rect 27252 8576 27304 8628
rect 27988 8576 28040 8628
rect 28172 8576 28224 8628
rect 28908 8576 28960 8628
rect 29184 8619 29236 8628
rect 29184 8585 29193 8619
rect 29193 8585 29227 8619
rect 29227 8585 29236 8619
rect 29184 8576 29236 8585
rect 29828 8508 29880 8560
rect 38016 8551 38068 8560
rect 38016 8517 38025 8551
rect 38025 8517 38059 8551
rect 38059 8517 38068 8551
rect 38016 8508 38068 8517
rect 14096 8440 14148 8492
rect 17316 8483 17368 8492
rect 17316 8449 17325 8483
rect 17325 8449 17359 8483
rect 17359 8449 17368 8483
rect 17316 8440 17368 8449
rect 19984 8483 20036 8492
rect 19984 8449 19993 8483
rect 19993 8449 20027 8483
rect 20027 8449 20036 8483
rect 19984 8440 20036 8449
rect 20812 8440 20864 8492
rect 21180 8483 21232 8492
rect 21180 8449 21189 8483
rect 21189 8449 21223 8483
rect 21223 8449 21232 8483
rect 21180 8440 21232 8449
rect 11060 8372 11112 8424
rect 12072 8372 12124 8424
rect 12532 8415 12584 8424
rect 12532 8381 12541 8415
rect 12541 8381 12575 8415
rect 12575 8381 12584 8415
rect 12532 8372 12584 8381
rect 14464 8415 14516 8424
rect 14464 8381 14473 8415
rect 14473 8381 14507 8415
rect 14507 8381 14516 8415
rect 14464 8372 14516 8381
rect 2780 8347 2832 8356
rect 2780 8313 2789 8347
rect 2789 8313 2823 8347
rect 2823 8313 2832 8347
rect 2780 8304 2832 8313
rect 15752 8304 15804 8356
rect 17500 8347 17552 8356
rect 17500 8313 17509 8347
rect 17509 8313 17543 8347
rect 17543 8313 17552 8347
rect 17500 8304 17552 8313
rect 13912 8236 13964 8288
rect 15292 8236 15344 8288
rect 16028 8236 16080 8288
rect 19248 8304 19300 8356
rect 20720 8372 20772 8424
rect 20904 8372 20956 8424
rect 21640 8440 21692 8492
rect 22284 8415 22336 8424
rect 22284 8381 22293 8415
rect 22293 8381 22327 8415
rect 22327 8381 22336 8415
rect 22284 8372 22336 8381
rect 22652 8372 22704 8424
rect 24768 8440 24820 8492
rect 25780 8440 25832 8492
rect 25964 8440 26016 8492
rect 26424 8440 26476 8492
rect 27620 8440 27672 8492
rect 27988 8483 28040 8492
rect 27988 8449 27997 8483
rect 27997 8449 28031 8483
rect 28031 8449 28040 8483
rect 27988 8440 28040 8449
rect 28632 8483 28684 8492
rect 28632 8449 28641 8483
rect 28641 8449 28675 8483
rect 28675 8449 28684 8483
rect 28632 8440 28684 8449
rect 28908 8440 28960 8492
rect 30012 8440 30064 8492
rect 38200 8483 38252 8492
rect 38200 8449 38209 8483
rect 38209 8449 38243 8483
rect 38243 8449 38252 8483
rect 38200 8440 38252 8449
rect 23664 8372 23716 8424
rect 23940 8372 23992 8424
rect 24492 8372 24544 8424
rect 19340 8236 19392 8288
rect 22008 8304 22060 8356
rect 23296 8304 23348 8356
rect 22376 8236 22428 8288
rect 24768 8304 24820 8356
rect 28724 8372 28776 8424
rect 29000 8304 29052 8356
rect 26240 8236 26292 8288
rect 26884 8236 26936 8288
rect 29920 8236 29972 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 10232 8032 10284 8084
rect 12072 8032 12124 8084
rect 12256 8032 12308 8084
rect 13268 8075 13320 8084
rect 13268 8041 13277 8075
rect 13277 8041 13311 8075
rect 13311 8041 13320 8075
rect 13268 8032 13320 8041
rect 10600 7896 10652 7948
rect 17040 8032 17092 8084
rect 17776 8032 17828 8084
rect 21824 8032 21876 8084
rect 22008 8032 22060 8084
rect 24768 8032 24820 8084
rect 25044 8032 25096 8084
rect 25596 8032 25648 8084
rect 26056 8032 26108 8084
rect 26792 8075 26844 8084
rect 26792 8041 26801 8075
rect 26801 8041 26835 8075
rect 26835 8041 26844 8075
rect 26792 8032 26844 8041
rect 27528 8032 27580 8084
rect 30288 8032 30340 8084
rect 19248 7964 19300 8016
rect 21088 7964 21140 8016
rect 19340 7896 19392 7948
rect 21640 7896 21692 7948
rect 23204 7964 23256 8016
rect 24032 7896 24084 7948
rect 3332 7828 3384 7880
rect 13268 7828 13320 7880
rect 14096 7828 14148 7880
rect 14556 7871 14608 7880
rect 14556 7837 14565 7871
rect 14565 7837 14599 7871
rect 14599 7837 14608 7871
rect 14556 7828 14608 7837
rect 18788 7828 18840 7880
rect 12624 7760 12676 7812
rect 11060 7692 11112 7744
rect 12072 7692 12124 7744
rect 17132 7692 17184 7744
rect 17316 7803 17368 7812
rect 17316 7769 17325 7803
rect 17325 7769 17359 7803
rect 17359 7769 17368 7803
rect 23756 7828 23808 7880
rect 26240 7871 26292 7880
rect 26240 7837 26249 7871
rect 26249 7837 26283 7871
rect 26283 7837 26292 7871
rect 26884 7871 26936 7880
rect 26240 7828 26292 7837
rect 26884 7837 26893 7871
rect 26893 7837 26927 7871
rect 26927 7837 26936 7871
rect 26884 7828 26936 7837
rect 27252 7828 27304 7880
rect 17316 7760 17368 7769
rect 18696 7692 18748 7744
rect 21272 7760 21324 7812
rect 21732 7760 21784 7812
rect 27436 7896 27488 7948
rect 28080 7828 28132 7880
rect 28172 7871 28224 7880
rect 28172 7837 28181 7871
rect 28181 7837 28215 7871
rect 28215 7837 28224 7871
rect 28816 7871 28868 7880
rect 28172 7828 28224 7837
rect 28816 7837 28825 7871
rect 28825 7837 28859 7871
rect 28859 7837 28868 7871
rect 28816 7828 28868 7837
rect 30012 7828 30064 7880
rect 30288 7828 30340 7880
rect 20720 7692 20772 7744
rect 21088 7692 21140 7744
rect 22192 7692 22244 7744
rect 24124 7692 24176 7744
rect 27252 7692 27304 7744
rect 27436 7735 27488 7744
rect 27436 7701 27445 7735
rect 27445 7701 27479 7735
rect 27479 7701 27488 7735
rect 27436 7692 27488 7701
rect 28448 7692 28500 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 13084 7488 13136 7540
rect 15384 7488 15436 7540
rect 17684 7488 17736 7540
rect 18236 7531 18288 7540
rect 18236 7497 18245 7531
rect 18245 7497 18279 7531
rect 18279 7497 18288 7531
rect 18236 7488 18288 7497
rect 18696 7488 18748 7540
rect 22008 7488 22060 7540
rect 23848 7488 23900 7540
rect 25320 7488 25372 7540
rect 25688 7531 25740 7540
rect 25688 7497 25697 7531
rect 25697 7497 25731 7531
rect 25731 7497 25740 7531
rect 25688 7488 25740 7497
rect 26332 7531 26384 7540
rect 26332 7497 26341 7531
rect 26341 7497 26375 7531
rect 26375 7497 26384 7531
rect 26332 7488 26384 7497
rect 27252 7488 27304 7540
rect 28632 7488 28684 7540
rect 29828 7531 29880 7540
rect 29828 7497 29837 7531
rect 29837 7497 29871 7531
rect 29871 7497 29880 7531
rect 29828 7488 29880 7497
rect 1860 7463 1912 7472
rect 1860 7429 1869 7463
rect 1869 7429 1903 7463
rect 1903 7429 1912 7463
rect 1860 7420 1912 7429
rect 15016 7420 15068 7472
rect 16120 7420 16172 7472
rect 1584 7352 1636 7404
rect 13360 7395 13412 7404
rect 13360 7361 13369 7395
rect 13369 7361 13403 7395
rect 13403 7361 13412 7395
rect 13360 7352 13412 7361
rect 11796 7284 11848 7336
rect 14280 7352 14332 7404
rect 14464 7327 14516 7336
rect 14464 7293 14473 7327
rect 14473 7293 14507 7327
rect 14507 7293 14516 7327
rect 14464 7284 14516 7293
rect 17316 7420 17368 7472
rect 17408 7352 17460 7404
rect 13820 7216 13872 7268
rect 16856 7284 16908 7336
rect 17684 7352 17736 7404
rect 17868 7352 17920 7404
rect 19340 7420 19392 7472
rect 22560 7420 22612 7472
rect 24216 7420 24268 7472
rect 25596 7420 25648 7472
rect 27896 7463 27948 7472
rect 27896 7429 27905 7463
rect 27905 7429 27939 7463
rect 27939 7429 27948 7463
rect 27896 7420 27948 7429
rect 29184 7463 29236 7472
rect 17776 7284 17828 7336
rect 21180 7352 21232 7404
rect 21640 7352 21692 7404
rect 23388 7352 23440 7404
rect 19616 7284 19668 7336
rect 20260 7284 20312 7336
rect 22376 7284 22428 7336
rect 22652 7284 22704 7336
rect 26240 7352 26292 7404
rect 26424 7395 26476 7404
rect 26424 7361 26433 7395
rect 26433 7361 26467 7395
rect 26467 7361 26476 7395
rect 26424 7352 26476 7361
rect 27528 7352 27580 7404
rect 29184 7429 29193 7463
rect 29193 7429 29227 7463
rect 29227 7429 29236 7463
rect 29184 7420 29236 7429
rect 28080 7352 28132 7404
rect 28816 7352 28868 7404
rect 16120 7216 16172 7268
rect 25688 7284 25740 7336
rect 30012 7352 30064 7404
rect 29184 7284 29236 7336
rect 30288 7284 30340 7336
rect 11060 7191 11112 7200
rect 11060 7157 11069 7191
rect 11069 7157 11103 7191
rect 11103 7157 11112 7191
rect 11060 7148 11112 7157
rect 11980 7148 12032 7200
rect 14188 7148 14240 7200
rect 14924 7148 14976 7200
rect 16028 7148 16080 7200
rect 18788 7148 18840 7200
rect 30472 7259 30524 7268
rect 30472 7225 30481 7259
rect 30481 7225 30515 7259
rect 30515 7225 30524 7259
rect 30472 7216 30524 7225
rect 21272 7148 21324 7200
rect 25044 7191 25096 7200
rect 25044 7157 25053 7191
rect 25053 7157 25087 7191
rect 25087 7157 25096 7191
rect 25044 7148 25096 7157
rect 27252 7191 27304 7200
rect 27252 7157 27261 7191
rect 27261 7157 27295 7191
rect 27295 7157 27304 7191
rect 27252 7148 27304 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 1584 6987 1636 6996
rect 1584 6953 1593 6987
rect 1593 6953 1627 6987
rect 1627 6953 1636 6987
rect 1584 6944 1636 6953
rect 9680 6808 9732 6860
rect 14096 6944 14148 6996
rect 15568 6944 15620 6996
rect 21088 6944 21140 6996
rect 21272 6944 21324 6996
rect 27252 6944 27304 6996
rect 17132 6876 17184 6928
rect 17592 6876 17644 6928
rect 17684 6876 17736 6928
rect 18788 6876 18840 6928
rect 12900 6808 12952 6860
rect 11980 6783 12032 6792
rect 11980 6749 11989 6783
rect 11989 6749 12023 6783
rect 12023 6749 12032 6783
rect 11980 6740 12032 6749
rect 14556 6808 14608 6860
rect 17776 6808 17828 6860
rect 17960 6851 18012 6860
rect 17960 6817 17969 6851
rect 17969 6817 18003 6851
rect 18003 6817 18012 6851
rect 17960 6808 18012 6817
rect 15016 6740 15068 6792
rect 17224 6740 17276 6792
rect 20628 6808 20680 6860
rect 21180 6851 21232 6860
rect 21180 6817 21189 6851
rect 21189 6817 21223 6851
rect 21223 6817 21232 6851
rect 21180 6808 21232 6817
rect 22468 6876 22520 6928
rect 25044 6876 25096 6928
rect 25596 6876 25648 6928
rect 21916 6808 21968 6860
rect 25136 6808 25188 6860
rect 18880 6783 18932 6792
rect 18880 6749 18889 6783
rect 18889 6749 18923 6783
rect 18923 6749 18932 6783
rect 19616 6783 19668 6792
rect 18880 6740 18932 6749
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 23204 6740 23256 6792
rect 23664 6740 23716 6792
rect 24492 6740 24544 6792
rect 24768 6740 24820 6792
rect 25596 6783 25648 6792
rect 25596 6749 25605 6783
rect 25605 6749 25639 6783
rect 25639 6749 25648 6783
rect 25596 6740 25648 6749
rect 25688 6783 25740 6792
rect 25688 6749 25697 6783
rect 25697 6749 25731 6783
rect 25731 6749 25740 6783
rect 29276 6808 29328 6860
rect 25688 6740 25740 6749
rect 26884 6740 26936 6792
rect 28080 6783 28132 6792
rect 28080 6749 28089 6783
rect 28089 6749 28123 6783
rect 28123 6749 28132 6783
rect 28080 6740 28132 6749
rect 29184 6783 29236 6792
rect 29184 6749 29193 6783
rect 29193 6749 29227 6783
rect 29227 6749 29236 6783
rect 29184 6740 29236 6749
rect 11060 6604 11112 6656
rect 12440 6604 12492 6656
rect 13544 6604 13596 6656
rect 15292 6604 15344 6656
rect 15752 6672 15804 6724
rect 19248 6672 19300 6724
rect 17224 6604 17276 6656
rect 17592 6604 17644 6656
rect 20168 6672 20220 6724
rect 27252 6672 27304 6724
rect 19984 6604 20036 6656
rect 23664 6604 23716 6656
rect 26516 6604 26568 6656
rect 27344 6647 27396 6656
rect 27344 6613 27353 6647
rect 27353 6613 27387 6647
rect 27387 6613 27396 6647
rect 27344 6604 27396 6613
rect 27988 6647 28040 6656
rect 27988 6613 27997 6647
rect 27997 6613 28031 6647
rect 28031 6613 28040 6647
rect 27988 6604 28040 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 12624 6400 12676 6452
rect 18144 6400 18196 6452
rect 20628 6443 20680 6452
rect 12900 6332 12952 6384
rect 15108 6332 15160 6384
rect 19340 6332 19392 6384
rect 20076 6332 20128 6384
rect 20628 6409 20637 6443
rect 20637 6409 20671 6443
rect 20671 6409 20680 6443
rect 20628 6400 20680 6409
rect 27988 6400 28040 6452
rect 29644 6332 29696 6384
rect 11704 6264 11756 6316
rect 12256 6264 12308 6316
rect 13728 6264 13780 6316
rect 16120 6264 16172 6316
rect 11888 6239 11940 6248
rect 11888 6205 11897 6239
rect 11897 6205 11931 6239
rect 11931 6205 11940 6239
rect 11888 6196 11940 6205
rect 11980 6196 12032 6248
rect 10416 6128 10468 6180
rect 14556 6239 14608 6248
rect 14556 6205 14565 6239
rect 14565 6205 14599 6239
rect 14599 6205 14608 6239
rect 14556 6196 14608 6205
rect 16488 6196 16540 6248
rect 17776 6307 17828 6316
rect 17776 6273 17785 6307
rect 17785 6273 17819 6307
rect 17819 6273 17828 6307
rect 17776 6264 17828 6273
rect 19156 6264 19208 6316
rect 18604 6196 18656 6248
rect 22284 6264 22336 6316
rect 16672 6128 16724 6180
rect 9864 6060 9916 6112
rect 11060 6103 11112 6112
rect 11060 6069 11069 6103
rect 11069 6069 11103 6103
rect 11103 6069 11112 6103
rect 11060 6060 11112 6069
rect 12256 6060 12308 6112
rect 15200 6060 15252 6112
rect 15292 6060 15344 6112
rect 17132 6060 17184 6112
rect 17224 6060 17276 6112
rect 19432 6196 19484 6248
rect 21732 6196 21784 6248
rect 23572 6239 23624 6248
rect 23572 6205 23581 6239
rect 23581 6205 23615 6239
rect 23615 6205 23624 6239
rect 23848 6239 23900 6248
rect 23572 6196 23624 6205
rect 23848 6205 23857 6239
rect 23857 6205 23891 6239
rect 23891 6205 23900 6239
rect 23848 6196 23900 6205
rect 25228 6264 25280 6316
rect 27252 6307 27304 6316
rect 25688 6196 25740 6248
rect 27252 6273 27261 6307
rect 27261 6273 27295 6307
rect 27295 6273 27304 6307
rect 27252 6264 27304 6273
rect 27804 6264 27856 6316
rect 28172 6264 28224 6316
rect 38200 6307 38252 6316
rect 38200 6273 38209 6307
rect 38209 6273 38243 6307
rect 38243 6273 38252 6307
rect 38200 6264 38252 6273
rect 33140 6196 33192 6248
rect 19248 6128 19300 6180
rect 22560 6128 22612 6180
rect 24768 6128 24820 6180
rect 27344 6128 27396 6180
rect 27896 6128 27948 6180
rect 30380 6128 30432 6180
rect 20904 6060 20956 6112
rect 24952 6060 25004 6112
rect 25412 6103 25464 6112
rect 25412 6069 25421 6103
rect 25421 6069 25455 6103
rect 25455 6069 25464 6103
rect 25412 6060 25464 6069
rect 27436 6060 27488 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 10416 5899 10468 5908
rect 10416 5865 10425 5899
rect 10425 5865 10459 5899
rect 10459 5865 10468 5899
rect 10416 5856 10468 5865
rect 13728 5856 13780 5908
rect 20260 5856 20312 5908
rect 20628 5856 20680 5908
rect 9956 5788 10008 5840
rect 10324 5788 10376 5840
rect 12256 5788 12308 5840
rect 16672 5831 16724 5840
rect 16672 5797 16681 5831
rect 16681 5797 16715 5831
rect 16715 5797 16724 5831
rect 16672 5788 16724 5797
rect 18420 5788 18472 5840
rect 11980 5720 12032 5772
rect 14556 5720 14608 5772
rect 15200 5763 15252 5772
rect 15200 5729 15209 5763
rect 15209 5729 15243 5763
rect 15243 5729 15252 5763
rect 15200 5720 15252 5729
rect 17776 5720 17828 5772
rect 18144 5720 18196 5772
rect 19432 5720 19484 5772
rect 20904 5720 20956 5772
rect 23112 5856 23164 5908
rect 25872 5856 25924 5908
rect 27528 5856 27580 5908
rect 27896 5899 27948 5908
rect 27896 5865 27905 5899
rect 27905 5865 27939 5899
rect 27939 5865 27948 5899
rect 27896 5856 27948 5865
rect 23388 5788 23440 5840
rect 29092 5788 29144 5840
rect 26700 5763 26752 5772
rect 26700 5729 26709 5763
rect 26709 5729 26743 5763
rect 26743 5729 26752 5763
rect 26700 5720 26752 5729
rect 12348 5652 12400 5704
rect 21272 5652 21324 5704
rect 24584 5695 24636 5704
rect 24584 5661 24593 5695
rect 24593 5661 24627 5695
rect 24627 5661 24636 5695
rect 24584 5652 24636 5661
rect 24676 5695 24728 5704
rect 24676 5661 24685 5695
rect 24685 5661 24719 5695
rect 24719 5661 24728 5695
rect 25872 5695 25924 5704
rect 24676 5652 24728 5661
rect 25872 5661 25881 5695
rect 25881 5661 25915 5695
rect 25915 5661 25924 5695
rect 25872 5652 25924 5661
rect 28172 5652 28224 5704
rect 29184 5652 29236 5704
rect 9864 5559 9916 5568
rect 9864 5525 9873 5559
rect 9873 5525 9907 5559
rect 9907 5525 9916 5559
rect 9864 5516 9916 5525
rect 13728 5584 13780 5636
rect 11520 5516 11572 5568
rect 17408 5627 17460 5636
rect 17408 5593 17417 5627
rect 17417 5593 17451 5627
rect 17451 5593 17460 5627
rect 17408 5584 17460 5593
rect 19984 5584 20036 5636
rect 20352 5516 20404 5568
rect 20536 5516 20588 5568
rect 23388 5584 23440 5636
rect 23664 5584 23716 5636
rect 23204 5516 23256 5568
rect 24032 5516 24084 5568
rect 25412 5584 25464 5636
rect 25504 5516 25556 5568
rect 25780 5559 25832 5568
rect 25780 5525 25789 5559
rect 25789 5525 25823 5559
rect 25823 5525 25832 5559
rect 25780 5516 25832 5525
rect 25964 5516 26016 5568
rect 30380 5559 30432 5568
rect 30380 5525 30389 5559
rect 30389 5525 30423 5559
rect 30423 5525 30432 5559
rect 30380 5516 30432 5525
rect 30840 5559 30892 5568
rect 30840 5525 30849 5559
rect 30849 5525 30883 5559
rect 30883 5525 30892 5559
rect 30840 5516 30892 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 8760 5312 8812 5364
rect 11520 5244 11572 5296
rect 14740 5312 14792 5364
rect 14924 5312 14976 5364
rect 20168 5312 20220 5364
rect 14464 5244 14516 5296
rect 14832 5287 14884 5296
rect 14832 5253 14841 5287
rect 14841 5253 14875 5287
rect 14875 5253 14884 5287
rect 14832 5244 14884 5253
rect 16488 5244 16540 5296
rect 2780 5176 2832 5228
rect 11980 5176 12032 5228
rect 13728 5176 13780 5228
rect 14556 5219 14608 5228
rect 14556 5185 14565 5219
rect 14565 5185 14599 5219
rect 14599 5185 14608 5219
rect 14556 5176 14608 5185
rect 17132 5176 17184 5228
rect 17776 5244 17828 5296
rect 25780 5312 25832 5364
rect 27252 5355 27304 5364
rect 27252 5321 27261 5355
rect 27261 5321 27295 5355
rect 27295 5321 27304 5355
rect 27252 5312 27304 5321
rect 28540 5312 28592 5364
rect 22376 5244 22428 5296
rect 24768 5244 24820 5296
rect 24400 5176 24452 5228
rect 25044 5176 25096 5228
rect 13820 5108 13872 5160
rect 16304 5108 16356 5160
rect 17040 5108 17092 5160
rect 18052 5108 18104 5160
rect 19616 5151 19668 5160
rect 1676 5015 1728 5024
rect 1676 4981 1685 5015
rect 1685 4981 1719 5015
rect 1719 4981 1728 5015
rect 1676 4972 1728 4981
rect 9312 4972 9364 5024
rect 9864 4972 9916 5024
rect 11060 5015 11112 5024
rect 11060 4981 11069 5015
rect 11069 4981 11103 5015
rect 11103 4981 11112 5015
rect 11060 4972 11112 4981
rect 14556 5040 14608 5092
rect 19616 5117 19625 5151
rect 19625 5117 19659 5151
rect 19659 5117 19668 5151
rect 19616 5108 19668 5117
rect 13728 4972 13780 5024
rect 16120 4972 16172 5024
rect 19064 5040 19116 5092
rect 20628 5108 20680 5160
rect 21824 5108 21876 5160
rect 22284 5151 22336 5160
rect 22284 5117 22293 5151
rect 22293 5117 22327 5151
rect 22327 5117 22336 5151
rect 22284 5108 22336 5117
rect 22376 5108 22428 5160
rect 25412 5108 25464 5160
rect 26884 5176 26936 5228
rect 27528 5176 27580 5228
rect 27988 5219 28040 5228
rect 27988 5185 27997 5219
rect 27997 5185 28031 5219
rect 28031 5185 28040 5219
rect 27988 5176 28040 5185
rect 28080 5176 28132 5228
rect 29920 5176 29972 5228
rect 30012 5176 30064 5228
rect 38016 5151 38068 5160
rect 38016 5117 38025 5151
rect 38025 5117 38059 5151
rect 38059 5117 38068 5151
rect 38016 5108 38068 5117
rect 38292 5151 38344 5160
rect 38292 5117 38301 5151
rect 38301 5117 38335 5151
rect 38335 5117 38344 5151
rect 38292 5108 38344 5117
rect 19248 4972 19300 5024
rect 21916 5040 21968 5092
rect 23572 5040 23624 5092
rect 30380 5040 30432 5092
rect 33600 5040 33652 5092
rect 21364 5015 21416 5024
rect 21364 4981 21373 5015
rect 21373 4981 21407 5015
rect 21407 4981 21416 5015
rect 21364 4972 21416 4981
rect 21456 4972 21508 5024
rect 23480 4972 23532 5024
rect 23756 5015 23808 5024
rect 23756 4981 23765 5015
rect 23765 4981 23799 5015
rect 23799 4981 23808 5015
rect 23756 4972 23808 4981
rect 24768 5015 24820 5024
rect 24768 4981 24777 5015
rect 24777 4981 24811 5015
rect 24811 4981 24820 5015
rect 24768 4972 24820 4981
rect 26424 5015 26476 5024
rect 26424 4981 26433 5015
rect 26433 4981 26467 5015
rect 26467 4981 26476 5015
rect 26424 4972 26476 4981
rect 28816 5015 28868 5024
rect 28816 4981 28825 5015
rect 28825 4981 28859 5015
rect 28859 4981 28868 5015
rect 28816 4972 28868 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 11060 4768 11112 4820
rect 10508 4700 10560 4752
rect 11060 4632 11112 4684
rect 11980 4675 12032 4684
rect 11980 4641 11989 4675
rect 11989 4641 12023 4675
rect 12023 4641 12032 4675
rect 11980 4632 12032 4641
rect 14924 4700 14976 4752
rect 16856 4700 16908 4752
rect 18788 4768 18840 4820
rect 19340 4768 19392 4820
rect 19616 4768 19668 4820
rect 20628 4768 20680 4820
rect 21180 4768 21232 4820
rect 23572 4768 23624 4820
rect 17132 4675 17184 4684
rect 17132 4641 17141 4675
rect 17141 4641 17175 4675
rect 17175 4641 17184 4675
rect 17132 4632 17184 4641
rect 20076 4675 20128 4684
rect 20076 4641 20085 4675
rect 20085 4641 20119 4675
rect 20119 4641 20128 4675
rect 20076 4632 20128 4641
rect 13636 4564 13688 4616
rect 21180 4564 21232 4616
rect 12348 4496 12400 4548
rect 9312 4471 9364 4480
rect 9312 4437 9321 4471
rect 9321 4437 9355 4471
rect 9355 4437 9364 4471
rect 9312 4428 9364 4437
rect 14832 4496 14884 4548
rect 14648 4471 14700 4480
rect 14648 4437 14657 4471
rect 14657 4437 14691 4471
rect 14691 4437 14700 4471
rect 14648 4428 14700 4437
rect 16212 4496 16264 4548
rect 16672 4496 16724 4548
rect 21456 4496 21508 4548
rect 21824 4632 21876 4684
rect 23848 4768 23900 4820
rect 24768 4768 24820 4820
rect 26240 4768 26292 4820
rect 27712 4811 27764 4820
rect 27712 4777 27721 4811
rect 27721 4777 27755 4811
rect 27755 4777 27764 4811
rect 27712 4768 27764 4777
rect 28632 4768 28684 4820
rect 33048 4811 33100 4820
rect 33048 4777 33057 4811
rect 33057 4777 33091 4811
rect 33091 4777 33100 4811
rect 33048 4768 33100 4777
rect 38292 4811 38344 4820
rect 38292 4777 38301 4811
rect 38301 4777 38335 4811
rect 38335 4777 38344 4811
rect 38292 4768 38344 4777
rect 27160 4700 27212 4752
rect 23480 4564 23532 4616
rect 27068 4607 27120 4616
rect 27068 4573 27077 4607
rect 27077 4573 27111 4607
rect 27111 4573 27120 4607
rect 27068 4564 27120 4573
rect 27436 4564 27488 4616
rect 28172 4564 28224 4616
rect 28448 4607 28500 4616
rect 28448 4573 28457 4607
rect 28457 4573 28491 4607
rect 28491 4573 28500 4607
rect 28448 4564 28500 4573
rect 29184 4607 29236 4616
rect 29184 4573 29193 4607
rect 29193 4573 29227 4607
rect 29227 4573 29236 4607
rect 29184 4564 29236 4573
rect 31208 4564 31260 4616
rect 31852 4564 31904 4616
rect 33048 4564 33100 4616
rect 22100 4428 22152 4480
rect 23112 4496 23164 4548
rect 23204 4496 23256 4548
rect 25596 4496 25648 4548
rect 26332 4496 26384 4548
rect 26976 4428 27028 4480
rect 27068 4428 27120 4480
rect 28448 4428 28500 4480
rect 38016 4632 38068 4684
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 10048 4267 10100 4276
rect 10048 4233 10057 4267
rect 10057 4233 10091 4267
rect 10091 4233 10100 4267
rect 10048 4224 10100 4233
rect 11060 4267 11112 4276
rect 11060 4233 11069 4267
rect 11069 4233 11103 4267
rect 11103 4233 11112 4267
rect 11060 4224 11112 4233
rect 12532 4224 12584 4276
rect 20536 4224 20588 4276
rect 20628 4224 20680 4276
rect 21456 4224 21508 4276
rect 26424 4224 26476 4276
rect 26976 4224 27028 4276
rect 30380 4224 30432 4276
rect 13820 4156 13872 4208
rect 16212 4156 16264 4208
rect 16304 4199 16356 4208
rect 16304 4165 16313 4199
rect 16313 4165 16347 4199
rect 16347 4165 16356 4199
rect 16304 4156 16356 4165
rect 16488 4156 16540 4208
rect 19156 4156 19208 4208
rect 22192 4156 22244 4208
rect 24400 4156 24452 4208
rect 24492 4199 24544 4208
rect 24492 4165 24501 4199
rect 24501 4165 24535 4199
rect 24535 4165 24544 4199
rect 24492 4156 24544 4165
rect 28816 4156 28868 4208
rect 16856 4131 16908 4140
rect 16856 4097 16865 4131
rect 16865 4097 16899 4131
rect 16899 4097 16908 4131
rect 16856 4088 16908 4097
rect 14556 4063 14608 4072
rect 8024 3884 8076 3936
rect 9312 3884 9364 3936
rect 12072 3884 12124 3936
rect 14556 4029 14565 4063
rect 14565 4029 14599 4063
rect 14599 4029 14608 4063
rect 14556 4020 14608 4029
rect 17132 4063 17184 4072
rect 17132 4029 17141 4063
rect 17141 4029 17175 4063
rect 17175 4029 17184 4063
rect 17132 4020 17184 4029
rect 17224 4020 17276 4072
rect 17868 4020 17920 4072
rect 18880 4063 18932 4072
rect 14556 3884 14608 3936
rect 14740 3884 14792 3936
rect 18512 3952 18564 4004
rect 18880 4029 18889 4063
rect 18889 4029 18923 4063
rect 18923 4029 18932 4063
rect 18880 4020 18932 4029
rect 18972 4020 19024 4072
rect 21272 4088 21324 4140
rect 23848 4088 23900 4140
rect 25780 4088 25832 4140
rect 27988 4088 28040 4140
rect 28172 4088 28224 4140
rect 29000 4088 29052 4140
rect 29092 4088 29144 4140
rect 30012 4156 30064 4208
rect 29828 4088 29880 4140
rect 30288 4088 30340 4140
rect 30564 4088 30616 4140
rect 31208 4131 31260 4140
rect 31208 4097 31217 4131
rect 31217 4097 31251 4131
rect 31251 4097 31260 4131
rect 31208 4088 31260 4097
rect 33048 4088 33100 4140
rect 20352 4020 20404 4072
rect 20812 4020 20864 4072
rect 22100 4020 22152 4072
rect 23480 4063 23532 4072
rect 23480 4029 23489 4063
rect 23489 4029 23523 4063
rect 23523 4029 23532 4063
rect 23480 4020 23532 4029
rect 15660 3884 15712 3936
rect 15936 3884 15988 3936
rect 16948 3884 17000 3936
rect 18604 3884 18656 3936
rect 19892 3952 19944 4004
rect 22376 3952 22428 4004
rect 19340 3884 19392 3936
rect 20352 3884 20404 3936
rect 26332 4020 26384 4072
rect 26424 4020 26476 4072
rect 32496 4063 32548 4072
rect 32496 4029 32505 4063
rect 32505 4029 32539 4063
rect 32539 4029 32548 4063
rect 32496 4020 32548 4029
rect 26516 3995 26568 4004
rect 26516 3961 26525 3995
rect 26525 3961 26559 3995
rect 26559 3961 26568 3995
rect 26516 3952 26568 3961
rect 27436 3952 27488 4004
rect 31116 3995 31168 4004
rect 31116 3961 31125 3995
rect 31125 3961 31159 3995
rect 31159 3961 31168 3995
rect 31116 3952 31168 3961
rect 31760 3952 31812 4004
rect 38016 3952 38068 4004
rect 24584 3884 24636 3936
rect 28172 3927 28224 3936
rect 28172 3893 28181 3927
rect 28181 3893 28215 3927
rect 28215 3893 28224 3927
rect 28172 3884 28224 3893
rect 28448 3884 28500 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 12440 3680 12492 3732
rect 12624 3680 12676 3732
rect 17132 3680 17184 3732
rect 17224 3680 17276 3732
rect 23296 3680 23348 3732
rect 28172 3680 28224 3732
rect 28724 3680 28776 3732
rect 30380 3680 30432 3732
rect 34796 3680 34848 3732
rect 4436 3612 4488 3664
rect 8116 3612 8168 3664
rect 11980 3612 12032 3664
rect 13268 3612 13320 3664
rect 14648 3612 14700 3664
rect 8576 3587 8628 3596
rect 8576 3553 8585 3587
rect 8585 3553 8619 3587
rect 8619 3553 8628 3587
rect 8576 3544 8628 3553
rect 11888 3544 11940 3596
rect 12256 3587 12308 3596
rect 12256 3553 12265 3587
rect 12265 3553 12299 3587
rect 12299 3553 12308 3587
rect 12256 3544 12308 3553
rect 12716 3544 12768 3596
rect 18788 3612 18840 3664
rect 20352 3612 20404 3664
rect 23756 3612 23808 3664
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 8208 3476 8260 3528
rect 11796 3476 11848 3528
rect 8576 3408 8628 3460
rect 13360 3476 13412 3528
rect 7472 3383 7524 3392
rect 7472 3349 7481 3383
rect 7481 3349 7515 3383
rect 7515 3349 7524 3383
rect 7472 3340 7524 3349
rect 8024 3383 8076 3392
rect 8024 3349 8033 3383
rect 8033 3349 8067 3383
rect 8067 3349 8076 3383
rect 8024 3340 8076 3349
rect 12348 3408 12400 3460
rect 15016 3544 15068 3596
rect 14556 3476 14608 3528
rect 15200 3408 15252 3460
rect 16212 3408 16264 3460
rect 17132 3544 17184 3596
rect 19892 3544 19944 3596
rect 20628 3544 20680 3596
rect 23848 3544 23900 3596
rect 26424 3612 26476 3664
rect 26608 3612 26660 3664
rect 31760 3612 31812 3664
rect 37924 3612 37976 3664
rect 25504 3544 25556 3596
rect 30012 3544 30064 3596
rect 32956 3587 33008 3596
rect 14832 3340 14884 3392
rect 17316 3340 17368 3392
rect 17500 3340 17552 3392
rect 20444 3519 20496 3528
rect 20444 3485 20453 3519
rect 20453 3485 20487 3519
rect 20487 3485 20496 3519
rect 20444 3476 20496 3485
rect 23204 3476 23256 3528
rect 23940 3476 23992 3528
rect 26792 3519 26844 3528
rect 26792 3485 26801 3519
rect 26801 3485 26835 3519
rect 26835 3485 26844 3519
rect 26792 3476 26844 3485
rect 27344 3476 27396 3528
rect 27528 3519 27580 3528
rect 27528 3485 27537 3519
rect 27537 3485 27571 3519
rect 27571 3485 27580 3519
rect 27528 3476 27580 3485
rect 28080 3476 28132 3528
rect 18604 3408 18656 3460
rect 18972 3408 19024 3460
rect 21180 3408 21232 3460
rect 21364 3408 21416 3460
rect 22928 3408 22980 3460
rect 28448 3408 28500 3460
rect 28816 3476 28868 3528
rect 29920 3519 29972 3528
rect 29920 3485 29929 3519
rect 29929 3485 29963 3519
rect 29963 3485 29972 3519
rect 29920 3476 29972 3485
rect 30288 3476 30340 3528
rect 31024 3476 31076 3528
rect 32956 3553 32965 3587
rect 32965 3553 32999 3587
rect 32999 3553 33008 3587
rect 32956 3544 33008 3553
rect 31852 3519 31904 3528
rect 31300 3408 31352 3460
rect 31852 3485 31861 3519
rect 31861 3485 31895 3519
rect 31895 3485 31904 3519
rect 31852 3476 31904 3485
rect 32496 3519 32548 3528
rect 32496 3485 32505 3519
rect 32505 3485 32539 3519
rect 32539 3485 32548 3519
rect 32496 3476 32548 3485
rect 39304 3408 39356 3460
rect 18696 3340 18748 3392
rect 21916 3340 21968 3392
rect 28264 3340 28316 3392
rect 30472 3383 30524 3392
rect 30472 3349 30481 3383
rect 30481 3349 30515 3383
rect 30515 3349 30524 3383
rect 30472 3340 30524 3349
rect 31760 3383 31812 3392
rect 31760 3349 31769 3383
rect 31769 3349 31803 3383
rect 31803 3349 31812 3383
rect 31760 3340 31812 3349
rect 33600 3383 33652 3392
rect 33600 3349 33609 3383
rect 33609 3349 33643 3383
rect 33643 3349 33652 3383
rect 33600 3340 33652 3349
rect 34060 3383 34112 3392
rect 34060 3349 34069 3383
rect 34069 3349 34103 3383
rect 34103 3349 34112 3383
rect 34060 3340 34112 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2872 3136 2924 3188
rect 3332 3179 3384 3188
rect 3332 3145 3341 3179
rect 3341 3145 3375 3179
rect 3375 3145 3384 3179
rect 3332 3136 3384 3145
rect 11152 3136 11204 3188
rect 12164 3136 12216 3188
rect 12256 3136 12308 3188
rect 4436 3043 4488 3052
rect 4436 3009 4445 3043
rect 4445 3009 4479 3043
rect 4479 3009 4488 3043
rect 4436 3000 4488 3009
rect 10048 3068 10100 3120
rect 10324 3111 10376 3120
rect 10324 3077 10333 3111
rect 10333 3077 10367 3111
rect 10367 3077 10376 3111
rect 10324 3068 10376 3077
rect 11612 3068 11664 3120
rect 12808 3136 12860 3188
rect 12900 3068 12952 3120
rect 13912 3068 13964 3120
rect 7472 3000 7524 3052
rect 8944 2932 8996 2984
rect 10968 3000 11020 3052
rect 12348 3043 12400 3052
rect 12348 3009 12357 3043
rect 12357 3009 12391 3043
rect 12391 3009 12400 3043
rect 12348 3000 12400 3009
rect 13728 3000 13780 3052
rect 12716 2932 12768 2984
rect 12992 2932 13044 2984
rect 14096 2975 14148 2984
rect 9864 2864 9916 2916
rect 10048 2864 10100 2916
rect 10968 2864 11020 2916
rect 11152 2864 11204 2916
rect 1676 2839 1728 2848
rect 1676 2805 1685 2839
rect 1685 2805 1719 2839
rect 1719 2805 1728 2839
rect 1676 2796 1728 2805
rect 4620 2839 4672 2848
rect 4620 2805 4629 2839
rect 4629 2805 4663 2839
rect 4663 2805 4672 2839
rect 4620 2796 4672 2805
rect 8024 2796 8076 2848
rect 8944 2796 8996 2848
rect 10876 2796 10928 2848
rect 11612 2796 11664 2848
rect 13636 2796 13688 2848
rect 14096 2941 14105 2975
rect 14105 2941 14139 2975
rect 14139 2941 14148 2975
rect 14096 2932 14148 2941
rect 17132 3136 17184 3188
rect 14556 2975 14608 2984
rect 14556 2941 14565 2975
rect 14565 2941 14599 2975
rect 14599 2941 14608 2975
rect 14556 2932 14608 2941
rect 16948 2932 17000 2984
rect 16120 2796 16172 2848
rect 19340 3136 19392 3188
rect 19800 3136 19852 3188
rect 18788 3068 18840 3120
rect 19616 3068 19668 3120
rect 22468 3068 22520 3120
rect 23296 3068 23348 3120
rect 23848 3068 23900 3120
rect 19340 3000 19392 3052
rect 25504 3068 25556 3120
rect 26240 3043 26292 3052
rect 26240 3009 26249 3043
rect 26249 3009 26283 3043
rect 26283 3009 26292 3043
rect 27436 3043 27488 3052
rect 26240 3000 26292 3009
rect 27436 3009 27445 3043
rect 27445 3009 27479 3043
rect 27479 3009 27488 3043
rect 27436 3000 27488 3009
rect 28448 3068 28500 3120
rect 28632 3068 28684 3120
rect 28540 3043 28592 3052
rect 28540 3009 28549 3043
rect 28549 3009 28583 3043
rect 28583 3009 28592 3043
rect 28540 3000 28592 3009
rect 17592 2932 17644 2984
rect 19156 2932 19208 2984
rect 20720 2864 20772 2916
rect 19800 2796 19852 2848
rect 20444 2796 20496 2848
rect 23388 2932 23440 2984
rect 23756 2975 23808 2984
rect 23756 2941 23765 2975
rect 23765 2941 23799 2975
rect 23799 2941 23808 2975
rect 24492 2975 24544 2984
rect 23756 2932 23808 2941
rect 24492 2941 24501 2975
rect 24501 2941 24535 2975
rect 24535 2941 24544 2975
rect 24492 2932 24544 2941
rect 25228 2932 25280 2984
rect 28632 2932 28684 2984
rect 24860 2864 24912 2916
rect 28908 3000 28960 3052
rect 29276 3000 29328 3052
rect 29736 3000 29788 3052
rect 30288 3000 30340 3052
rect 32496 3043 32548 3052
rect 32496 3009 32505 3043
rect 32505 3009 32539 3043
rect 32539 3009 32548 3043
rect 32496 3000 32548 3009
rect 33140 3000 33192 3052
rect 38016 3043 38068 3052
rect 38016 3009 38025 3043
rect 38025 3009 38059 3043
rect 38059 3009 38068 3043
rect 38016 3000 38068 3009
rect 31024 2932 31076 2984
rect 34336 2932 34388 2984
rect 30840 2864 30892 2916
rect 36636 2864 36688 2916
rect 27068 2796 27120 2848
rect 27896 2839 27948 2848
rect 27896 2805 27905 2839
rect 27905 2805 27939 2839
rect 27939 2805 27948 2839
rect 27896 2796 27948 2805
rect 28908 2796 28960 2848
rect 29276 2839 29328 2848
rect 29276 2805 29285 2839
rect 29285 2805 29319 2839
rect 29319 2805 29328 2839
rect 29276 2796 29328 2805
rect 29920 2839 29972 2848
rect 29920 2805 29929 2839
rect 29929 2805 29963 2839
rect 29963 2805 29972 2839
rect 29920 2796 29972 2805
rect 30564 2839 30616 2848
rect 30564 2805 30573 2839
rect 30573 2805 30607 2839
rect 30607 2805 30616 2839
rect 30564 2796 30616 2805
rect 31208 2839 31260 2848
rect 31208 2805 31217 2839
rect 31217 2805 31251 2839
rect 31251 2805 31260 2839
rect 31208 2796 31260 2805
rect 32312 2796 32364 2848
rect 35440 2796 35492 2848
rect 38200 2839 38252 2848
rect 38200 2805 38209 2839
rect 38209 2805 38243 2839
rect 38243 2805 38252 2839
rect 38200 2796 38252 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 2136 2592 2188 2644
rect 8024 2635 8076 2644
rect 8024 2601 8033 2635
rect 8033 2601 8067 2635
rect 8067 2601 8076 2635
rect 8024 2592 8076 2601
rect 10048 2635 10100 2644
rect 10048 2601 10057 2635
rect 10057 2601 10091 2635
rect 10091 2601 10100 2635
rect 10048 2592 10100 2601
rect 11704 2592 11756 2644
rect 13268 2592 13320 2644
rect 20 2524 72 2576
rect 3332 2524 3384 2576
rect 10784 2524 10836 2576
rect 12348 2524 12400 2576
rect 2872 2388 2924 2440
rect 3240 2388 3292 2440
rect 7196 2456 7248 2508
rect 14556 2499 14608 2508
rect 14556 2465 14565 2499
rect 14565 2465 14599 2499
rect 14599 2465 14608 2499
rect 17132 2499 17184 2508
rect 14556 2456 14608 2465
rect 17132 2465 17141 2499
rect 17141 2465 17175 2499
rect 17175 2465 17184 2499
rect 17132 2456 17184 2465
rect 8208 2388 8260 2440
rect 9864 2431 9916 2440
rect 9864 2397 9873 2431
rect 9873 2397 9907 2431
rect 9907 2397 9916 2431
rect 9864 2388 9916 2397
rect 11152 2388 11204 2440
rect 12348 2388 12400 2440
rect 22008 2592 22060 2644
rect 29552 2592 29604 2644
rect 31300 2592 31352 2644
rect 33600 2592 33652 2644
rect 23480 2524 23532 2576
rect 26516 2524 26568 2576
rect 29276 2524 29328 2576
rect 30932 2524 30984 2576
rect 18604 2456 18656 2508
rect 24400 2456 24452 2508
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 25044 2456 25096 2508
rect 26332 2499 26384 2508
rect 26332 2465 26341 2499
rect 26341 2465 26375 2499
rect 26375 2465 26384 2499
rect 26332 2456 26384 2465
rect 29828 2499 29880 2508
rect 29828 2465 29837 2499
rect 29837 2465 29871 2499
rect 29871 2465 29880 2499
rect 29828 2456 29880 2465
rect 8392 2320 8444 2372
rect 13544 2320 13596 2372
rect 17316 2320 17368 2372
rect 17684 2320 17736 2372
rect 19984 2320 20036 2372
rect 21364 2320 21416 2372
rect 21456 2363 21508 2372
rect 21456 2329 21465 2363
rect 21465 2329 21499 2363
rect 21499 2329 21508 2363
rect 21456 2320 21508 2329
rect 1308 2252 1360 2304
rect 4528 2252 4580 2304
rect 6460 2252 6512 2304
rect 8576 2295 8628 2304
rect 8576 2261 8585 2295
rect 8585 2261 8619 2295
rect 8619 2261 8628 2295
rect 8576 2252 8628 2261
rect 9312 2295 9364 2304
rect 9312 2261 9321 2295
rect 9321 2261 9355 2295
rect 9355 2261 9364 2295
rect 9312 2252 9364 2261
rect 11336 2252 11388 2304
rect 18420 2252 18472 2304
rect 19892 2252 19944 2304
rect 27896 2388 27948 2440
rect 27988 2388 28040 2440
rect 28816 2431 28868 2440
rect 28816 2397 28825 2431
rect 28825 2397 28859 2431
rect 28859 2397 28868 2431
rect 28816 2388 28868 2397
rect 29736 2431 29788 2440
rect 29736 2397 29745 2431
rect 29745 2397 29779 2431
rect 29779 2397 29788 2431
rect 29736 2388 29788 2397
rect 25596 2320 25648 2372
rect 26424 2320 26476 2372
rect 28080 2363 28132 2372
rect 28080 2329 28089 2363
rect 28089 2329 28123 2363
rect 28123 2329 28132 2363
rect 28080 2320 28132 2329
rect 23756 2295 23808 2304
rect 23756 2261 23765 2295
rect 23765 2261 23799 2295
rect 23799 2261 23808 2295
rect 23756 2252 23808 2261
rect 23848 2252 23900 2304
rect 28724 2295 28776 2304
rect 28724 2261 28733 2295
rect 28733 2261 28767 2295
rect 28767 2261 28776 2295
rect 28724 2252 28776 2261
rect 30288 2252 30340 2304
rect 31300 2431 31352 2440
rect 31300 2397 31309 2431
rect 31309 2397 31343 2431
rect 31343 2397 31352 2431
rect 31300 2388 31352 2397
rect 34060 2456 34112 2508
rect 32312 2431 32364 2440
rect 32312 2397 32321 2431
rect 32321 2397 32355 2431
rect 32355 2397 32364 2431
rect 32312 2388 32364 2397
rect 32220 2320 32272 2372
rect 34336 2388 34388 2440
rect 34796 2388 34848 2440
rect 36636 2431 36688 2440
rect 36636 2397 36645 2431
rect 36645 2397 36679 2431
rect 36679 2397 36688 2431
rect 36636 2388 36688 2397
rect 37464 2431 37516 2440
rect 37464 2397 37473 2431
rect 37473 2397 37507 2431
rect 37507 2397 37516 2431
rect 37464 2388 37516 2397
rect 35440 2320 35492 2372
rect 33140 2252 33192 2304
rect 33600 2295 33652 2304
rect 33600 2261 33609 2295
rect 33609 2261 33643 2295
rect 33643 2261 33652 2295
rect 33600 2252 33652 2261
rect 34152 2252 34204 2304
rect 37188 2252 37240 2304
rect 37372 2252 37424 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 17316 2048 17368 2100
rect 8576 1980 8628 2032
rect 18604 1980 18656 2032
rect 18880 1980 18932 2032
rect 21456 1980 21508 2032
rect 22192 2048 22244 2100
rect 28724 2048 28776 2100
rect 28908 2048 28960 2100
rect 37464 2048 37516 2100
rect 31208 1980 31260 2032
rect 16212 1912 16264 1964
rect 31760 1912 31812 1964
rect 13360 1844 13412 1896
rect 25504 1844 25556 1896
rect 25596 1844 25648 1896
rect 30564 1844 30616 1896
rect 21364 1776 21416 1828
rect 33600 1776 33652 1828
rect 25136 1708 25188 1760
rect 28080 1708 28132 1760
rect 29000 1708 29052 1760
rect 32312 1708 32364 1760
rect 9312 1640 9364 1692
rect 26792 1640 26844 1692
rect 25504 1572 25556 1624
rect 30472 1572 30524 1624
<< metal2 >>
rect 1306 39200 1362 39800
rect 2594 39200 2650 39800
rect 2962 39536 3018 39545
rect 2962 39471 3018 39480
rect 1320 37126 1348 39200
rect 2320 37256 2372 37262
rect 2320 37198 2372 37204
rect 2608 37210 2636 39200
rect 2870 37496 2926 37505
rect 2870 37431 2926 37440
rect 1308 37120 1360 37126
rect 1308 37062 1360 37068
rect 1860 36168 1912 36174
rect 1674 36136 1730 36145
rect 1860 36110 1912 36116
rect 1674 36071 1730 36080
rect 1688 36038 1716 36071
rect 1676 36032 1728 36038
rect 1676 35974 1728 35980
rect 1872 35834 1900 36110
rect 1860 35828 1912 35834
rect 1860 35770 1912 35776
rect 2228 34536 2280 34542
rect 2228 34478 2280 34484
rect 1676 34400 1728 34406
rect 1676 34342 1728 34348
rect 1688 34105 1716 34342
rect 1674 34096 1730 34105
rect 1674 34031 1730 34040
rect 1584 32428 1636 32434
rect 1584 32370 1636 32376
rect 1596 32065 1624 32370
rect 1582 32056 1638 32065
rect 1582 31991 1584 32000
rect 1636 31991 1638 32000
rect 1584 31962 1636 31968
rect 1674 30696 1730 30705
rect 1674 30631 1676 30640
rect 1728 30631 1730 30640
rect 1676 30602 1728 30608
rect 1688 30394 1716 30602
rect 1768 30592 1820 30598
rect 1768 30534 1820 30540
rect 1676 30388 1728 30394
rect 1676 30330 1728 30336
rect 1584 29096 1636 29102
rect 1584 29038 1636 29044
rect 1596 28694 1624 29038
rect 1584 28688 1636 28694
rect 1582 28656 1584 28665
rect 1636 28656 1638 28665
rect 1582 28591 1638 28600
rect 1676 26784 1728 26790
rect 1676 26726 1728 26732
rect 1688 26625 1716 26726
rect 1674 26616 1730 26625
rect 1674 26551 1730 26560
rect 1584 25288 1636 25294
rect 1582 25256 1584 25265
rect 1636 25256 1638 25265
rect 1582 25191 1638 25200
rect 1596 24954 1624 25191
rect 1584 24948 1636 24954
rect 1584 24890 1636 24896
rect 1780 23882 1808 30534
rect 2044 25288 2096 25294
rect 2044 25230 2096 25236
rect 1780 23854 1992 23882
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 1676 23520 1728 23526
rect 1676 23462 1728 23468
rect 1688 23225 1716 23462
rect 1674 23216 1730 23225
rect 1674 23151 1730 23160
rect 1768 21548 1820 21554
rect 1768 21490 1820 21496
rect 1676 21344 1728 21350
rect 1676 21286 1728 21292
rect 1688 21185 1716 21286
rect 1674 21176 1730 21185
rect 1780 21146 1808 21490
rect 1674 21111 1730 21120
rect 1768 21140 1820 21146
rect 1768 21082 1820 21088
rect 1674 19816 1730 19825
rect 1674 19751 1730 19760
rect 1688 19718 1716 19751
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1872 19514 1900 23666
rect 1964 19922 1992 23854
rect 2056 20942 2084 25230
rect 2044 20936 2096 20942
rect 2044 20878 2096 20884
rect 1952 19916 2004 19922
rect 1952 19858 2004 19864
rect 1860 19508 1912 19514
rect 1860 19450 1912 19456
rect 2056 19446 2084 20878
rect 2044 19440 2096 19446
rect 2044 19382 2096 19388
rect 2136 19372 2188 19378
rect 2136 19314 2188 19320
rect 1768 18828 1820 18834
rect 1768 18770 1820 18776
rect 1780 18426 1808 18770
rect 1768 18420 1820 18426
rect 1768 18362 1820 18368
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 1596 17814 1624 18226
rect 1584 17808 1636 17814
rect 1582 17776 1584 17785
rect 1636 17776 1638 17785
rect 1582 17711 1638 17720
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1688 15745 1716 15846
rect 1674 15736 1730 15745
rect 1674 15671 1730 15680
rect 1674 14376 1730 14385
rect 1674 14311 1730 14320
rect 1688 14278 1716 14311
rect 1676 14272 1728 14278
rect 1676 14214 1728 14220
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1688 12345 1716 12582
rect 1674 12336 1730 12345
rect 1674 12271 1730 12280
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1596 10305 1624 10610
rect 1582 10296 1638 10305
rect 1582 10231 1584 10240
rect 1636 10231 1638 10240
rect 1584 10202 1636 10208
rect 1584 8968 1636 8974
rect 1582 8936 1584 8945
rect 1636 8936 1638 8945
rect 1582 8871 1638 8880
rect 1596 8634 1624 8871
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1872 7478 1900 12038
rect 1860 7472 1912 7478
rect 1860 7414 1912 7420
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1596 7002 1624 7346
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1596 6905 1624 6938
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1688 4865 1716 4966
rect 1674 4856 1730 4865
rect 1674 4791 1730 4800
rect 1584 3528 1636 3534
rect 1582 3496 1584 3505
rect 1636 3496 1638 3505
rect 1582 3431 1638 3440
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 20 2576 72 2582
rect 20 2518 72 2524
rect 32 800 60 2518
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 1320 800 1348 2246
rect 1688 1465 1716 2790
rect 2148 2650 2176 19314
rect 2240 16794 2268 34478
rect 2332 20058 2360 37198
rect 2608 37182 2820 37210
rect 2792 37126 2820 37182
rect 2780 37120 2832 37126
rect 2780 37062 2832 37068
rect 2884 36854 2912 37431
rect 2872 36848 2924 36854
rect 2872 36790 2924 36796
rect 2504 36576 2556 36582
rect 2504 36518 2556 36524
rect 2320 20052 2372 20058
rect 2320 19994 2372 20000
rect 2516 19514 2544 36518
rect 2884 36378 2912 36790
rect 2976 36786 3004 39471
rect 4526 39200 4582 39800
rect 6458 39200 6514 39800
rect 7746 39200 7802 39800
rect 9678 39200 9734 39800
rect 11610 39200 11666 39800
rect 12898 39200 12954 39800
rect 14830 39200 14886 39800
rect 16762 39200 16818 39800
rect 18050 39200 18106 39800
rect 19982 39200 20038 39800
rect 21914 39200 21970 39800
rect 23202 39200 23258 39800
rect 25134 39200 25190 39800
rect 27066 39200 27122 39800
rect 28354 39200 28410 39800
rect 30286 39200 30342 39800
rect 32218 39200 32274 39800
rect 33506 39200 33562 39800
rect 35438 39200 35494 39800
rect 37370 39200 37426 39800
rect 38658 39200 38714 39800
rect 4540 37754 4568 39200
rect 4540 37726 4660 37754
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4632 37126 4660 37726
rect 5448 37256 5500 37262
rect 5448 37198 5500 37204
rect 5460 37126 5488 37198
rect 6472 37126 6500 39200
rect 7760 37262 7788 39200
rect 7288 37256 7340 37262
rect 7288 37198 7340 37204
rect 7748 37256 7800 37262
rect 7748 37198 7800 37204
rect 6736 37188 6788 37194
rect 6736 37130 6788 37136
rect 4620 37120 4672 37126
rect 4620 37062 4672 37068
rect 5448 37120 5500 37126
rect 5448 37062 5500 37068
rect 6460 37120 6512 37126
rect 6460 37062 6512 37068
rect 5460 36922 5488 37062
rect 5448 36916 5500 36922
rect 5448 36858 5500 36864
rect 2964 36780 3016 36786
rect 2964 36722 3016 36728
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 2872 36372 2924 36378
rect 2872 36314 2924 36320
rect 3424 35488 3476 35494
rect 3424 35430 3476 35436
rect 2596 19848 2648 19854
rect 2596 19790 2648 19796
rect 2504 19508 2556 19514
rect 2504 19450 2556 19456
rect 2228 16788 2280 16794
rect 2228 16730 2280 16736
rect 2608 12102 2636 19790
rect 3436 14618 3464 35430
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 6748 34202 6776 37130
rect 7300 36582 7328 37198
rect 9692 37126 9720 39200
rect 11624 37126 11652 39200
rect 12072 37256 12124 37262
rect 12072 37198 12124 37204
rect 8024 37120 8076 37126
rect 8024 37062 8076 37068
rect 9680 37120 9732 37126
rect 9680 37062 9732 37068
rect 11612 37120 11664 37126
rect 11612 37062 11664 37068
rect 7288 36576 7340 36582
rect 7288 36518 7340 36524
rect 6736 34196 6788 34202
rect 6736 34138 6788 34144
rect 7104 33992 7156 33998
rect 7104 33934 7156 33940
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 6552 26988 6604 26994
rect 6552 26930 6604 26936
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 6564 21690 6592 26930
rect 7116 24138 7144 33934
rect 7104 24132 7156 24138
rect 7104 24074 7156 24080
rect 6552 21684 6604 21690
rect 6552 21626 6604 21632
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4620 19780 4672 19786
rect 4620 19722 4672 19728
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4632 18426 4660 19722
rect 4620 18420 4672 18426
rect 4620 18362 4672 18368
rect 8036 18086 8064 37062
rect 10048 21344 10100 21350
rect 10048 21286 10100 21292
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 8024 18080 8076 18086
rect 8024 18022 8076 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 8208 16516 8260 16522
rect 8208 16458 8260 16464
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 8128 15706 8156 16050
rect 8116 15700 8168 15706
rect 8116 15642 8168 15648
rect 8220 15502 8248 16458
rect 9692 15706 9720 19110
rect 9772 15972 9824 15978
rect 9772 15914 9824 15920
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9692 15502 9720 15642
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9312 14884 9364 14890
rect 9312 14826 9364 14832
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 9324 14414 9352 14826
rect 9404 14476 9456 14482
rect 9404 14418 9456 14424
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 5552 12442 5580 12786
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 7760 12170 7788 12786
rect 7748 12164 7800 12170
rect 7748 12106 7800 12112
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 2872 11076 2924 11082
rect 2872 11018 2924 11024
rect 2780 8356 2832 8362
rect 2780 8298 2832 8304
rect 2792 5234 2820 8298
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2884 3194 2912 11018
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3344 3194 3372 7822
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4436 3664 4488 3670
rect 4436 3606 4488 3612
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 2136 2644 2188 2650
rect 2136 2586 2188 2592
rect 2884 2446 2912 3130
rect 3344 2582 3372 3130
rect 4448 3058 4476 3606
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4618 2952 4674 2961
rect 4618 2887 4674 2896
rect 4632 2854 4660 2887
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 3332 2576 3384 2582
rect 3332 2518 3384 2524
rect 7208 2514 7236 9386
rect 7300 9042 7328 11494
rect 7852 11082 7880 13806
rect 7932 13728 7984 13734
rect 7932 13670 7984 13676
rect 7944 12986 7972 13670
rect 9128 13456 9180 13462
rect 9128 13398 9180 13404
rect 8852 13320 8904 13326
rect 8852 13262 8904 13268
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 8864 12434 8892 13262
rect 9140 12986 9168 13398
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 8864 12406 8984 12434
rect 8760 12164 8812 12170
rect 8760 12106 8812 12112
rect 8116 11756 8168 11762
rect 8116 11698 8168 11704
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 8128 10470 8156 11698
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 8036 3398 8064 3878
rect 8128 3670 8156 10406
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 8588 3602 8616 11018
rect 8772 10810 8800 12106
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 8772 10266 8800 10746
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8864 10538 8892 10610
rect 8852 10532 8904 10538
rect 8852 10474 8904 10480
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8772 10062 8800 10202
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8864 9874 8892 10474
rect 8772 9846 8892 9874
rect 8772 9382 8800 9846
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8772 5370 8800 9318
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 7484 3058 7512 3334
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 8036 2854 8064 3334
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 8036 2650 8064 2790
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 8220 2446 8248 3470
rect 8576 3460 8628 3466
rect 8576 3402 8628 3408
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 1674 1456 1730 1465
rect 1674 1391 1730 1400
rect 3252 800 3280 2382
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 4540 800 4568 2246
rect 6472 800 6500 2246
rect 8404 800 8432 2314
rect 8588 2310 8616 3402
rect 8956 2990 8984 12406
rect 9048 12238 9076 12786
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 9048 11898 9076 12174
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 9048 10198 9076 11834
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9036 10192 9088 10198
rect 9036 10134 9088 10140
rect 9140 9722 9168 11494
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9232 10810 9260 10950
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 9324 9217 9352 14350
rect 9416 9926 9444 14418
rect 9784 14414 9812 15914
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9784 14006 9812 14350
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9876 13138 9904 13194
rect 9876 13110 9996 13138
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 9586 12336 9642 12345
rect 9586 12271 9642 12280
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 9508 11082 9536 12174
rect 9600 12170 9628 12271
rect 9588 12164 9640 12170
rect 9588 12106 9640 12112
rect 9496 11076 9548 11082
rect 9496 11018 9548 11024
rect 9692 10266 9720 12854
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9772 12368 9824 12374
rect 9772 12310 9824 12316
rect 9784 12209 9812 12310
rect 9770 12200 9826 12209
rect 9770 12135 9826 12144
rect 9876 11257 9904 12786
rect 9862 11248 9918 11257
rect 9862 11183 9918 11192
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9692 9654 9720 10202
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9310 9208 9366 9217
rect 9310 9143 9366 9152
rect 9692 6866 9720 9590
rect 9784 9178 9812 11018
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 9876 10130 9904 10950
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9784 8498 9812 9114
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9876 5574 9904 6054
rect 9968 5846 9996 13110
rect 10060 9042 10088 21286
rect 11520 19168 11572 19174
rect 11520 19110 11572 19116
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 10968 15564 11020 15570
rect 10968 15506 11020 15512
rect 10782 15056 10838 15065
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 10416 15020 10468 15026
rect 10980 15026 11008 15506
rect 11072 15162 11100 16186
rect 11164 16114 11192 18022
rect 11244 17604 11296 17610
rect 11244 17546 11296 17552
rect 11256 16454 11284 17546
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11152 15496 11204 15502
rect 11150 15464 11152 15473
rect 11256 15484 11284 16390
rect 11204 15464 11284 15484
rect 11206 15456 11284 15464
rect 11150 15399 11206 15408
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10782 14991 10838 15000
rect 10968 15020 11020 15026
rect 10416 14962 10468 14968
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10152 10985 10180 12378
rect 10138 10976 10194 10985
rect 10138 10911 10194 10920
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 10244 8090 10272 14962
rect 10324 14884 10376 14890
rect 10324 14826 10376 14832
rect 10336 14006 10364 14826
rect 10324 14000 10376 14006
rect 10324 13942 10376 13948
rect 10322 13832 10378 13841
rect 10322 13767 10378 13776
rect 10336 11898 10364 13767
rect 10428 12186 10456 14962
rect 10508 14408 10560 14414
rect 10506 14376 10508 14385
rect 10560 14376 10562 14385
rect 10506 14311 10562 14320
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10612 12322 10640 13126
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10704 12753 10732 12786
rect 10690 12744 10746 12753
rect 10690 12679 10746 12688
rect 10796 12646 10824 14991
rect 10968 14962 11020 14968
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 10876 13864 10928 13870
rect 11164 13818 11192 13874
rect 10876 13806 10928 13812
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10782 12472 10838 12481
rect 10782 12407 10784 12416
rect 10836 12407 10838 12416
rect 10784 12378 10836 12384
rect 10612 12294 10824 12322
rect 10692 12232 10744 12238
rect 10428 12158 10640 12186
rect 10692 12174 10744 12180
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10428 11558 10456 12038
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10520 11098 10548 11698
rect 10428 11082 10548 11098
rect 10324 11076 10376 11082
rect 10324 11018 10376 11024
rect 10416 11076 10548 11082
rect 10468 11070 10548 11076
rect 10416 11018 10468 11024
rect 10336 9654 10364 11018
rect 10612 10198 10640 12158
rect 10508 10192 10560 10198
rect 10508 10134 10560 10140
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 10520 10033 10548 10134
rect 10506 10024 10562 10033
rect 10506 9959 10562 9968
rect 10324 9648 10376 9654
rect 10324 9590 10376 9596
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10428 8922 10456 9318
rect 10428 8894 10548 8922
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10416 6180 10468 6186
rect 10416 6122 10468 6128
rect 10428 5914 10456 6122
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 9956 5840 10008 5846
rect 9956 5782 10008 5788
rect 10324 5840 10376 5846
rect 10324 5782 10376 5788
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 9876 5030 9904 5510
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9324 4486 9352 4966
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9324 3942 9352 4422
rect 10046 4312 10102 4321
rect 10046 4247 10048 4256
rect 10100 4247 10102 4256
rect 10048 4218 10100 4224
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 10336 3126 10364 5782
rect 10520 4758 10548 8894
rect 10612 7954 10640 10134
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 10704 6089 10732 12174
rect 10796 9382 10824 12294
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10888 9081 10916 13806
rect 10980 13790 11192 13818
rect 11256 13802 11284 13942
rect 11440 13938 11468 14758
rect 11428 13932 11480 13938
rect 11428 13874 11480 13880
rect 11244 13796 11296 13802
rect 10980 13530 11008 13790
rect 11244 13738 11296 13744
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 11058 13424 11114 13433
rect 11058 13359 11060 13368
rect 11112 13359 11114 13368
rect 11060 13330 11112 13336
rect 11256 13326 11284 13738
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10980 12850 11008 13126
rect 11152 12912 11204 12918
rect 11072 12860 11152 12866
rect 11072 12854 11204 12860
rect 11242 12880 11298 12889
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 11072 12838 11192 12854
rect 11072 11778 11100 12838
rect 11242 12815 11298 12824
rect 11256 12442 11284 12815
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11152 12368 11204 12374
rect 11440 12345 11468 13874
rect 11532 12918 11560 19110
rect 12084 16153 12112 37198
rect 12912 37126 12940 39200
rect 14844 37330 14872 39200
rect 16776 37482 16804 39200
rect 16684 37454 16804 37482
rect 18064 37466 18092 39200
rect 18052 37460 18104 37466
rect 16684 37330 16712 37454
rect 18052 37402 18104 37408
rect 14832 37324 14884 37330
rect 14832 37266 14884 37272
rect 16672 37324 16724 37330
rect 16672 37266 16724 37272
rect 16764 37324 16816 37330
rect 16764 37266 16816 37272
rect 13268 37256 13320 37262
rect 13268 37198 13320 37204
rect 13360 37256 13412 37262
rect 13360 37198 13412 37204
rect 13176 37188 13228 37194
rect 13176 37130 13228 37136
rect 12900 37120 12952 37126
rect 12900 37062 12952 37068
rect 12716 33516 12768 33522
rect 12716 33458 12768 33464
rect 12256 19508 12308 19514
rect 12256 19450 12308 19456
rect 12268 19378 12296 19450
rect 12256 19372 12308 19378
rect 12256 19314 12308 19320
rect 12728 19310 12756 33458
rect 12992 32224 13044 32230
rect 12992 32166 13044 32172
rect 13004 25498 13032 32166
rect 13188 28218 13216 37130
rect 13176 28212 13228 28218
rect 13176 28154 13228 28160
rect 13280 26042 13308 37198
rect 13372 36786 13400 37198
rect 13360 36780 13412 36786
rect 13360 36722 13412 36728
rect 13372 28558 13400 36722
rect 16304 36644 16356 36650
rect 16304 36586 16356 36592
rect 14740 30252 14792 30258
rect 14740 30194 14792 30200
rect 14752 30054 14780 30194
rect 14740 30048 14792 30054
rect 14740 29990 14792 29996
rect 14752 29102 14780 29990
rect 14740 29096 14792 29102
rect 14740 29038 14792 29044
rect 13360 28552 13412 28558
rect 13360 28494 13412 28500
rect 14280 28416 14332 28422
rect 14280 28358 14332 28364
rect 13268 26036 13320 26042
rect 13268 25978 13320 25984
rect 12992 25492 13044 25498
rect 12992 25434 13044 25440
rect 13004 25294 13032 25434
rect 12992 25288 13044 25294
rect 12992 25230 13044 25236
rect 12900 25152 12952 25158
rect 12900 25094 12952 25100
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 12808 17264 12860 17270
rect 12808 17206 12860 17212
rect 12624 16516 12676 16522
rect 12624 16458 12676 16464
rect 12070 16144 12126 16153
rect 12070 16079 12126 16088
rect 12636 15978 12664 16458
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12532 15972 12584 15978
rect 12532 15914 12584 15920
rect 12624 15972 12676 15978
rect 12624 15914 12676 15920
rect 12544 15881 12572 15914
rect 12530 15872 12586 15881
rect 12530 15807 12586 15816
rect 12728 15502 12756 16390
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 11796 15360 11848 15366
rect 11796 15302 11848 15308
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11624 12918 11652 14010
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11716 13462 11744 13670
rect 11704 13456 11756 13462
rect 11704 13398 11756 13404
rect 11808 13326 11836 15302
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 12072 14884 12124 14890
rect 12072 14826 12124 14832
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 11992 14521 12020 14554
rect 11978 14512 12034 14521
rect 11978 14447 12034 14456
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11900 14074 11928 14214
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11520 12912 11572 12918
rect 11520 12854 11572 12860
rect 11612 12912 11664 12918
rect 11612 12854 11664 12860
rect 11152 12310 11204 12316
rect 11426 12336 11482 12345
rect 11164 11898 11192 12310
rect 11426 12271 11482 12280
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11428 12164 11480 12170
rect 11256 12124 11428 12152
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 10980 11762 11100 11778
rect 10968 11756 11100 11762
rect 11020 11750 11100 11756
rect 11152 11756 11204 11762
rect 10968 11698 11020 11704
rect 11152 11698 11204 11704
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 11072 10554 11100 11562
rect 10980 10538 11100 10554
rect 10968 10532 11100 10538
rect 11020 10526 11100 10532
rect 10968 10474 11020 10480
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 11072 10266 11100 10406
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 10980 10062 11008 10202
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10874 9072 10930 9081
rect 10784 9036 10836 9042
rect 10874 9007 10930 9016
rect 10784 8978 10836 8984
rect 10690 6080 10746 6089
rect 10690 6015 10746 6024
rect 10508 4752 10560 4758
rect 10508 4694 10560 4700
rect 10048 3120 10100 3126
rect 10048 3062 10100 3068
rect 10324 3120 10376 3126
rect 10324 3062 10376 3068
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 8956 2854 8984 2926
rect 10060 2922 10088 3062
rect 9864 2916 9916 2922
rect 9864 2858 9916 2864
rect 10048 2916 10100 2922
rect 10048 2858 10100 2864
rect 8944 2848 8996 2854
rect 8944 2790 8996 2796
rect 9876 2446 9904 2858
rect 10060 2650 10088 2858
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 10796 2582 10824 8978
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 10980 8634 11008 8910
rect 11060 8900 11112 8906
rect 11060 8842 11112 8848
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 11072 8430 11100 8842
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 11072 7750 11100 8366
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 11072 7206 11100 7686
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11072 6662 11100 7142
rect 11164 7041 11192 11698
rect 11256 11626 11284 12124
rect 11428 12106 11480 12112
rect 11244 11620 11296 11626
rect 11244 11562 11296 11568
rect 11336 11620 11388 11626
rect 11336 11562 11388 11568
rect 11348 11150 11376 11562
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11336 11144 11388 11150
rect 11624 11121 11652 11222
rect 11336 11086 11388 11092
rect 11610 11112 11666 11121
rect 11428 11076 11480 11082
rect 11428 11018 11480 11024
rect 11520 11076 11572 11082
rect 11610 11047 11666 11056
rect 11520 11018 11572 11024
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 11256 10169 11284 10610
rect 11242 10160 11298 10169
rect 11242 10095 11298 10104
rect 11348 10062 11376 10610
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11244 9920 11296 9926
rect 11242 9888 11244 9897
rect 11296 9888 11298 9897
rect 11242 9823 11298 9832
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11256 8786 11284 9590
rect 11348 9178 11376 9998
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11256 8758 11376 8786
rect 11244 8560 11296 8566
rect 11242 8528 11244 8537
rect 11296 8528 11298 8537
rect 11242 8463 11298 8472
rect 11150 7032 11206 7041
rect 11150 6967 11206 6976
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11072 6118 11100 6598
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 11072 4826 11100 4966
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 11072 4690 11100 4762
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 11072 4282 11100 4626
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 10980 2922 11008 2994
rect 11164 2922 11192 3130
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 11152 2916 11204 2922
rect 11152 2858 11204 2864
rect 10876 2848 10928 2854
rect 10874 2816 10876 2825
rect 10928 2816 10930 2825
rect 10874 2751 10930 2760
rect 10784 2576 10836 2582
rect 10784 2518 10836 2524
rect 11164 2446 11192 2858
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 8576 2304 8628 2310
rect 8576 2246 8628 2252
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 8588 2038 8616 2246
rect 8576 2032 8628 2038
rect 8576 1974 8628 1980
rect 9324 1698 9352 2246
rect 9876 1986 9904 2382
rect 11348 2310 11376 8758
rect 11440 5658 11468 11018
rect 11532 10577 11560 11018
rect 11518 10568 11574 10577
rect 11518 10503 11574 10512
rect 11612 10532 11664 10538
rect 11532 9178 11560 10503
rect 11612 10474 11664 10480
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11440 5630 11560 5658
rect 11532 5574 11560 5630
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11532 5302 11560 5510
rect 11520 5296 11572 5302
rect 11520 5238 11572 5244
rect 11624 3126 11652 10474
rect 11716 6322 11744 12174
rect 11808 9178 11836 13126
rect 11992 12986 12020 14350
rect 12084 13326 12112 14826
rect 12176 14618 12204 14962
rect 12452 14958 12480 15302
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12164 14612 12216 14618
rect 12164 14554 12216 14560
rect 12256 14544 12308 14550
rect 12256 14486 12308 14492
rect 12164 13456 12216 13462
rect 12164 13398 12216 13404
rect 12176 13326 12204 13398
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12268 13190 12296 14486
rect 12532 14408 12584 14414
rect 12584 14368 12664 14396
rect 12532 14350 12584 14356
rect 12438 14104 12494 14113
rect 12438 14039 12440 14048
rect 12492 14039 12494 14048
rect 12440 14010 12492 14016
rect 12346 13832 12402 13841
rect 12346 13767 12348 13776
rect 12400 13767 12402 13776
rect 12440 13796 12492 13802
rect 12348 13738 12400 13744
rect 12440 13738 12492 13744
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 12256 13184 12308 13190
rect 12360 13161 12388 13194
rect 12256 13126 12308 13132
rect 12346 13152 12402 13161
rect 12346 13087 12402 13096
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 12072 12912 12124 12918
rect 12452 12866 12480 13738
rect 12532 13728 12584 13734
rect 12530 13696 12532 13705
rect 12584 13696 12586 13705
rect 12530 13631 12586 13640
rect 12636 13025 12664 14368
rect 12622 13016 12678 13025
rect 12622 12951 12678 12960
rect 12072 12854 12124 12860
rect 12084 12714 12112 12854
rect 12360 12838 12664 12866
rect 12360 12714 12388 12838
rect 12072 12708 12124 12714
rect 12072 12650 12124 12656
rect 12348 12708 12400 12714
rect 12348 12650 12400 12656
rect 11980 12164 12032 12170
rect 11980 12106 12032 12112
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 11992 11234 12020 12106
rect 12544 11914 12572 12106
rect 12360 11886 12572 11914
rect 12256 11824 12308 11830
rect 12256 11766 12308 11772
rect 11992 11206 12204 11234
rect 12268 11218 12296 11766
rect 12176 10198 12204 11206
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 12360 11121 12388 11886
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 12440 11620 12492 11626
rect 12440 11562 12492 11568
rect 12346 11112 12402 11121
rect 12346 11047 12402 11056
rect 12256 10736 12308 10742
rect 12256 10678 12308 10684
rect 12268 10606 12296 10678
rect 12256 10600 12308 10606
rect 12256 10542 12308 10548
rect 12164 10192 12216 10198
rect 12164 10134 12216 10140
rect 12256 9988 12308 9994
rect 12256 9930 12308 9936
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 12072 8560 12124 8566
rect 12072 8502 12124 8508
rect 12084 8430 12112 8502
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12084 7750 12112 8026
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11808 3534 11836 7278
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11992 6798 12020 7142
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11992 6254 12020 6734
rect 11888 6248 11940 6254
rect 11886 6216 11888 6225
rect 11980 6248 12032 6254
rect 11940 6216 11942 6225
rect 11980 6190 12032 6196
rect 11886 6151 11942 6160
rect 11992 5778 12020 6190
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11992 5234 12020 5714
rect 11980 5228 12032 5234
rect 11980 5170 12032 5176
rect 11992 4690 12020 5170
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 11978 3768 12034 3777
rect 11978 3703 12034 3712
rect 11992 3670 12020 3703
rect 11980 3664 12032 3670
rect 11980 3606 12032 3612
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11612 3120 11664 3126
rect 11900 3097 11928 3538
rect 11612 3062 11664 3068
rect 11886 3088 11942 3097
rect 11624 2938 11652 3062
rect 12084 3074 12112 3878
rect 12176 3194 12204 8842
rect 12268 8090 12296 9930
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12360 8838 12388 9454
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12452 6662 12480 11562
rect 12544 10606 12572 11766
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12544 8430 12572 10406
rect 12636 9518 12664 12838
rect 12728 12170 12756 15438
rect 12820 13802 12848 17206
rect 12912 16046 12940 25094
rect 13176 16992 13228 16998
rect 13176 16934 13228 16940
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 13188 16590 13216 16934
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 12992 16448 13044 16454
rect 12992 16390 13044 16396
rect 13004 16182 13032 16390
rect 12992 16176 13044 16182
rect 12992 16118 13044 16124
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12912 15502 12940 15982
rect 13544 15972 13596 15978
rect 13544 15914 13596 15920
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 13556 15094 13584 15914
rect 13636 15360 13688 15366
rect 13636 15302 13688 15308
rect 13084 15088 13136 15094
rect 13004 15048 13084 15076
rect 12808 13796 12860 13802
rect 12808 13738 12860 13744
rect 12806 12744 12862 12753
rect 12806 12679 12862 12688
rect 12716 12164 12768 12170
rect 12716 12106 12768 12112
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12636 9042 12664 9454
rect 12624 9036 12676 9042
rect 12624 8978 12676 8984
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 12268 6118 12296 6258
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 12256 5840 12308 5846
rect 12256 5782 12308 5788
rect 12346 5808 12402 5817
rect 12268 5545 12296 5782
rect 12346 5743 12402 5752
rect 12360 5710 12388 5743
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12254 5536 12310 5545
rect 12254 5471 12310 5480
rect 12348 4548 12400 4554
rect 12348 4490 12400 4496
rect 12254 4448 12310 4457
rect 12254 4383 12310 4392
rect 12268 3602 12296 4383
rect 12360 4185 12388 4490
rect 12544 4282 12572 8366
rect 12728 7834 12756 10950
rect 12820 10470 12848 12679
rect 12900 12300 12952 12306
rect 12900 12242 12952 12248
rect 12912 11830 12940 12242
rect 12900 11824 12952 11830
rect 12900 11766 12952 11772
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12808 9988 12860 9994
rect 12808 9930 12860 9936
rect 12820 9722 12848 9930
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 12912 9450 12940 11766
rect 13004 10198 13032 15048
rect 13084 15030 13136 15036
rect 13544 15088 13596 15094
rect 13544 15030 13596 15036
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 13096 14346 13124 14894
rect 13174 14376 13230 14385
rect 13084 14340 13136 14346
rect 13174 14311 13176 14320
rect 13084 14282 13136 14288
rect 13228 14311 13230 14320
rect 13176 14282 13228 14288
rect 13648 13870 13676 15302
rect 13832 14414 13860 16934
rect 14200 15094 14228 16934
rect 14292 15638 14320 28358
rect 14752 26234 14780 29038
rect 16316 26382 16344 36586
rect 16488 28076 16540 28082
rect 16488 28018 16540 28024
rect 16500 26518 16528 28018
rect 16488 26512 16540 26518
rect 16488 26454 16540 26460
rect 16304 26376 16356 26382
rect 16304 26318 16356 26324
rect 14752 26206 14872 26234
rect 14844 22642 14872 26206
rect 16316 25294 16344 26318
rect 16304 25288 16356 25294
rect 16304 25230 16356 25236
rect 14832 22636 14884 22642
rect 14832 22578 14884 22584
rect 14372 22432 14424 22438
rect 14372 22374 14424 22380
rect 14384 16658 14412 22374
rect 16120 19712 16172 19718
rect 16120 19654 16172 19660
rect 15476 19508 15528 19514
rect 15476 19450 15528 19456
rect 14924 17672 14976 17678
rect 14924 17614 14976 17620
rect 14936 17202 14964 17614
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 14924 17196 14976 17202
rect 14924 17138 14976 17144
rect 14936 17105 14964 17138
rect 14922 17096 14978 17105
rect 14922 17031 14978 17040
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 14384 16046 14412 16594
rect 14464 16516 14516 16522
rect 14464 16458 14516 16464
rect 15016 16516 15068 16522
rect 15016 16458 15068 16464
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14476 15706 14504 16458
rect 14556 16448 14608 16454
rect 14556 16390 14608 16396
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 14280 15632 14332 15638
rect 14280 15574 14332 15580
rect 14568 15434 14596 16390
rect 14556 15428 14608 15434
rect 14556 15370 14608 15376
rect 14922 15328 14978 15337
rect 14922 15263 14978 15272
rect 14188 15088 14240 15094
rect 14188 15030 14240 15036
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14648 14884 14700 14890
rect 14648 14826 14700 14832
rect 14002 14512 14058 14521
rect 14002 14447 14058 14456
rect 14462 14512 14518 14521
rect 14462 14447 14518 14456
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13372 13462 13400 13806
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13360 13456 13412 13462
rect 13360 13398 13412 13404
rect 13084 13252 13136 13258
rect 13084 13194 13136 13200
rect 13360 13252 13412 13258
rect 13360 13194 13412 13200
rect 13096 12782 13124 13194
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 13174 12744 13230 12753
rect 13174 12679 13230 12688
rect 13188 12374 13216 12679
rect 13176 12368 13228 12374
rect 13176 12310 13228 12316
rect 13188 11694 13216 12310
rect 13372 12306 13400 13194
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13464 12374 13492 12922
rect 13452 12368 13504 12374
rect 13452 12310 13504 12316
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 13084 10736 13136 10742
rect 13084 10678 13136 10684
rect 12992 10192 13044 10198
rect 12992 10134 13044 10140
rect 12900 9444 12952 9450
rect 12900 9386 12952 9392
rect 12636 7818 12756 7834
rect 12624 7812 12756 7818
rect 12676 7806 12756 7812
rect 12624 7754 12676 7760
rect 13096 7546 13124 10678
rect 13188 9926 13216 11018
rect 13266 10976 13322 10985
rect 13266 10911 13322 10920
rect 13280 10742 13308 10911
rect 13268 10736 13320 10742
rect 13268 10678 13320 10684
rect 13268 10600 13320 10606
rect 13266 10568 13268 10577
rect 13320 10568 13322 10577
rect 13266 10503 13322 10512
rect 13372 9994 13400 11494
rect 13464 11354 13492 12038
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13556 11218 13584 13466
rect 13648 11354 13676 13806
rect 13740 13530 13768 14282
rect 13818 14104 13874 14113
rect 13818 14039 13874 14048
rect 13832 13870 13860 14039
rect 13912 14000 13964 14006
rect 13910 13968 13912 13977
rect 13964 13968 13966 13977
rect 13910 13903 13966 13912
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13910 13832 13966 13841
rect 13910 13767 13912 13776
rect 13964 13767 13966 13776
rect 13912 13738 13964 13744
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13726 12608 13782 12617
rect 13726 12543 13782 12552
rect 13740 12306 13768 12543
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13740 11830 13768 12106
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13450 11112 13506 11121
rect 13450 11047 13452 11056
rect 13504 11047 13506 11056
rect 13452 11018 13504 11024
rect 13832 11014 13860 13126
rect 14016 12306 14044 14447
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14200 13161 14228 14214
rect 14186 13152 14242 13161
rect 14186 13087 14242 13096
rect 14094 13016 14150 13025
rect 14094 12951 14150 12960
rect 14004 12300 14056 12306
rect 14004 12242 14056 12248
rect 13912 11824 13964 11830
rect 13912 11766 13964 11772
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13634 10160 13690 10169
rect 13634 10095 13690 10104
rect 13360 9988 13412 9994
rect 13360 9930 13412 9936
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13280 8090 13308 9522
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12636 5545 12664 6394
rect 12912 6390 12940 6802
rect 12900 6384 12952 6390
rect 12900 6326 12952 6332
rect 12622 5536 12678 5545
rect 12622 5471 12678 5480
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12346 4176 12402 4185
rect 12346 4111 12402 4120
rect 12438 4040 12494 4049
rect 12438 3975 12494 3984
rect 12452 3738 12480 3975
rect 12622 3768 12678 3777
rect 12440 3732 12492 3738
rect 12622 3703 12624 3712
rect 12440 3674 12492 3680
rect 12676 3703 12678 3712
rect 12624 3674 12676 3680
rect 13280 3670 13308 7822
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13372 4457 13400 7346
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13358 4448 13414 4457
rect 13358 4383 13414 4392
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12348 3460 12400 3466
rect 12348 3402 12400 3408
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 12268 3074 12296 3130
rect 12084 3046 12296 3074
rect 12360 3058 12388 3402
rect 12348 3052 12400 3058
rect 11886 3023 11942 3032
rect 12348 2994 12400 3000
rect 11624 2910 11744 2938
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11336 2304 11388 2310
rect 11336 2246 11388 2252
rect 9692 1958 9904 1986
rect 9312 1692 9364 1698
rect 9312 1634 9364 1640
rect 9692 800 9720 1958
rect 11624 800 11652 2790
rect 11716 2650 11744 2910
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 12360 2582 12388 2994
rect 12728 2990 12756 3538
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12820 2825 12848 3130
rect 12900 3120 12952 3126
rect 12952 3080 13032 3108
rect 12900 3062 12952 3068
rect 13004 2990 13032 3080
rect 12992 2984 13044 2990
rect 12992 2926 13044 2932
rect 12806 2816 12862 2825
rect 12806 2751 12862 2760
rect 13280 2650 13308 3606
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 12348 2576 12400 2582
rect 12348 2518 12400 2524
rect 12348 2440 12400 2446
rect 12346 2408 12348 2417
rect 12400 2408 12402 2417
rect 12346 2343 12402 2352
rect 13372 1902 13400 3470
rect 13556 2378 13584 6598
rect 13648 5624 13676 10095
rect 13924 9382 13952 11766
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 14016 11150 14044 11630
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 14016 10742 14044 11086
rect 14004 10736 14056 10742
rect 14004 10678 14056 10684
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 14016 9722 14044 10542
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 13832 7274 13860 9046
rect 14016 8974 14044 9318
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 13912 8628 13964 8634
rect 14108 8616 14136 12951
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14200 12434 14228 12718
rect 14200 12406 14320 12434
rect 14188 8628 14240 8634
rect 14108 8588 14188 8616
rect 13912 8570 13964 8576
rect 14188 8570 14240 8576
rect 13924 8294 13952 8570
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 14108 7993 14136 8434
rect 14094 7984 14150 7993
rect 14094 7919 14150 7928
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 14108 7002 14136 7822
rect 14200 7206 14228 8570
rect 14292 7410 14320 12406
rect 14384 9110 14412 14350
rect 14476 13870 14504 14447
rect 14660 13870 14688 14826
rect 14740 14340 14792 14346
rect 14740 14282 14792 14288
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14752 13802 14780 14282
rect 14740 13796 14792 13802
rect 14740 13738 14792 13744
rect 14556 13728 14608 13734
rect 14648 13728 14700 13734
rect 14556 13670 14608 13676
rect 14646 13696 14648 13705
rect 14700 13696 14702 13705
rect 14464 13456 14516 13462
rect 14462 13424 14464 13433
rect 14516 13424 14518 13433
rect 14462 13359 14518 13368
rect 14476 13326 14504 13359
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14568 13258 14596 13670
rect 14646 13631 14702 13640
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14752 12782 14780 13738
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 14844 12434 14872 14894
rect 14936 14414 14964 15263
rect 15028 15162 15056 16458
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15120 15706 15148 15982
rect 15108 15700 15160 15706
rect 15108 15642 15160 15648
rect 15108 15428 15160 15434
rect 15108 15370 15160 15376
rect 15016 15156 15068 15162
rect 15016 15098 15068 15104
rect 14924 14408 14976 14414
rect 14924 14350 14976 14356
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 14936 12714 14964 13806
rect 15014 13424 15070 13433
rect 15014 13359 15070 13368
rect 15028 12782 15056 13359
rect 15016 12776 15068 12782
rect 15120 12753 15148 15370
rect 15016 12718 15068 12724
rect 15106 12744 15162 12753
rect 14924 12708 14976 12714
rect 14924 12650 14976 12656
rect 15028 12617 15056 12718
rect 15106 12679 15162 12688
rect 15014 12608 15070 12617
rect 15014 12543 15070 12552
rect 14752 12406 14872 12434
rect 14556 12368 14608 12374
rect 14556 12310 14608 12316
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14476 9518 14504 9998
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14372 9104 14424 9110
rect 14372 9046 14424 9052
rect 14372 8968 14424 8974
rect 14476 8922 14504 9454
rect 14424 8916 14504 8922
rect 14372 8910 14504 8916
rect 14384 8894 14504 8910
rect 14568 8906 14596 12310
rect 14752 10810 14780 12406
rect 14924 12300 14976 12306
rect 14924 12242 14976 12248
rect 14936 11830 14964 12242
rect 14924 11824 14976 11830
rect 14924 11766 14976 11772
rect 15016 11280 15068 11286
rect 15016 11222 15068 11228
rect 14924 11144 14976 11150
rect 14924 11086 14976 11092
rect 14740 10804 14792 10810
rect 14740 10746 14792 10752
rect 14648 10736 14700 10742
rect 14648 10678 14700 10684
rect 14660 9042 14688 10678
rect 14936 10606 14964 11086
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 14832 10532 14884 10538
rect 14832 10474 14884 10480
rect 14844 9722 14872 10474
rect 14936 10130 14964 10542
rect 15028 10538 15056 11222
rect 15016 10532 15068 10538
rect 15016 10474 15068 10480
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 15212 10033 15240 10066
rect 15198 10024 15254 10033
rect 14924 9988 14976 9994
rect 15198 9959 15254 9968
rect 14924 9930 14976 9936
rect 14936 9897 14964 9930
rect 14922 9888 14978 9897
rect 14922 9823 14978 9832
rect 14832 9716 14884 9722
rect 14832 9658 14884 9664
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 14648 9036 14700 9042
rect 14648 8978 14700 8984
rect 14476 8430 14504 8894
rect 14556 8900 14608 8906
rect 14556 8842 14608 8848
rect 14752 8566 14780 9590
rect 14740 8560 14792 8566
rect 14740 8502 14792 8508
rect 14464 8424 14516 8430
rect 14516 8384 14596 8412
rect 14464 8366 14516 8372
rect 14568 7886 14596 8384
rect 14556 7880 14608 7886
rect 14556 7822 14608 7828
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14464 7336 14516 7342
rect 14568 7290 14596 7822
rect 14516 7284 14596 7290
rect 14464 7278 14596 7284
rect 14476 7262 14596 7278
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13740 5914 13768 6258
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13728 5636 13780 5642
rect 13648 5596 13728 5624
rect 13648 4978 13676 5596
rect 13728 5578 13780 5584
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13740 5137 13768 5170
rect 13820 5160 13872 5166
rect 13726 5128 13782 5137
rect 13820 5102 13872 5108
rect 13726 5063 13782 5072
rect 13728 5024 13780 5030
rect 13648 4972 13728 4978
rect 13648 4966 13780 4972
rect 13648 4950 13768 4966
rect 13636 4616 13688 4622
rect 13634 4584 13636 4593
rect 13688 4584 13690 4593
rect 13634 4519 13690 4528
rect 13832 4214 13860 5102
rect 13820 4208 13872 4214
rect 13820 4150 13872 4156
rect 13912 3120 13964 3126
rect 13910 3088 13912 3097
rect 13964 3088 13966 3097
rect 13728 3052 13780 3058
rect 13910 3023 13966 3032
rect 13728 2994 13780 3000
rect 13636 2848 13688 2854
rect 13636 2790 13688 2796
rect 13544 2372 13596 2378
rect 13544 2314 13596 2320
rect 13360 1896 13412 1902
rect 13360 1838 13412 1844
rect 13648 1714 13676 2790
rect 13740 2553 13768 2994
rect 14108 2990 14136 6938
rect 14568 6866 14596 7262
rect 14556 6860 14608 6866
rect 14556 6802 14608 6808
rect 14568 6254 14596 6802
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14568 5778 14596 6190
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 14464 5296 14516 5302
rect 14464 5238 14516 5244
rect 14476 4842 14504 5238
rect 14568 5234 14596 5714
rect 14752 5370 14780 8502
rect 15304 8294 15332 16594
rect 15396 15094 15424 17478
rect 15384 15088 15436 15094
rect 15384 15030 15436 15036
rect 15488 14958 15516 19450
rect 16132 18290 16160 19654
rect 16212 18692 16264 18698
rect 16212 18634 16264 18640
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 15936 17808 15988 17814
rect 15936 17750 15988 17756
rect 15948 17134 15976 17750
rect 16028 17264 16080 17270
rect 16028 17206 16080 17212
rect 15844 17128 15896 17134
rect 15844 17070 15896 17076
rect 15936 17128 15988 17134
rect 15936 17070 15988 17076
rect 15660 17060 15712 17066
rect 15660 17002 15712 17008
rect 15568 15972 15620 15978
rect 15568 15914 15620 15920
rect 15580 15638 15608 15914
rect 15568 15632 15620 15638
rect 15568 15574 15620 15580
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15488 13190 15516 14894
rect 15672 13410 15700 17002
rect 15856 16726 15884 17070
rect 16040 17066 16068 17206
rect 16028 17060 16080 17066
rect 16028 17002 16080 17008
rect 15844 16720 15896 16726
rect 15844 16662 15896 16668
rect 15752 16448 15804 16454
rect 15752 16390 15804 16396
rect 15764 16182 15792 16390
rect 15752 16176 15804 16182
rect 15752 16118 15804 16124
rect 15752 15904 15804 15910
rect 15750 15872 15752 15881
rect 15804 15872 15806 15881
rect 15750 15807 15806 15816
rect 15672 13382 15792 13410
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15384 12912 15436 12918
rect 15384 12854 15436 12860
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 15396 7546 15424 12854
rect 15476 12776 15528 12782
rect 15764 12764 15792 13382
rect 15476 12718 15528 12724
rect 15580 12736 15792 12764
rect 15488 11626 15516 12718
rect 15580 12209 15608 12736
rect 15856 12434 15884 16662
rect 16028 15088 16080 15094
rect 16028 15030 16080 15036
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 15764 12406 15884 12434
rect 15566 12200 15622 12209
rect 15566 12135 15568 12144
rect 15620 12135 15622 12144
rect 15568 12106 15620 12112
rect 15580 12075 15608 12106
rect 15476 11620 15528 11626
rect 15476 11562 15528 11568
rect 15488 11218 15516 11562
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15580 11082 15608 11290
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15764 9382 15792 12406
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15764 8362 15792 9318
rect 15752 8356 15804 8362
rect 15752 8298 15804 8304
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15016 7472 15068 7478
rect 15016 7414 15068 7420
rect 14924 7200 14976 7206
rect 15028 7177 15056 7414
rect 14924 7142 14976 7148
rect 15014 7168 15070 7177
rect 14936 6338 14964 7142
rect 15014 7103 15070 7112
rect 15568 6996 15620 7002
rect 15568 6938 15620 6944
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 15580 6746 15608 6938
rect 15028 6474 15056 6734
rect 15580 6730 15792 6746
rect 15580 6724 15804 6730
rect 15580 6718 15752 6724
rect 15752 6666 15804 6672
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15106 6488 15162 6497
rect 15028 6446 15106 6474
rect 15106 6423 15162 6432
rect 15120 6390 15148 6423
rect 15108 6384 15160 6390
rect 14936 6310 15056 6338
rect 15108 6326 15160 6332
rect 14740 5364 14792 5370
rect 14740 5306 14792 5312
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 14832 5296 14884 5302
rect 14832 5238 14884 5244
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14556 5092 14608 5098
rect 14556 5034 14608 5040
rect 14568 5001 14596 5034
rect 14554 4992 14610 5001
rect 14554 4927 14610 4936
rect 14476 4814 14780 4842
rect 14648 4480 14700 4486
rect 14646 4448 14648 4457
rect 14700 4448 14702 4457
rect 14646 4383 14702 4392
rect 14554 4176 14610 4185
rect 14554 4111 14610 4120
rect 14568 4078 14596 4111
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 14646 4040 14702 4049
rect 14646 3975 14702 3984
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14568 3534 14596 3878
rect 14660 3670 14688 3975
rect 14752 3942 14780 4814
rect 14844 4554 14872 5238
rect 14936 4758 14964 5306
rect 14924 4752 14976 4758
rect 14924 4694 14976 4700
rect 14832 4548 14884 4554
rect 14832 4490 14884 4496
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14648 3664 14700 3670
rect 14648 3606 14700 3612
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14568 2990 14596 3470
rect 14844 3398 14872 4490
rect 14922 4312 14978 4321
rect 14922 4247 14978 4256
rect 14832 3392 14884 3398
rect 14832 3334 14884 3340
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 14556 2984 14608 2990
rect 14556 2926 14608 2932
rect 13726 2544 13782 2553
rect 14568 2514 14596 2926
rect 14936 2632 14964 4247
rect 15028 3602 15056 6310
rect 15304 6118 15332 6598
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15212 5778 15240 6054
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15948 3942 15976 12582
rect 16040 12481 16068 15030
rect 16026 12472 16082 12481
rect 16026 12407 16082 12416
rect 16132 11370 16160 18226
rect 16224 16658 16252 18634
rect 16776 17610 16804 37266
rect 18064 37262 18092 37402
rect 18144 37324 18196 37330
rect 18144 37266 18196 37272
rect 18052 37256 18104 37262
rect 18052 37198 18104 37204
rect 17592 27872 17644 27878
rect 17592 27814 17644 27820
rect 16948 25220 17000 25226
rect 16948 25162 17000 25168
rect 16960 18222 16988 25162
rect 17132 18896 17184 18902
rect 17132 18838 17184 18844
rect 17144 18630 17172 18838
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 17144 17678 17172 18566
rect 17408 18148 17460 18154
rect 17408 18090 17460 18096
rect 17132 17672 17184 17678
rect 17132 17614 17184 17620
rect 16764 17604 16816 17610
rect 16764 17546 16816 17552
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16580 17264 16632 17270
rect 16580 17206 16632 17212
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16212 16652 16264 16658
rect 16212 16594 16264 16600
rect 16408 16182 16436 16934
rect 16592 16590 16620 17206
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16396 16176 16448 16182
rect 16396 16118 16448 16124
rect 16304 15428 16356 15434
rect 16304 15370 16356 15376
rect 16316 15065 16344 15370
rect 16302 15056 16358 15065
rect 16302 14991 16358 15000
rect 16304 14884 16356 14890
rect 16304 14826 16356 14832
rect 16316 14414 16344 14826
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16396 14408 16448 14414
rect 16396 14350 16448 14356
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16224 13530 16252 13670
rect 16316 13530 16344 13874
rect 16408 13705 16436 14350
rect 16684 14006 16712 17478
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16776 16046 16804 17070
rect 16764 16040 16816 16046
rect 16948 16040 17000 16046
rect 16764 15982 16816 15988
rect 16868 16000 16948 16028
rect 16868 15366 16896 16000
rect 16948 15982 17000 15988
rect 16948 15632 17000 15638
rect 16948 15574 17000 15580
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 16672 14000 16724 14006
rect 16672 13942 16724 13948
rect 16394 13696 16450 13705
rect 16394 13631 16450 13640
rect 16212 13524 16264 13530
rect 16212 13466 16264 13472
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16408 12850 16436 13631
rect 16776 13258 16804 14418
rect 16868 13852 16896 15302
rect 16960 14482 16988 15574
rect 17144 15450 17172 17614
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 17236 15638 17264 16390
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17224 15632 17276 15638
rect 17224 15574 17276 15580
rect 17144 15422 17264 15450
rect 17040 14816 17092 14822
rect 17040 14758 17092 14764
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 17052 14006 17080 14758
rect 17236 14226 17264 15422
rect 17144 14198 17264 14226
rect 17040 14000 17092 14006
rect 17040 13942 17092 13948
rect 16948 13864 17000 13870
rect 16868 13824 16948 13852
rect 16948 13806 17000 13812
rect 16764 13252 16816 13258
rect 16764 13194 16816 13200
rect 16396 12844 16448 12850
rect 16316 12804 16396 12832
rect 16316 11762 16344 12804
rect 16396 12786 16448 12792
rect 16396 12368 16448 12374
rect 16396 12310 16448 12316
rect 17040 12368 17092 12374
rect 17040 12310 17092 12316
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16132 11342 16344 11370
rect 16212 11280 16264 11286
rect 16212 11222 16264 11228
rect 16028 8288 16080 8294
rect 16028 8230 16080 8236
rect 16040 7206 16068 8230
rect 16120 7472 16172 7478
rect 16120 7414 16172 7420
rect 16132 7274 16160 7414
rect 16120 7268 16172 7274
rect 16120 7210 16172 7216
rect 16028 7200 16080 7206
rect 16028 7142 16080 7148
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 16132 6225 16160 6258
rect 16118 6216 16174 6225
rect 16118 6151 16174 6160
rect 16132 5030 16160 6151
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16224 4554 16252 11222
rect 16316 5166 16344 11342
rect 16408 10198 16436 12310
rect 16672 12164 16724 12170
rect 16672 12106 16724 12112
rect 16578 11112 16634 11121
rect 16578 11047 16634 11056
rect 16592 10742 16620 11047
rect 16580 10736 16632 10742
rect 16580 10678 16632 10684
rect 16684 10266 16712 12106
rect 17052 11762 17080 12310
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16396 10192 16448 10198
rect 16396 10134 16448 10140
rect 17052 10130 17080 10610
rect 17040 10124 17092 10130
rect 16960 10084 17040 10112
rect 16486 10024 16542 10033
rect 16486 9959 16488 9968
rect 16540 9959 16542 9968
rect 16764 9988 16816 9994
rect 16488 9930 16540 9936
rect 16764 9930 16816 9936
rect 16488 9648 16540 9654
rect 16488 9590 16540 9596
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 16408 9081 16436 9386
rect 16500 9110 16528 9590
rect 16776 9518 16804 9930
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16868 9194 16896 9454
rect 16684 9166 16896 9194
rect 16488 9104 16540 9110
rect 16394 9072 16450 9081
rect 16488 9046 16540 9052
rect 16394 9007 16396 9016
rect 16448 9007 16450 9016
rect 16396 8978 16448 8984
rect 16486 6624 16542 6633
rect 16486 6559 16542 6568
rect 16500 6254 16528 6559
rect 16488 6248 16540 6254
rect 16488 6190 16540 6196
rect 16684 6186 16712 9166
rect 16960 9058 16988 10084
rect 17040 10066 17092 10072
rect 17144 9194 17172 14198
rect 17224 12912 17276 12918
rect 17224 12854 17276 12860
rect 16868 9042 16988 9058
rect 16856 9036 16988 9042
rect 16908 9030 16988 9036
rect 17052 9166 17172 9194
rect 16856 8978 16908 8984
rect 17052 8242 17080 9166
rect 17132 9036 17184 9042
rect 17132 8978 17184 8984
rect 16960 8214 17080 8242
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16672 6180 16724 6186
rect 16672 6122 16724 6128
rect 16670 6080 16726 6089
rect 16670 6015 16726 6024
rect 16684 5846 16712 6015
rect 16672 5840 16724 5846
rect 16672 5782 16724 5788
rect 16488 5296 16540 5302
rect 16486 5264 16488 5273
rect 16540 5264 16542 5273
rect 16486 5199 16542 5208
rect 16304 5160 16356 5166
rect 16304 5102 16356 5108
rect 16212 4548 16264 4554
rect 16132 4508 16212 4536
rect 15660 3936 15712 3942
rect 15212 3896 15660 3924
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 15212 3466 15240 3896
rect 15660 3878 15712 3884
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 15200 3460 15252 3466
rect 15200 3402 15252 3408
rect 16132 2854 16160 4508
rect 16212 4490 16264 4496
rect 16316 4214 16344 5102
rect 16684 4554 16712 5782
rect 16868 4758 16896 7278
rect 16856 4752 16908 4758
rect 16856 4694 16908 4700
rect 16672 4548 16724 4554
rect 16672 4490 16724 4496
rect 16854 4312 16910 4321
rect 16854 4247 16910 4256
rect 16212 4208 16264 4214
rect 16212 4150 16264 4156
rect 16304 4208 16356 4214
rect 16304 4150 16356 4156
rect 16488 4208 16540 4214
rect 16488 4150 16540 4156
rect 16224 4060 16252 4150
rect 16500 4060 16528 4150
rect 16868 4146 16896 4247
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 16224 4032 16528 4060
rect 16960 3942 16988 8214
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 17052 5166 17080 8026
rect 17144 7750 17172 8978
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 17132 6928 17184 6934
rect 17132 6870 17184 6876
rect 17144 6118 17172 6870
rect 17236 6798 17264 12854
rect 17328 12170 17356 16186
rect 17420 15366 17448 18090
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 17512 15434 17540 17478
rect 17604 16726 17632 27814
rect 17776 24132 17828 24138
rect 17776 24074 17828 24080
rect 17788 22094 17816 24074
rect 17696 22066 17816 22094
rect 17592 16720 17644 16726
rect 17592 16662 17644 16668
rect 17696 16538 17724 22066
rect 17776 21548 17828 21554
rect 17776 21490 17828 21496
rect 17604 16510 17724 16538
rect 17500 15428 17552 15434
rect 17500 15370 17552 15376
rect 17408 15360 17460 15366
rect 17408 15302 17460 15308
rect 17420 14482 17448 15302
rect 17604 14958 17632 16510
rect 17684 16448 17736 16454
rect 17684 16390 17736 16396
rect 17592 14952 17644 14958
rect 17590 14920 17592 14929
rect 17644 14920 17646 14929
rect 17590 14855 17646 14864
rect 17500 14544 17552 14550
rect 17500 14486 17552 14492
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17512 14346 17540 14486
rect 17500 14340 17552 14346
rect 17500 14282 17552 14288
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 17316 12164 17368 12170
rect 17316 12106 17368 12112
rect 17328 11898 17356 12106
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17314 11248 17370 11257
rect 17314 11183 17370 11192
rect 17328 10130 17356 11183
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17328 9994 17356 10066
rect 17316 9988 17368 9994
rect 17316 9930 17368 9936
rect 17420 9761 17448 12786
rect 17590 12336 17646 12345
rect 17590 12271 17646 12280
rect 17604 11694 17632 12271
rect 17592 11688 17644 11694
rect 17592 11630 17644 11636
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17406 9752 17462 9761
rect 17406 9687 17462 9696
rect 17512 8922 17540 10202
rect 17420 8906 17632 8922
rect 17408 8900 17632 8906
rect 17460 8894 17632 8900
rect 17408 8842 17460 8848
rect 17314 8528 17370 8537
rect 17314 8463 17316 8472
rect 17368 8463 17370 8472
rect 17316 8434 17368 8440
rect 17500 8356 17552 8362
rect 17500 8298 17552 8304
rect 17316 7812 17368 7818
rect 17316 7754 17368 7760
rect 17328 7478 17356 7754
rect 17316 7472 17368 7478
rect 17316 7414 17368 7420
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17236 6118 17264 6598
rect 17132 6112 17184 6118
rect 17132 6054 17184 6060
rect 17224 6112 17276 6118
rect 17224 6054 17276 6060
rect 17132 5228 17184 5234
rect 17132 5170 17184 5176
rect 17040 5160 17092 5166
rect 17040 5102 17092 5108
rect 17144 4690 17172 5170
rect 17132 4684 17184 4690
rect 17132 4626 17184 4632
rect 17052 4134 17264 4162
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 17052 3754 17080 4134
rect 17236 4078 17264 4134
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 16960 3726 17080 3754
rect 17144 3738 17172 4014
rect 17328 3913 17356 7414
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17420 5642 17448 7346
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 17314 3904 17370 3913
rect 17314 3839 17370 3848
rect 17132 3732 17184 3738
rect 16212 3460 16264 3466
rect 16212 3402 16264 3408
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 14844 2604 14964 2632
rect 13726 2479 13782 2488
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 13556 1686 13676 1714
rect 13556 800 13584 1686
rect 14844 800 14872 2604
rect 16224 1970 16252 3402
rect 16960 2990 16988 3726
rect 17132 3674 17184 3680
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 17132 3596 17184 3602
rect 17132 3538 17184 3544
rect 17144 3194 17172 3538
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 16948 2984 17000 2990
rect 16948 2926 17000 2932
rect 17144 2514 17172 3130
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 16212 1964 16264 1970
rect 16212 1906 16264 1912
rect 16776 870 16896 898
rect 16776 800 16804 870
rect 18 200 74 800
rect 1306 200 1362 800
rect 3238 200 3294 800
rect 4526 200 4582 800
rect 6458 200 6514 800
rect 8390 200 8446 800
rect 9678 200 9734 800
rect 11610 200 11666 800
rect 13542 200 13598 800
rect 14830 200 14886 800
rect 16762 200 16818 800
rect 16868 762 16896 870
rect 17236 762 17264 3674
rect 17314 3496 17370 3505
rect 17314 3431 17370 3440
rect 17328 3398 17356 3431
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 17420 3210 17448 5578
rect 17512 3398 17540 8298
rect 17604 6934 17632 8894
rect 17696 7546 17724 16390
rect 17788 12850 17816 21490
rect 17868 17060 17920 17066
rect 17868 17002 17920 17008
rect 17880 16658 17908 17002
rect 18052 16720 18104 16726
rect 18052 16662 18104 16668
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 18064 16522 18092 16662
rect 18052 16516 18104 16522
rect 18052 16458 18104 16464
rect 17960 15972 18012 15978
rect 17960 15914 18012 15920
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 17880 15026 17908 15642
rect 17972 15434 18000 15914
rect 18156 15910 18184 37266
rect 19996 37126 20024 39200
rect 21928 37330 21956 39200
rect 21916 37324 21968 37330
rect 21916 37266 21968 37272
rect 20076 37256 20128 37262
rect 20076 37198 20128 37204
rect 20536 37256 20588 37262
rect 20536 37198 20588 37204
rect 23020 37256 23072 37262
rect 23020 37198 23072 37204
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19984 35080 20036 35086
rect 19984 35022 20036 35028
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19996 32434 20024 35022
rect 19984 32428 20036 32434
rect 19984 32370 20036 32376
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 20088 26234 20116 37198
rect 20548 29170 20576 37198
rect 20720 37188 20772 37194
rect 20720 37130 20772 37136
rect 20732 35290 20760 37130
rect 22100 36916 22152 36922
rect 22100 36858 22152 36864
rect 20720 35284 20772 35290
rect 20720 35226 20772 35232
rect 20536 29164 20588 29170
rect 20536 29106 20588 29112
rect 20260 29028 20312 29034
rect 20260 28970 20312 28976
rect 19996 26206 20116 26234
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 18236 25900 18288 25906
rect 18236 25842 18288 25848
rect 18248 18970 18276 25842
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19996 21690 20024 26206
rect 19984 21684 20036 21690
rect 19984 21626 20036 21632
rect 19432 20800 19484 20806
rect 19432 20742 19484 20748
rect 19444 20534 19472 20742
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 19432 20528 19484 20534
rect 19432 20470 19484 20476
rect 19156 20392 19208 20398
rect 19156 20334 19208 20340
rect 18236 18964 18288 18970
rect 18236 18906 18288 18912
rect 18512 18964 18564 18970
rect 18512 18906 18564 18912
rect 18236 18760 18288 18766
rect 18236 18702 18288 18708
rect 18248 18086 18276 18702
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 18248 17678 18276 18022
rect 18420 17740 18472 17746
rect 18420 17682 18472 17688
rect 18236 17672 18288 17678
rect 18236 17614 18288 17620
rect 18328 17264 18380 17270
rect 18328 17206 18380 17212
rect 18340 16250 18368 17206
rect 18432 17202 18460 17682
rect 18420 17196 18472 17202
rect 18420 17138 18472 17144
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 18144 15904 18196 15910
rect 18144 15846 18196 15852
rect 18524 15502 18552 18906
rect 18788 18624 18840 18630
rect 18788 18566 18840 18572
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18512 15496 18564 15502
rect 18512 15438 18564 15444
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 18144 15360 18196 15366
rect 18142 15328 18144 15337
rect 18196 15328 18198 15337
rect 18142 15263 18198 15272
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 17868 15020 17920 15026
rect 17868 14962 17920 14968
rect 17972 14414 18000 15098
rect 18156 15094 18184 15263
rect 18616 15094 18644 17478
rect 18708 15586 18736 17614
rect 18800 17270 18828 18566
rect 19168 18086 19196 20334
rect 19352 20058 19380 20470
rect 19616 20256 19668 20262
rect 19616 20198 19668 20204
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19628 19854 19656 20198
rect 19616 19848 19668 19854
rect 19616 19790 19668 19796
rect 19984 19780 20036 19786
rect 19984 19722 20036 19728
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19892 19236 19944 19242
rect 19892 19178 19944 19184
rect 19904 18873 19932 19178
rect 19890 18864 19946 18873
rect 19432 18828 19484 18834
rect 19890 18799 19946 18808
rect 19432 18770 19484 18776
rect 19340 18148 19392 18154
rect 19340 18090 19392 18096
rect 19156 18080 19208 18086
rect 19156 18022 19208 18028
rect 18788 17264 18840 17270
rect 18788 17206 18840 17212
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18800 15706 18828 15982
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 18708 15558 18828 15586
rect 18144 15088 18196 15094
rect 18144 15030 18196 15036
rect 18604 15088 18656 15094
rect 18604 15030 18656 15036
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 17866 13968 17922 13977
rect 17866 13903 17922 13912
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17880 11778 17908 13903
rect 17788 11750 17908 11778
rect 17788 9518 17816 11750
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17880 11121 17908 11630
rect 17866 11112 17922 11121
rect 17866 11047 17922 11056
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17776 8084 17828 8090
rect 17776 8026 17828 8032
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17788 7426 17816 8026
rect 17696 7410 17816 7426
rect 17880 7410 17908 10066
rect 17972 9722 18000 14350
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18144 13796 18196 13802
rect 18144 13738 18196 13744
rect 18236 13796 18288 13802
rect 18236 13738 18288 13744
rect 18156 11082 18184 13738
rect 18248 13530 18276 13738
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18236 13252 18288 13258
rect 18236 13194 18288 13200
rect 18248 12986 18276 13194
rect 18236 12980 18288 12986
rect 18236 12922 18288 12928
rect 18248 12782 18276 12922
rect 18328 12912 18380 12918
rect 18326 12880 18328 12889
rect 18380 12880 18382 12889
rect 18326 12815 18382 12824
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 18144 11076 18196 11082
rect 18144 11018 18196 11024
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 18064 7857 18092 10950
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 18156 9110 18184 9590
rect 18144 9104 18196 9110
rect 18144 9046 18196 9052
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 18156 8634 18184 8774
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 18050 7848 18106 7857
rect 18050 7783 18106 7792
rect 18248 7546 18276 11766
rect 18432 10198 18460 14010
rect 18708 13938 18736 14486
rect 18696 13932 18748 13938
rect 18696 13874 18748 13880
rect 18604 13524 18656 13530
rect 18604 13466 18656 13472
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18524 12782 18552 13330
rect 18512 12776 18564 12782
rect 18512 12718 18564 12724
rect 18524 12646 18552 12718
rect 18512 12640 18564 12646
rect 18512 12582 18564 12588
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18524 10810 18552 11086
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18420 10192 18472 10198
rect 18326 10160 18382 10169
rect 18420 10134 18472 10140
rect 18326 10095 18382 10104
rect 18340 9994 18368 10095
rect 18328 9988 18380 9994
rect 18328 9930 18380 9936
rect 18512 8560 18564 8566
rect 18512 8502 18564 8508
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18524 7449 18552 8502
rect 18510 7440 18566 7449
rect 17684 7404 17816 7410
rect 17736 7398 17816 7404
rect 17868 7404 17920 7410
rect 17684 7346 17736 7352
rect 18510 7375 18566 7384
rect 17868 7346 17920 7352
rect 17776 7336 17828 7342
rect 17776 7278 17828 7284
rect 17682 7032 17738 7041
rect 17682 6967 17738 6976
rect 17696 6934 17724 6967
rect 17592 6928 17644 6934
rect 17592 6870 17644 6876
rect 17684 6928 17736 6934
rect 17684 6870 17736 6876
rect 17788 6866 17816 7278
rect 17958 6896 18014 6905
rect 17776 6860 17828 6866
rect 17958 6831 17960 6840
rect 17776 6802 17828 6808
rect 18012 6831 18014 6840
rect 17960 6802 18012 6808
rect 17592 6656 17644 6662
rect 17590 6624 17592 6633
rect 17644 6624 17646 6633
rect 17646 6582 17724 6610
rect 17590 6559 17646 6568
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17420 3182 17632 3210
rect 17604 2990 17632 3182
rect 17592 2984 17644 2990
rect 17592 2926 17644 2932
rect 17696 2378 17724 6582
rect 17788 6322 17816 6802
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 17776 6316 17828 6322
rect 17776 6258 17828 6264
rect 17788 5778 17816 6258
rect 18156 5778 18184 6394
rect 18616 6254 18644 13466
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18708 12646 18736 12922
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18696 11688 18748 11694
rect 18696 11630 18748 11636
rect 18708 11082 18736 11630
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18800 9926 18828 15558
rect 18880 15088 18932 15094
rect 18880 15030 18932 15036
rect 18892 12374 18920 15030
rect 18970 14920 19026 14929
rect 18970 14855 19026 14864
rect 18984 14346 19012 14855
rect 18972 14340 19024 14346
rect 18972 14282 19024 14288
rect 19076 14006 19104 16050
rect 19168 15978 19196 18022
rect 19352 17066 19380 18090
rect 19444 17320 19472 18770
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 18222 20024 19722
rect 20076 19712 20128 19718
rect 20076 19654 20128 19660
rect 20088 18358 20116 19654
rect 20168 19168 20220 19174
rect 20168 19110 20220 19116
rect 20180 18698 20208 19110
rect 20168 18692 20220 18698
rect 20168 18634 20220 18640
rect 20076 18352 20128 18358
rect 20076 18294 20128 18300
rect 19984 18216 20036 18222
rect 19984 18158 20036 18164
rect 19890 17776 19946 17785
rect 19890 17711 19892 17720
rect 19944 17711 19946 17720
rect 19892 17682 19944 17688
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19892 17332 19944 17338
rect 19444 17292 19564 17320
rect 19340 17060 19392 17066
rect 19340 17002 19392 17008
rect 19156 15972 19208 15978
rect 19156 15914 19208 15920
rect 19352 15094 19380 17002
rect 19536 16436 19564 17292
rect 19892 17274 19944 17280
rect 19708 17264 19760 17270
rect 19708 17206 19760 17212
rect 19616 17128 19668 17134
rect 19616 17070 19668 17076
rect 19628 16522 19656 17070
rect 19720 16726 19748 17206
rect 19904 17134 19932 17274
rect 19892 17128 19944 17134
rect 19892 17070 19944 17076
rect 19708 16720 19760 16726
rect 19708 16662 19760 16668
rect 19616 16516 19668 16522
rect 19616 16458 19668 16464
rect 19444 16408 19564 16436
rect 19340 15088 19392 15094
rect 19340 15030 19392 15036
rect 19444 15026 19472 16408
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19890 15736 19946 15745
rect 19890 15671 19946 15680
rect 19524 15632 19576 15638
rect 19522 15600 19524 15609
rect 19576 15600 19578 15609
rect 19522 15535 19578 15544
rect 19904 15502 19932 15671
rect 19996 15638 20024 18158
rect 20272 17746 20300 28970
rect 22112 27062 22140 36858
rect 23032 36786 23060 37198
rect 23216 37126 23244 39200
rect 23296 37256 23348 37262
rect 23296 37198 23348 37204
rect 23204 37120 23256 37126
rect 23204 37062 23256 37068
rect 23308 36922 23336 37198
rect 25148 37126 25176 39200
rect 25872 37256 25924 37262
rect 25872 37198 25924 37204
rect 25136 37120 25188 37126
rect 25136 37062 25188 37068
rect 23296 36916 23348 36922
rect 23296 36858 23348 36864
rect 22284 36780 22336 36786
rect 22284 36722 22336 36728
rect 22744 36780 22796 36786
rect 22744 36722 22796 36728
rect 23020 36780 23072 36786
rect 23020 36722 23072 36728
rect 22296 28762 22324 36722
rect 22756 36582 22784 36722
rect 22744 36576 22796 36582
rect 22744 36518 22796 36524
rect 22756 36378 22784 36518
rect 22744 36372 22796 36378
rect 22744 36314 22796 36320
rect 22284 28756 22336 28762
rect 22284 28698 22336 28704
rect 22296 28558 22324 28698
rect 22284 28552 22336 28558
rect 22284 28494 22336 28500
rect 22652 28416 22704 28422
rect 22652 28358 22704 28364
rect 22100 27056 22152 27062
rect 22100 26998 22152 27004
rect 22100 19848 22152 19854
rect 22100 19790 22152 19796
rect 20352 19372 20404 19378
rect 20352 19314 20404 19320
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 20076 17672 20128 17678
rect 20128 17620 20208 17626
rect 20076 17614 20208 17620
rect 20088 17598 20208 17614
rect 20180 16794 20208 17598
rect 20364 17338 20392 19314
rect 21088 19236 21140 19242
rect 21088 19178 21140 19184
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 20352 17332 20404 17338
rect 20352 17274 20404 17280
rect 20168 16788 20220 16794
rect 20168 16730 20220 16736
rect 20076 16516 20128 16522
rect 20076 16458 20128 16464
rect 20088 15910 20116 16458
rect 20076 15904 20128 15910
rect 20076 15846 20128 15852
rect 19984 15632 20036 15638
rect 19984 15574 20036 15580
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 20074 15464 20130 15473
rect 20074 15399 20076 15408
rect 20128 15399 20130 15408
rect 20076 15370 20128 15376
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19892 15088 19944 15094
rect 20076 15088 20128 15094
rect 19944 15048 20076 15076
rect 19892 15030 19944 15036
rect 20076 15030 20128 15036
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19248 14952 19300 14958
rect 19248 14894 19300 14900
rect 19064 14000 19116 14006
rect 19064 13942 19116 13948
rect 19076 13394 19104 13942
rect 19156 13864 19208 13870
rect 19154 13832 19156 13841
rect 19208 13832 19210 13841
rect 19154 13767 19210 13776
rect 19260 13433 19288 14894
rect 19432 14816 19484 14822
rect 19812 14793 19840 14962
rect 19432 14758 19484 14764
rect 19798 14784 19854 14793
rect 19444 14482 19472 14758
rect 19798 14719 19854 14728
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19246 13424 19302 13433
rect 19064 13388 19116 13394
rect 19246 13359 19302 13368
rect 19064 13330 19116 13336
rect 19246 13288 19302 13297
rect 19246 13223 19302 13232
rect 19260 12764 19288 13223
rect 19352 12866 19380 14350
rect 19444 14056 19472 14418
rect 20180 14362 20208 16730
rect 20456 16658 20484 18770
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 20536 18148 20588 18154
rect 20536 18090 20588 18096
rect 20444 16652 20496 16658
rect 20444 16594 20496 16600
rect 20260 16516 20312 16522
rect 20260 16458 20312 16464
rect 20272 15570 20300 16458
rect 20352 16176 20404 16182
rect 20352 16118 20404 16124
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 19996 14334 20208 14362
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19444 14028 19564 14056
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19444 12986 19472 13806
rect 19536 13394 19564 14028
rect 19614 13560 19670 13569
rect 19614 13495 19670 13504
rect 19524 13388 19576 13394
rect 19524 13330 19576 13336
rect 19628 13258 19656 13495
rect 19996 13444 20024 14334
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 19996 13416 20116 13444
rect 19892 13388 19944 13394
rect 19944 13348 20024 13376
rect 19892 13330 19944 13336
rect 19616 13252 19668 13258
rect 19616 13194 19668 13200
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19352 12838 19472 12866
rect 19340 12776 19392 12782
rect 19260 12736 19340 12764
rect 19340 12718 19392 12724
rect 18880 12368 18932 12374
rect 18880 12310 18932 12316
rect 18972 12300 19024 12306
rect 18972 12242 19024 12248
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 18984 11694 19012 12242
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 19076 11830 19104 12038
rect 19064 11824 19116 11830
rect 19064 11766 19116 11772
rect 18972 11688 19024 11694
rect 18972 11630 19024 11636
rect 18880 10600 18932 10606
rect 18880 10542 18932 10548
rect 18788 9920 18840 9926
rect 18788 9862 18840 9868
rect 18786 8936 18842 8945
rect 18786 8871 18788 8880
rect 18840 8871 18842 8880
rect 18788 8842 18840 8848
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18708 7546 18736 7686
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18800 7206 18828 7822
rect 18788 7200 18840 7206
rect 18788 7142 18840 7148
rect 18788 6928 18840 6934
rect 18788 6870 18840 6876
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18420 5840 18472 5846
rect 18420 5782 18472 5788
rect 17776 5772 17828 5778
rect 17776 5714 17828 5720
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 17788 5302 17816 5714
rect 18432 5658 18460 5782
rect 17880 5630 18460 5658
rect 17776 5296 17828 5302
rect 17776 5238 17828 5244
rect 17880 4078 17908 5630
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 18064 5001 18092 5102
rect 18050 4992 18106 5001
rect 18050 4927 18106 4936
rect 18800 4826 18828 6870
rect 18892 6798 18920 10542
rect 18984 9110 19012 11630
rect 19156 11620 19208 11626
rect 19156 11562 19208 11568
rect 19168 11286 19196 11562
rect 19156 11280 19208 11286
rect 19156 11222 19208 11228
rect 19260 11218 19288 12242
rect 19444 12238 19472 12838
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19432 12232 19484 12238
rect 19430 12200 19432 12209
rect 19484 12200 19486 12209
rect 19340 12164 19392 12170
rect 19430 12135 19486 12144
rect 19340 12106 19392 12112
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 19064 11008 19116 11014
rect 19064 10950 19116 10956
rect 19076 10606 19104 10950
rect 19156 10804 19208 10810
rect 19156 10746 19208 10752
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 19076 9722 19104 10542
rect 19168 10266 19196 10746
rect 19352 10305 19380 12106
rect 19536 12084 19564 12718
rect 19708 12436 19760 12442
rect 19708 12378 19760 12384
rect 19720 12170 19748 12378
rect 19708 12164 19760 12170
rect 19708 12106 19760 12112
rect 19444 12056 19564 12084
rect 19444 11880 19472 12056
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19444 11852 19564 11880
rect 19432 11280 19484 11286
rect 19430 11248 19432 11257
rect 19484 11248 19486 11257
rect 19430 11183 19486 11192
rect 19536 11014 19564 11852
rect 19996 11694 20024 13348
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 20088 11506 20116 13416
rect 20180 11830 20208 14214
rect 20272 14006 20300 15302
rect 20364 15162 20392 16118
rect 20456 15978 20484 16594
rect 20444 15972 20496 15978
rect 20444 15914 20496 15920
rect 20548 15706 20576 18090
rect 20626 17776 20682 17785
rect 20626 17711 20628 17720
rect 20680 17711 20682 17720
rect 20628 17682 20680 17688
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20732 16522 20760 17478
rect 21008 17338 21036 18362
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 21100 17202 21128 19178
rect 22112 18766 22140 19790
rect 22100 18760 22152 18766
rect 22100 18702 22152 18708
rect 22664 18358 22692 28358
rect 23388 26784 23440 26790
rect 23388 26726 23440 26732
rect 23400 26586 23428 26726
rect 23388 26580 23440 26586
rect 23388 26522 23440 26528
rect 23400 20058 23428 26522
rect 25228 25152 25280 25158
rect 25228 25094 25280 25100
rect 24124 24132 24176 24138
rect 24124 24074 24176 24080
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 23400 19854 23428 19994
rect 23388 19848 23440 19854
rect 23388 19790 23440 19796
rect 23112 19712 23164 19718
rect 23112 19654 23164 19660
rect 23020 19168 23072 19174
rect 23020 19110 23072 19116
rect 22560 18352 22612 18358
rect 22560 18294 22612 18300
rect 22652 18352 22704 18358
rect 22652 18294 22704 18300
rect 21180 18080 21232 18086
rect 21180 18022 21232 18028
rect 22284 18080 22336 18086
rect 22284 18022 22336 18028
rect 21192 17270 21220 18022
rect 22296 17678 22324 18022
rect 22572 17882 22600 18294
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 22664 17746 22692 18294
rect 22376 17740 22428 17746
rect 22376 17682 22428 17688
rect 22652 17740 22704 17746
rect 22652 17682 22704 17688
rect 21640 17672 21692 17678
rect 21640 17614 21692 17620
rect 22284 17672 22336 17678
rect 22284 17614 22336 17620
rect 21180 17264 21232 17270
rect 21180 17206 21232 17212
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 21456 17060 21508 17066
rect 21456 17002 21508 17008
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 20904 16720 20956 16726
rect 20904 16662 20956 16668
rect 20720 16516 20772 16522
rect 20720 16458 20772 16464
rect 20628 16448 20680 16454
rect 20628 16390 20680 16396
rect 20812 16448 20864 16454
rect 20812 16390 20864 16396
rect 20640 15978 20668 16390
rect 20628 15972 20680 15978
rect 20628 15914 20680 15920
rect 20536 15700 20588 15706
rect 20536 15642 20588 15648
rect 20444 15632 20496 15638
rect 20444 15574 20496 15580
rect 20534 15600 20590 15609
rect 20456 15434 20484 15574
rect 20534 15535 20590 15544
rect 20548 15502 20576 15535
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 20444 15428 20496 15434
rect 20444 15370 20496 15376
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20456 15042 20484 15370
rect 20718 15328 20774 15337
rect 20718 15263 20774 15272
rect 20364 15014 20484 15042
rect 20536 15020 20588 15026
rect 20364 14482 20392 15014
rect 20536 14962 20588 14968
rect 20548 14929 20576 14962
rect 20534 14920 20590 14929
rect 20732 14890 20760 15263
rect 20534 14855 20590 14864
rect 20720 14884 20772 14890
rect 20720 14826 20772 14832
rect 20720 14544 20772 14550
rect 20720 14486 20772 14492
rect 20352 14476 20404 14482
rect 20352 14418 20404 14424
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 20260 14000 20312 14006
rect 20260 13942 20312 13948
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20272 12306 20300 13262
rect 20352 13252 20404 13258
rect 20352 13194 20404 13200
rect 20364 12442 20392 13194
rect 20456 12918 20484 14010
rect 20628 13728 20680 13734
rect 20628 13670 20680 13676
rect 20640 13433 20668 13670
rect 20626 13424 20682 13433
rect 20626 13359 20682 13368
rect 20536 13184 20588 13190
rect 20536 13126 20588 13132
rect 20444 12912 20496 12918
rect 20444 12854 20496 12860
rect 20456 12442 20484 12854
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 20444 12436 20496 12442
rect 20444 12378 20496 12384
rect 20364 12306 20392 12378
rect 20260 12300 20312 12306
rect 20260 12242 20312 12248
rect 20352 12300 20404 12306
rect 20352 12242 20404 12248
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 20088 11478 20392 11506
rect 20258 11384 20314 11393
rect 19892 11348 19944 11354
rect 20258 11319 20314 11328
rect 19892 11290 19944 11296
rect 19904 11218 19932 11290
rect 19892 11212 19944 11218
rect 19892 11154 19944 11160
rect 19524 11008 19576 11014
rect 19524 10950 19576 10956
rect 20076 11008 20128 11014
rect 20076 10950 20128 10956
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19522 10704 19578 10713
rect 19522 10639 19524 10648
rect 19576 10639 19578 10648
rect 19524 10610 19576 10616
rect 19338 10296 19394 10305
rect 19156 10260 19208 10266
rect 19338 10231 19394 10240
rect 19706 10296 19762 10305
rect 19706 10231 19762 10240
rect 19156 10202 19208 10208
rect 19248 10192 19300 10198
rect 19616 10192 19668 10198
rect 19300 10140 19616 10146
rect 19248 10134 19668 10140
rect 19260 10118 19656 10134
rect 19616 9988 19668 9994
rect 19260 9948 19616 9976
rect 19156 9920 19208 9926
rect 19260 9897 19288 9948
rect 19616 9930 19668 9936
rect 19720 9926 19748 10231
rect 19708 9920 19760 9926
rect 19156 9862 19208 9868
rect 19246 9888 19302 9897
rect 19064 9716 19116 9722
rect 19064 9658 19116 9664
rect 19168 9602 19196 9862
rect 19708 9862 19760 9868
rect 19246 9823 19302 9832
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19430 9752 19486 9761
rect 19574 9755 19882 9764
rect 19430 9687 19486 9696
rect 19076 9574 19196 9602
rect 18972 9104 19024 9110
rect 18972 9046 19024 9052
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 18892 4162 18920 6734
rect 19076 5098 19104 9574
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 19352 8412 19380 9454
rect 19444 8537 19472 9687
rect 20088 9674 20116 10950
rect 20168 10736 20220 10742
rect 20168 10678 20220 10684
rect 20180 9761 20208 10678
rect 20166 9752 20222 9761
rect 20166 9687 20222 9696
rect 19996 9646 20116 9674
rect 19614 9072 19670 9081
rect 19614 9007 19670 9016
rect 19628 8974 19656 9007
rect 19616 8968 19668 8974
rect 19616 8910 19668 8916
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19430 8528 19486 8537
rect 19996 8498 20024 9646
rect 20180 9586 20208 9687
rect 20168 9580 20220 9586
rect 20168 9522 20220 9528
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 19430 8463 19486 8472
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19352 8384 19472 8412
rect 19248 8356 19300 8362
rect 19248 8298 19300 8304
rect 19260 8022 19288 8298
rect 19340 8288 19392 8294
rect 19340 8230 19392 8236
rect 19248 8016 19300 8022
rect 19248 7958 19300 7964
rect 19352 7954 19380 8230
rect 19340 7948 19392 7954
rect 19340 7890 19392 7896
rect 19352 7478 19380 7890
rect 19340 7472 19392 7478
rect 19340 7414 19392 7420
rect 19444 6905 19472 8384
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19628 7041 19656 7278
rect 19614 7032 19670 7041
rect 19614 6967 19670 6976
rect 19430 6896 19486 6905
rect 19430 6831 19486 6840
rect 19628 6798 19656 6967
rect 19616 6792 19668 6798
rect 19444 6740 19616 6746
rect 19444 6734 19668 6740
rect 19996 6746 20024 8434
rect 20088 7313 20116 9318
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 20074 7304 20130 7313
rect 20074 7239 20130 7248
rect 19248 6724 19300 6730
rect 19248 6666 19300 6672
rect 19444 6718 19656 6734
rect 19996 6718 20116 6746
rect 20180 6730 20208 8910
rect 20272 8809 20300 11319
rect 20364 10996 20392 11478
rect 20456 11150 20484 12378
rect 20444 11144 20496 11150
rect 20444 11086 20496 11092
rect 20364 10968 20484 10996
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 20364 9897 20392 9998
rect 20350 9888 20406 9897
rect 20350 9823 20406 9832
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 20258 8800 20314 8809
rect 20258 8735 20314 8744
rect 20272 7342 20300 8735
rect 20260 7336 20312 7342
rect 20260 7278 20312 7284
rect 19154 6352 19210 6361
rect 19154 6287 19156 6296
rect 19208 6287 19210 6296
rect 19156 6258 19208 6264
rect 19260 6186 19288 6666
rect 19338 6488 19394 6497
rect 19338 6423 19394 6432
rect 19352 6390 19380 6423
rect 19340 6384 19392 6390
rect 19340 6326 19392 6332
rect 19444 6254 19472 6718
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 19248 6180 19300 6186
rect 19248 6122 19300 6128
rect 19432 5772 19484 5778
rect 19432 5714 19484 5720
rect 19064 5092 19116 5098
rect 19064 5034 19116 5040
rect 19248 5024 19300 5030
rect 19248 4966 19300 4972
rect 19156 4208 19208 4214
rect 18892 4134 19104 4162
rect 19260 4196 19288 4966
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19208 4168 19288 4196
rect 19156 4150 19208 4156
rect 18432 4100 18828 4128
rect 17868 4072 17920 4078
rect 17868 4014 17920 4020
rect 17316 2372 17368 2378
rect 17316 2314 17368 2320
rect 17684 2372 17736 2378
rect 17684 2314 17736 2320
rect 17328 2106 17356 2314
rect 18432 2310 18460 4100
rect 18800 4060 18828 4100
rect 18880 4072 18932 4078
rect 18800 4032 18880 4060
rect 18524 4010 18736 4026
rect 18972 4072 19024 4078
rect 18880 4014 18932 4020
rect 18970 4040 18972 4049
rect 19024 4040 19026 4049
rect 18512 4004 18736 4010
rect 18564 3998 18736 4004
rect 18512 3946 18564 3952
rect 18604 3936 18656 3942
rect 18604 3878 18656 3884
rect 18708 3890 18736 3998
rect 18970 3975 19026 3984
rect 18616 3466 18644 3878
rect 18708 3862 19012 3890
rect 18788 3664 18840 3670
rect 18788 3606 18840 3612
rect 18604 3460 18656 3466
rect 18604 3402 18656 3408
rect 18696 3392 18748 3398
rect 18696 3334 18748 3340
rect 18604 2508 18656 2514
rect 18604 2450 18656 2456
rect 18420 2304 18472 2310
rect 18420 2246 18472 2252
rect 17316 2100 17368 2106
rect 17316 2042 17368 2048
rect 18616 2038 18644 2450
rect 18604 2032 18656 2038
rect 18604 1974 18656 1980
rect 18708 800 18736 3334
rect 18800 3126 18828 3606
rect 18984 3466 19012 3862
rect 18972 3460 19024 3466
rect 18972 3402 19024 3408
rect 18788 3120 18840 3126
rect 18788 3062 18840 3068
rect 19076 2774 19104 4134
rect 19352 3942 19380 4762
rect 19340 3936 19392 3942
rect 19154 3904 19210 3913
rect 19340 3878 19392 3884
rect 19154 3839 19210 3848
rect 19168 2990 19196 3839
rect 19352 3194 19380 3878
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19352 3058 19380 3130
rect 19444 3108 19472 5714
rect 19996 5642 20024 6598
rect 20088 6390 20116 6718
rect 20168 6724 20220 6730
rect 20168 6666 20220 6672
rect 20076 6384 20128 6390
rect 20076 6326 20128 6332
rect 20258 5944 20314 5953
rect 20258 5879 20260 5888
rect 20312 5879 20314 5888
rect 20260 5850 20312 5856
rect 20364 5658 20392 9522
rect 20456 7177 20484 10968
rect 20548 8906 20576 13126
rect 20626 13016 20682 13025
rect 20626 12951 20682 12960
rect 20640 11286 20668 12951
rect 20732 12434 20760 14486
rect 20824 14346 20852 16390
rect 20812 14340 20864 14346
rect 20812 14282 20864 14288
rect 20810 13968 20866 13977
rect 20810 13903 20812 13912
rect 20864 13903 20866 13912
rect 20812 13874 20864 13880
rect 20824 12986 20852 13874
rect 20916 13326 20944 16662
rect 21008 15434 21036 16934
rect 21364 16516 21416 16522
rect 21364 16458 21416 16464
rect 20996 15428 21048 15434
rect 20996 15370 21048 15376
rect 21376 15162 21404 16458
rect 21364 15156 21416 15162
rect 21364 15098 21416 15104
rect 21270 15056 21326 15065
rect 21192 15000 21270 15008
rect 21192 14980 21272 15000
rect 20996 14340 21048 14346
rect 20996 14282 21048 14288
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 20812 12980 20864 12986
rect 20812 12922 20864 12928
rect 21008 12782 21036 14282
rect 21192 13938 21220 14980
rect 21324 14991 21326 15000
rect 21364 15020 21416 15026
rect 21272 14962 21324 14968
rect 21364 14962 21416 14968
rect 21376 14618 21404 14962
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21364 14272 21416 14278
rect 21364 14214 21416 14220
rect 21180 13932 21232 13938
rect 21180 13874 21232 13880
rect 21088 13252 21140 13258
rect 21088 13194 21140 13200
rect 20996 12776 21048 12782
rect 20996 12718 21048 12724
rect 20732 12406 20944 12434
rect 20720 12368 20772 12374
rect 20718 12336 20720 12345
rect 20772 12336 20774 12345
rect 20718 12271 20774 12280
rect 20812 12096 20864 12102
rect 20812 12038 20864 12044
rect 20824 11830 20852 12038
rect 20812 11824 20864 11830
rect 20812 11766 20864 11772
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 20732 11082 20760 11494
rect 20916 11393 20944 12406
rect 20902 11384 20958 11393
rect 20902 11319 20958 11328
rect 20720 11076 20772 11082
rect 20720 11018 20772 11024
rect 20904 11008 20956 11014
rect 20904 10950 20956 10956
rect 20916 10130 20944 10950
rect 20996 10668 21048 10674
rect 20996 10610 21048 10616
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 20904 9988 20956 9994
rect 20904 9930 20956 9936
rect 20628 9920 20680 9926
rect 20628 9862 20680 9868
rect 20536 8900 20588 8906
rect 20536 8842 20588 8848
rect 20640 8786 20668 9862
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 20732 9110 20760 9318
rect 20720 9104 20772 9110
rect 20720 9046 20772 9052
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 20548 8758 20668 8786
rect 20442 7168 20498 7177
rect 20442 7103 20498 7112
rect 19984 5636 20036 5642
rect 19984 5578 20036 5584
rect 20180 5630 20392 5658
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 20180 5370 20208 5630
rect 20352 5568 20404 5574
rect 20352 5510 20404 5516
rect 20168 5364 20220 5370
rect 20168 5306 20220 5312
rect 19616 5160 19668 5166
rect 19616 5102 19668 5108
rect 19628 4826 19656 5102
rect 20074 4856 20130 4865
rect 19616 4820 19668 4826
rect 20074 4791 20130 4800
rect 19616 4762 19668 4768
rect 20088 4690 20116 4791
rect 20076 4684 20128 4690
rect 20076 4626 20128 4632
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19892 4004 19944 4010
rect 19892 3946 19944 3952
rect 19904 3602 19932 3946
rect 19892 3596 19944 3602
rect 19892 3538 19944 3544
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19800 3188 19852 3194
rect 19800 3130 19852 3136
rect 19616 3120 19668 3126
rect 19444 3080 19616 3108
rect 19616 3062 19668 3068
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19156 2984 19208 2990
rect 19156 2926 19208 2932
rect 18892 2746 19104 2774
rect 19352 2774 19380 2994
rect 19812 2854 19840 3130
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 19352 2746 19472 2774
rect 18892 2038 18920 2746
rect 19444 2446 19472 2746
rect 20180 2666 20208 5306
rect 20364 4078 20392 5510
rect 20456 4162 20484 7103
rect 20548 5574 20576 8758
rect 20732 8430 20760 8842
rect 20824 8498 20852 9318
rect 20916 8906 20944 9930
rect 21008 9722 21036 10610
rect 20996 9716 21048 9722
rect 20996 9658 21048 9664
rect 21100 9042 21128 13194
rect 21192 9450 21220 13874
rect 21272 13864 21324 13870
rect 21272 13806 21324 13812
rect 21284 11354 21312 13806
rect 21376 12918 21404 14214
rect 21364 12912 21416 12918
rect 21364 12854 21416 12860
rect 21364 12232 21416 12238
rect 21364 12174 21416 12180
rect 21376 11762 21404 12174
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 21272 11076 21324 11082
rect 21272 11018 21324 11024
rect 21284 10810 21312 11018
rect 21376 11014 21404 11290
rect 21364 11008 21416 11014
rect 21364 10950 21416 10956
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 21272 10600 21324 10606
rect 21272 10542 21324 10548
rect 21180 9444 21232 9450
rect 21180 9386 21232 9392
rect 21284 9382 21312 10542
rect 21364 10260 21416 10266
rect 21364 10202 21416 10208
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21088 9036 21140 9042
rect 21088 8978 21140 8984
rect 20996 8968 21048 8974
rect 20996 8910 21048 8916
rect 20904 8900 20956 8906
rect 20904 8842 20956 8848
rect 20812 8492 20864 8498
rect 20812 8434 20864 8440
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20718 8256 20774 8265
rect 20718 8191 20774 8200
rect 20732 7750 20760 8191
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20640 6458 20668 6802
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 20640 5914 20668 6394
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20536 5568 20588 5574
rect 20536 5510 20588 5516
rect 20640 5166 20668 5850
rect 20628 5160 20680 5166
rect 20628 5102 20680 5108
rect 20640 4826 20668 5102
rect 20628 4820 20680 4826
rect 20628 4762 20680 4768
rect 20534 4720 20590 4729
rect 20534 4655 20590 4664
rect 20548 4282 20576 4655
rect 20640 4282 20668 4762
rect 20536 4276 20588 4282
rect 20536 4218 20588 4224
rect 20628 4276 20680 4282
rect 20628 4218 20680 4224
rect 20456 4134 20576 4162
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 20352 3936 20404 3942
rect 20352 3878 20404 3884
rect 20364 3670 20392 3878
rect 20352 3664 20404 3670
rect 20352 3606 20404 3612
rect 20444 3528 20496 3534
rect 20444 3470 20496 3476
rect 20456 2854 20484 3470
rect 20548 2938 20576 4134
rect 20640 3602 20668 4218
rect 20824 4078 20852 8434
rect 20904 8424 20956 8430
rect 21008 8412 21036 8910
rect 21178 8528 21234 8537
rect 21178 8463 21180 8472
rect 21232 8463 21234 8472
rect 21180 8434 21232 8440
rect 20956 8384 21036 8412
rect 20904 8366 20956 8372
rect 20916 6118 20944 8366
rect 21088 8016 21140 8022
rect 21088 7958 21140 7964
rect 21100 7750 21128 7958
rect 21272 7812 21324 7818
rect 21272 7754 21324 7760
rect 21088 7744 21140 7750
rect 21088 7686 21140 7692
rect 21100 7002 21128 7686
rect 21284 7585 21312 7754
rect 21270 7576 21326 7585
rect 21270 7511 21326 7520
rect 21180 7404 21232 7410
rect 21180 7346 21232 7352
rect 21088 6996 21140 7002
rect 21088 6938 21140 6944
rect 21192 6866 21220 7346
rect 21272 7200 21324 7206
rect 21272 7142 21324 7148
rect 21284 7002 21312 7142
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 21180 6860 21232 6866
rect 21180 6802 21232 6808
rect 20904 6112 20956 6118
rect 20904 6054 20956 6060
rect 20916 5778 20944 6054
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 21272 5704 21324 5710
rect 21272 5646 21324 5652
rect 21284 5545 21312 5646
rect 21270 5536 21326 5545
rect 21270 5471 21326 5480
rect 21376 5030 21404 10202
rect 21468 9994 21496 17002
rect 21548 16584 21600 16590
rect 21548 16526 21600 16532
rect 21560 16250 21588 16526
rect 21548 16244 21600 16250
rect 21548 16186 21600 16192
rect 21548 15428 21600 15434
rect 21548 15370 21600 15376
rect 21560 12646 21588 15370
rect 21548 12640 21600 12646
rect 21548 12582 21600 12588
rect 21546 11928 21602 11937
rect 21546 11863 21602 11872
rect 21560 11762 21588 11863
rect 21548 11756 21600 11762
rect 21548 11698 21600 11704
rect 21652 10810 21680 17614
rect 22388 17134 22416 17682
rect 22376 17128 22428 17134
rect 22376 17070 22428 17076
rect 22836 17128 22888 17134
rect 22836 17070 22888 17076
rect 22192 16992 22244 16998
rect 22192 16934 22244 16940
rect 22652 16992 22704 16998
rect 22652 16934 22704 16940
rect 22204 16250 22232 16934
rect 22560 16652 22612 16658
rect 22560 16594 22612 16600
rect 22192 16244 22244 16250
rect 22192 16186 22244 16192
rect 22006 16144 22062 16153
rect 22006 16079 22008 16088
rect 22060 16079 22062 16088
rect 22008 16050 22060 16056
rect 22100 15972 22152 15978
rect 22100 15914 22152 15920
rect 21914 15600 21970 15609
rect 21914 15535 21970 15544
rect 21928 15502 21956 15535
rect 21916 15496 21968 15502
rect 21916 15438 21968 15444
rect 21916 14952 21968 14958
rect 21916 14894 21968 14900
rect 22112 14940 22140 15914
rect 22376 15088 22428 15094
rect 22376 15030 22428 15036
rect 22468 15088 22520 15094
rect 22468 15030 22520 15036
rect 22388 14958 22416 15030
rect 22192 14952 22244 14958
rect 22112 14912 22192 14940
rect 21928 14618 21956 14894
rect 22008 14884 22060 14890
rect 22008 14826 22060 14832
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 22020 14550 22048 14826
rect 22008 14544 22060 14550
rect 22008 14486 22060 14492
rect 22112 14226 22140 14912
rect 22192 14894 22244 14900
rect 22376 14952 22428 14958
rect 22376 14894 22428 14900
rect 22376 14340 22428 14346
rect 22376 14282 22428 14288
rect 21928 14198 22140 14226
rect 21824 13864 21876 13870
rect 21824 13806 21876 13812
rect 21732 13796 21784 13802
rect 21732 13738 21784 13744
rect 21744 13705 21772 13738
rect 21730 13696 21786 13705
rect 21730 13631 21786 13640
rect 21730 13560 21786 13569
rect 21730 13495 21732 13504
rect 21784 13495 21786 13504
rect 21732 13466 21784 13472
rect 21732 12912 21784 12918
rect 21732 12854 21784 12860
rect 21744 12170 21772 12854
rect 21836 12434 21864 13806
rect 21928 13394 21956 14198
rect 22008 13728 22060 13734
rect 22388 13705 22416 14282
rect 22008 13670 22060 13676
rect 22374 13696 22430 13705
rect 22020 13530 22048 13670
rect 22374 13631 22430 13640
rect 22008 13524 22060 13530
rect 22008 13466 22060 13472
rect 21916 13388 21968 13394
rect 21916 13330 21968 13336
rect 22284 12776 22336 12782
rect 22282 12744 22284 12753
rect 22336 12744 22338 12753
rect 22282 12679 22338 12688
rect 21836 12406 21956 12434
rect 21732 12164 21784 12170
rect 21732 12106 21784 12112
rect 21824 11756 21876 11762
rect 21824 11698 21876 11704
rect 21640 10804 21692 10810
rect 21640 10746 21692 10752
rect 21652 10690 21680 10746
rect 21560 10662 21680 10690
rect 21456 9988 21508 9994
rect 21456 9930 21508 9936
rect 21560 9602 21588 10662
rect 21640 10600 21692 10606
rect 21640 10542 21692 10548
rect 21652 10130 21680 10542
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 21652 9761 21680 10066
rect 21638 9752 21694 9761
rect 21638 9687 21694 9696
rect 21468 9574 21588 9602
rect 21652 9586 21680 9687
rect 21640 9580 21692 9586
rect 21468 5030 21496 9574
rect 21640 9522 21692 9528
rect 21548 9444 21600 9450
rect 21548 9386 21600 9392
rect 21560 7721 21588 9386
rect 21652 9042 21680 9522
rect 21730 9344 21786 9353
rect 21730 9279 21786 9288
rect 21640 9036 21692 9042
rect 21640 8978 21692 8984
rect 21652 8498 21680 8978
rect 21744 8838 21772 9279
rect 21732 8832 21784 8838
rect 21732 8774 21784 8780
rect 21640 8492 21692 8498
rect 21640 8434 21692 8440
rect 21652 7954 21680 8434
rect 21836 8242 21864 11698
rect 21928 11082 21956 12406
rect 22284 12232 22336 12238
rect 22284 12174 22336 12180
rect 22100 11688 22152 11694
rect 22100 11630 22152 11636
rect 22112 11218 22140 11630
rect 22296 11218 22324 12174
rect 22376 11824 22428 11830
rect 22376 11766 22428 11772
rect 22388 11286 22416 11766
rect 22376 11280 22428 11286
rect 22376 11222 22428 11228
rect 22100 11212 22152 11218
rect 22100 11154 22152 11160
rect 22284 11212 22336 11218
rect 22284 11154 22336 11160
rect 21916 11076 21968 11082
rect 21916 11018 21968 11024
rect 22284 11076 22336 11082
rect 22284 11018 22336 11024
rect 22296 10130 22324 11018
rect 22284 10124 22336 10130
rect 22284 10066 22336 10072
rect 21916 9988 21968 9994
rect 21916 9930 21968 9936
rect 21744 8214 21864 8242
rect 21640 7948 21692 7954
rect 21640 7890 21692 7896
rect 21546 7712 21602 7721
rect 21546 7647 21602 7656
rect 21652 7410 21680 7890
rect 21744 7818 21772 8214
rect 21822 8120 21878 8129
rect 21822 8055 21824 8064
rect 21876 8055 21878 8064
rect 21824 8026 21876 8032
rect 21732 7812 21784 7818
rect 21732 7754 21784 7760
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 21744 6254 21772 7754
rect 21928 6866 21956 9930
rect 22192 9648 22244 9654
rect 22190 9616 22192 9625
rect 22244 9616 22246 9625
rect 22480 9602 22508 15030
rect 22572 12356 22600 16594
rect 22664 16522 22692 16934
rect 22652 16516 22704 16522
rect 22652 16458 22704 16464
rect 22664 12434 22692 16458
rect 22848 15484 22876 17070
rect 23032 16522 23060 19110
rect 23020 16516 23072 16522
rect 23020 16458 23072 16464
rect 23124 15570 23152 19654
rect 23756 19168 23808 19174
rect 23756 19110 23808 19116
rect 23480 18624 23532 18630
rect 23480 18566 23532 18572
rect 23388 18216 23440 18222
rect 23388 18158 23440 18164
rect 23296 18080 23348 18086
rect 23296 18022 23348 18028
rect 23308 17882 23336 18022
rect 23296 17876 23348 17882
rect 23296 17818 23348 17824
rect 23400 17762 23428 18158
rect 23204 17740 23256 17746
rect 23204 17682 23256 17688
rect 23308 17734 23428 17762
rect 23216 16794 23244 17682
rect 23204 16788 23256 16794
rect 23204 16730 23256 16736
rect 23204 16040 23256 16046
rect 23204 15982 23256 15988
rect 23216 15910 23244 15982
rect 23204 15904 23256 15910
rect 23204 15846 23256 15852
rect 23112 15564 23164 15570
rect 23112 15506 23164 15512
rect 22756 15456 22876 15484
rect 22928 15496 22980 15502
rect 22756 12986 22784 15456
rect 22980 15456 23060 15484
rect 22928 15438 22980 15444
rect 22928 15360 22980 15366
rect 22928 15302 22980 15308
rect 22836 14952 22888 14958
rect 22836 14894 22888 14900
rect 22848 14385 22876 14894
rect 22834 14376 22890 14385
rect 22940 14346 22968 15302
rect 23032 14822 23060 15456
rect 23020 14816 23072 14822
rect 23020 14758 23072 14764
rect 23124 14482 23152 15506
rect 23216 15473 23244 15846
rect 23202 15464 23258 15473
rect 23202 15399 23258 15408
rect 23112 14476 23164 14482
rect 23112 14418 23164 14424
rect 22834 14311 22890 14320
rect 22928 14340 22980 14346
rect 22744 12980 22796 12986
rect 22744 12922 22796 12928
rect 22664 12406 22784 12434
rect 22572 12328 22692 12356
rect 22560 11620 22612 11626
rect 22560 11562 22612 11568
rect 22572 11286 22600 11562
rect 22560 11280 22612 11286
rect 22560 11222 22612 11228
rect 22664 11132 22692 12328
rect 22190 9551 22246 9560
rect 22296 9574 22508 9602
rect 22572 11104 22692 11132
rect 22054 9500 22106 9506
rect 22190 9480 22246 9489
rect 22106 9448 22190 9466
rect 22054 9442 22190 9448
rect 22066 9438 22190 9442
rect 22190 9415 22246 9424
rect 22008 9376 22060 9382
rect 22008 9318 22060 9324
rect 22020 8362 22048 9318
rect 22296 9110 22324 9574
rect 22376 9512 22428 9518
rect 22376 9454 22428 9460
rect 22284 9104 22336 9110
rect 22284 9046 22336 9052
rect 22284 8832 22336 8838
rect 22282 8800 22284 8809
rect 22336 8800 22338 8809
rect 22282 8735 22338 8744
rect 22284 8424 22336 8430
rect 22284 8366 22336 8372
rect 22008 8356 22060 8362
rect 22008 8298 22060 8304
rect 22296 8129 22324 8366
rect 22388 8294 22416 9454
rect 22572 8786 22600 11104
rect 22650 9616 22706 9625
rect 22650 9551 22706 9560
rect 22664 9518 22692 9551
rect 22652 9512 22704 9518
rect 22652 9454 22704 9460
rect 22756 9382 22784 12406
rect 22848 10470 22876 14311
rect 22928 14282 22980 14288
rect 23124 14006 23152 14418
rect 23112 14000 23164 14006
rect 23112 13942 23164 13948
rect 23018 13424 23074 13433
rect 23018 13359 23020 13368
rect 23072 13359 23074 13368
rect 23020 13330 23072 13336
rect 22926 13152 22982 13161
rect 22926 13087 22982 13096
rect 22940 12918 22968 13087
rect 22928 12912 22980 12918
rect 22928 12854 22980 12860
rect 23110 12880 23166 12889
rect 23110 12815 23166 12824
rect 22928 12640 22980 12646
rect 22928 12582 22980 12588
rect 22940 12288 22968 12582
rect 22940 12260 23060 12288
rect 22928 12164 22980 12170
rect 22928 12106 22980 12112
rect 22836 10464 22888 10470
rect 22836 10406 22888 10412
rect 22744 9376 22796 9382
rect 22744 9318 22796 9324
rect 22480 8758 22600 8786
rect 22376 8288 22428 8294
rect 22376 8230 22428 8236
rect 22282 8120 22338 8129
rect 22008 8084 22060 8090
rect 22480 8106 22508 8758
rect 22560 8628 22612 8634
rect 22560 8570 22612 8576
rect 22572 8514 22600 8570
rect 22572 8486 22692 8514
rect 22664 8430 22692 8486
rect 22652 8424 22704 8430
rect 22558 8392 22614 8401
rect 22652 8366 22704 8372
rect 22558 8327 22614 8336
rect 22338 8078 22508 8106
rect 22282 8055 22338 8064
rect 22008 8026 22060 8032
rect 22020 7546 22048 8026
rect 22192 7744 22244 7750
rect 22190 7712 22192 7721
rect 22244 7712 22246 7721
rect 22190 7647 22246 7656
rect 22008 7540 22060 7546
rect 22008 7482 22060 7488
rect 22296 6905 22324 8055
rect 22572 7478 22600 8327
rect 22560 7472 22612 7478
rect 22560 7414 22612 7420
rect 22376 7336 22428 7342
rect 22376 7278 22428 7284
rect 22652 7336 22704 7342
rect 22652 7278 22704 7284
rect 22388 7177 22416 7278
rect 22374 7168 22430 7177
rect 22374 7103 22430 7112
rect 22468 6928 22520 6934
rect 22098 6896 22154 6905
rect 21916 6860 21968 6866
rect 22282 6896 22338 6905
rect 22154 6854 22232 6882
rect 22098 6831 22154 6840
rect 21916 6802 21968 6808
rect 21732 6248 21784 6254
rect 21732 6190 21784 6196
rect 22204 5681 22232 6854
rect 22468 6870 22520 6876
rect 22282 6831 22338 6840
rect 22284 6316 22336 6322
rect 22284 6258 22336 6264
rect 22190 5672 22246 5681
rect 22190 5607 22246 5616
rect 21824 5160 21876 5166
rect 22204 5148 22232 5607
rect 22296 5409 22324 6258
rect 22282 5400 22338 5409
rect 22282 5335 22338 5344
rect 22376 5296 22428 5302
rect 22376 5238 22428 5244
rect 22388 5166 22416 5238
rect 22284 5160 22336 5166
rect 22204 5120 22284 5148
rect 21824 5102 21876 5108
rect 21364 5024 21416 5030
rect 21364 4966 21416 4972
rect 21456 5024 21508 5030
rect 21456 4966 21508 4972
rect 21376 4842 21404 4966
rect 21180 4820 21232 4826
rect 21180 4762 21232 4768
rect 21284 4814 21404 4842
rect 21192 4622 21220 4762
rect 21180 4616 21232 4622
rect 21180 4558 21232 4564
rect 21284 4146 21312 4814
rect 21468 4706 21496 4966
rect 21376 4678 21496 4706
rect 21836 4690 21864 5102
rect 21928 5098 22140 5114
rect 22284 5102 22336 5108
rect 22376 5160 22428 5166
rect 22376 5102 22428 5108
rect 21916 5092 22140 5098
rect 21968 5086 22140 5092
rect 21916 5034 21968 5040
rect 22112 4978 22140 5086
rect 22480 4978 22508 6870
rect 22560 6180 22612 6186
rect 22560 6122 22612 6128
rect 22572 6089 22600 6122
rect 22558 6080 22614 6089
rect 22558 6015 22614 6024
rect 22112 4950 22508 4978
rect 21824 4684 21876 4690
rect 21272 4140 21324 4146
rect 21272 4082 21324 4088
rect 20812 4072 20864 4078
rect 20812 4014 20864 4020
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 21376 3466 21404 4678
rect 21824 4626 21876 4632
rect 22664 4570 22692 7278
rect 22848 7177 22876 10406
rect 22834 7168 22890 7177
rect 22834 7103 22890 7112
rect 21456 4548 21508 4554
rect 21456 4490 21508 4496
rect 22388 4542 22692 4570
rect 21468 4282 21496 4490
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 21456 4276 21508 4282
rect 21456 4218 21508 4224
rect 22112 4078 22140 4422
rect 22192 4208 22244 4214
rect 22192 4150 22244 4156
rect 22100 4072 22152 4078
rect 22100 4014 22152 4020
rect 21180 3460 21232 3466
rect 21180 3402 21232 3408
rect 21364 3460 21416 3466
rect 21364 3402 21416 3408
rect 21192 3233 21220 3402
rect 21916 3392 21968 3398
rect 21916 3334 21968 3340
rect 21178 3224 21234 3233
rect 21178 3159 21234 3168
rect 20548 2922 20760 2938
rect 20548 2916 20772 2922
rect 20548 2910 20720 2916
rect 20720 2858 20772 2864
rect 20444 2848 20496 2854
rect 20444 2790 20496 2796
rect 20088 2638 20208 2666
rect 20088 2496 20116 2638
rect 19904 2468 20116 2496
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19904 2310 19932 2468
rect 19984 2372 20036 2378
rect 19984 2314 20036 2320
rect 21364 2372 21416 2378
rect 21364 2314 21416 2320
rect 21456 2372 21508 2378
rect 21456 2314 21508 2320
rect 19892 2304 19944 2310
rect 19892 2246 19944 2252
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 18880 2032 18932 2038
rect 18880 1974 18932 1980
rect 19996 800 20024 2314
rect 21376 1834 21404 2314
rect 21468 2038 21496 2314
rect 21456 2032 21508 2038
rect 21456 1974 21508 1980
rect 21364 1828 21416 1834
rect 21364 1770 21416 1776
rect 21928 800 21956 3334
rect 22006 2680 22062 2689
rect 22006 2615 22008 2624
rect 22060 2615 22062 2624
rect 22008 2586 22060 2592
rect 22204 2106 22232 4150
rect 22388 4010 22416 4542
rect 22940 4185 22968 12106
rect 23032 11830 23060 12260
rect 23020 11824 23072 11830
rect 23020 11766 23072 11772
rect 23124 5914 23152 12815
rect 23308 12730 23336 17734
rect 23492 17610 23520 18566
rect 23768 18290 23796 19110
rect 23756 18284 23808 18290
rect 23756 18226 23808 18232
rect 23768 17746 23796 18226
rect 24032 18080 24084 18086
rect 24032 18022 24084 18028
rect 23756 17740 23808 17746
rect 23756 17682 23808 17688
rect 23480 17604 23532 17610
rect 23480 17546 23532 17552
rect 23388 17128 23440 17134
rect 23388 17070 23440 17076
rect 23400 16454 23428 17070
rect 23388 16448 23440 16454
rect 23388 16390 23440 16396
rect 24044 16182 24072 18022
rect 23572 16176 23624 16182
rect 23572 16118 23624 16124
rect 24032 16176 24084 16182
rect 24032 16118 24084 16124
rect 23480 15972 23532 15978
rect 23480 15914 23532 15920
rect 23388 15564 23440 15570
rect 23388 15506 23440 15512
rect 23400 15337 23428 15506
rect 23386 15328 23442 15337
rect 23386 15263 23442 15272
rect 23400 14482 23428 15263
rect 23388 14476 23440 14482
rect 23388 14418 23440 14424
rect 23386 14104 23442 14113
rect 23386 14039 23442 14048
rect 23400 14006 23428 14039
rect 23388 14000 23440 14006
rect 23388 13942 23440 13948
rect 23388 13864 23440 13870
rect 23388 13806 23440 13812
rect 23400 13462 23428 13806
rect 23388 13456 23440 13462
rect 23388 13398 23440 13404
rect 23400 12850 23428 13398
rect 23492 13190 23520 15914
rect 23584 15570 23612 16118
rect 23756 16040 23808 16046
rect 23808 15988 23980 15994
rect 23756 15982 23980 15988
rect 23768 15966 23980 15982
rect 23664 15904 23716 15910
rect 23664 15846 23716 15852
rect 23572 15564 23624 15570
rect 23572 15506 23624 15512
rect 23584 15094 23612 15506
rect 23572 15088 23624 15094
rect 23572 15030 23624 15036
rect 23480 13184 23532 13190
rect 23480 13126 23532 13132
rect 23492 12918 23520 13126
rect 23480 12912 23532 12918
rect 23480 12854 23532 12860
rect 23388 12844 23440 12850
rect 23388 12786 23440 12792
rect 23216 12702 23336 12730
rect 23388 12708 23440 12714
rect 23216 12170 23244 12702
rect 23388 12650 23440 12656
rect 23296 12368 23348 12374
rect 23296 12310 23348 12316
rect 23308 12209 23336 12310
rect 23400 12306 23428 12650
rect 23676 12374 23704 15846
rect 23952 15706 23980 15966
rect 23940 15700 23992 15706
rect 23940 15642 23992 15648
rect 23754 15328 23810 15337
rect 23754 15263 23810 15272
rect 23664 12368 23716 12374
rect 23664 12310 23716 12316
rect 23388 12300 23440 12306
rect 23388 12242 23440 12248
rect 23572 12300 23624 12306
rect 23572 12242 23624 12248
rect 23294 12200 23350 12209
rect 23204 12164 23256 12170
rect 23294 12135 23350 12144
rect 23478 12200 23534 12209
rect 23478 12135 23480 12144
rect 23204 12106 23256 12112
rect 23202 11792 23258 11801
rect 23202 11727 23204 11736
rect 23256 11727 23258 11736
rect 23204 11698 23256 11704
rect 23308 10266 23336 12135
rect 23532 12135 23534 12144
rect 23480 12106 23532 12112
rect 23584 11694 23612 12242
rect 23664 12164 23716 12170
rect 23664 12106 23716 12112
rect 23676 11898 23704 12106
rect 23664 11892 23716 11898
rect 23664 11834 23716 11840
rect 23572 11688 23624 11694
rect 23572 11630 23624 11636
rect 23388 11620 23440 11626
rect 23388 11562 23440 11568
rect 23400 11014 23428 11562
rect 23480 11552 23532 11558
rect 23480 11494 23532 11500
rect 23492 11082 23520 11494
rect 23570 11248 23626 11257
rect 23570 11183 23626 11192
rect 23480 11076 23532 11082
rect 23480 11018 23532 11024
rect 23388 11008 23440 11014
rect 23388 10950 23440 10956
rect 23296 10260 23348 10266
rect 23296 10202 23348 10208
rect 23308 9926 23336 10202
rect 23296 9920 23348 9926
rect 23296 9862 23348 9868
rect 23388 9920 23440 9926
rect 23388 9862 23440 9868
rect 23294 9480 23350 9489
rect 23294 9415 23296 9424
rect 23348 9415 23350 9424
rect 23296 9386 23348 9392
rect 23400 9382 23428 9862
rect 23388 9376 23440 9382
rect 23388 9318 23440 9324
rect 23204 8900 23256 8906
rect 23204 8842 23256 8848
rect 23216 8022 23244 8842
rect 23296 8356 23348 8362
rect 23296 8298 23348 8304
rect 23204 8016 23256 8022
rect 23204 7958 23256 7964
rect 23204 6792 23256 6798
rect 23204 6734 23256 6740
rect 23112 5908 23164 5914
rect 23112 5850 23164 5856
rect 23124 4554 23152 5850
rect 23216 5574 23244 6734
rect 23204 5568 23256 5574
rect 23204 5510 23256 5516
rect 23202 4720 23258 4729
rect 23202 4655 23258 4664
rect 23216 4554 23244 4655
rect 23112 4548 23164 4554
rect 23112 4490 23164 4496
rect 23204 4548 23256 4554
rect 23204 4490 23256 4496
rect 22926 4176 22982 4185
rect 22926 4111 22982 4120
rect 22376 4004 22428 4010
rect 22376 3946 22428 3952
rect 22940 3466 22968 4111
rect 23308 3890 23336 8298
rect 23386 7712 23442 7721
rect 23386 7647 23442 7656
rect 23400 7410 23428 7647
rect 23388 7404 23440 7410
rect 23388 7346 23440 7352
rect 23584 6254 23612 11183
rect 23768 10606 23796 15263
rect 23848 14816 23900 14822
rect 23848 14758 23900 14764
rect 23860 12434 23888 14758
rect 23940 14612 23992 14618
rect 23940 14554 23992 14560
rect 23952 14006 23980 14554
rect 24032 14272 24084 14278
rect 24032 14214 24084 14220
rect 23940 14000 23992 14006
rect 23940 13942 23992 13948
rect 24044 13938 24072 14214
rect 24032 13932 24084 13938
rect 24032 13874 24084 13880
rect 24032 13796 24084 13802
rect 24032 13738 24084 13744
rect 23940 13388 23992 13394
rect 23940 13330 23992 13336
rect 23952 12646 23980 13330
rect 24044 13258 24072 13738
rect 24136 13394 24164 24074
rect 24860 24064 24912 24070
rect 24860 24006 24912 24012
rect 24492 19304 24544 19310
rect 24492 19246 24544 19252
rect 24400 19236 24452 19242
rect 24400 19178 24452 19184
rect 24216 18760 24268 18766
rect 24216 18702 24268 18708
rect 24228 18426 24256 18702
rect 24216 18420 24268 18426
rect 24216 18362 24268 18368
rect 24228 15337 24256 18362
rect 24412 17649 24440 19178
rect 24398 17640 24454 17649
rect 24308 17604 24360 17610
rect 24398 17575 24454 17584
rect 24308 17546 24360 17552
rect 24320 17134 24348 17546
rect 24412 17202 24440 17575
rect 24400 17196 24452 17202
rect 24400 17138 24452 17144
rect 24308 17128 24360 17134
rect 24308 17070 24360 17076
rect 24214 15328 24270 15337
rect 24214 15263 24270 15272
rect 24320 13841 24348 17070
rect 24412 16028 24440 17138
rect 24504 16182 24532 19246
rect 24584 18624 24636 18630
rect 24584 18566 24636 18572
rect 24596 18290 24624 18566
rect 24584 18284 24636 18290
rect 24584 18226 24636 18232
rect 24872 16658 24900 24006
rect 25044 18148 25096 18154
rect 25044 18090 25096 18096
rect 25056 17610 25084 18090
rect 25136 18080 25188 18086
rect 25136 18022 25188 18028
rect 25044 17604 25096 17610
rect 25044 17546 25096 17552
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 25044 16652 25096 16658
rect 25044 16594 25096 16600
rect 24584 16516 24636 16522
rect 24584 16458 24636 16464
rect 24492 16176 24544 16182
rect 24492 16118 24544 16124
rect 24412 16000 24532 16028
rect 24400 15156 24452 15162
rect 24400 15098 24452 15104
rect 24412 14890 24440 15098
rect 24400 14884 24452 14890
rect 24400 14826 24452 14832
rect 24306 13832 24362 13841
rect 24306 13767 24362 13776
rect 24124 13388 24176 13394
rect 24124 13330 24176 13336
rect 24032 13252 24084 13258
rect 24032 13194 24084 13200
rect 24124 13184 24176 13190
rect 24124 13126 24176 13132
rect 24136 12918 24164 13126
rect 24124 12912 24176 12918
rect 24124 12854 24176 12860
rect 23940 12640 23992 12646
rect 23940 12582 23992 12588
rect 23860 12406 24072 12434
rect 23940 11824 23992 11830
rect 23940 11766 23992 11772
rect 23756 10600 23808 10606
rect 23756 10542 23808 10548
rect 23768 9382 23796 10542
rect 23952 9674 23980 11766
rect 24044 11665 24072 12406
rect 24030 11656 24086 11665
rect 24030 11591 24086 11600
rect 23860 9646 23980 9674
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23664 8424 23716 8430
rect 23664 8366 23716 8372
rect 23676 6798 23704 8366
rect 23756 7880 23808 7886
rect 23756 7822 23808 7828
rect 23664 6792 23716 6798
rect 23664 6734 23716 6740
rect 23664 6656 23716 6662
rect 23664 6598 23716 6604
rect 23572 6248 23624 6254
rect 23572 6190 23624 6196
rect 23388 5840 23440 5846
rect 23388 5782 23440 5788
rect 23400 5642 23428 5782
rect 23388 5636 23440 5642
rect 23388 5578 23440 5584
rect 23584 5250 23612 6190
rect 23676 5642 23704 6598
rect 23664 5636 23716 5642
rect 23664 5578 23716 5584
rect 23584 5222 23704 5250
rect 23572 5092 23624 5098
rect 23572 5034 23624 5040
rect 23480 5024 23532 5030
rect 23480 4966 23532 4972
rect 23492 4622 23520 4966
rect 23584 4826 23612 5034
rect 23572 4820 23624 4826
rect 23572 4762 23624 4768
rect 23480 4616 23532 4622
rect 23480 4558 23532 4564
rect 23480 4072 23532 4078
rect 23478 4040 23480 4049
rect 23532 4040 23534 4049
rect 23478 3975 23534 3984
rect 23216 3862 23336 3890
rect 23216 3534 23244 3862
rect 23296 3732 23348 3738
rect 23296 3674 23348 3680
rect 23204 3528 23256 3534
rect 23204 3470 23256 3476
rect 22928 3460 22980 3466
rect 22928 3402 22980 3408
rect 22466 3360 22522 3369
rect 22466 3295 22522 3304
rect 22480 3126 22508 3295
rect 23308 3126 23336 3674
rect 22468 3120 22520 3126
rect 22468 3062 22520 3068
rect 23296 3120 23348 3126
rect 23296 3062 23348 3068
rect 23386 3088 23442 3097
rect 23386 3023 23442 3032
rect 23400 2990 23428 3023
rect 23388 2984 23440 2990
rect 23388 2926 23440 2932
rect 23676 2774 23704 5222
rect 23768 5030 23796 7822
rect 23860 7546 23888 9646
rect 24044 9568 24072 11591
rect 24216 9648 24268 9654
rect 24216 9590 24268 9596
rect 23952 9540 24072 9568
rect 24124 9580 24176 9586
rect 23952 8430 23980 9540
rect 24124 9522 24176 9528
rect 24136 9382 24164 9522
rect 24124 9376 24176 9382
rect 24124 9318 24176 9324
rect 24136 8786 24164 9318
rect 24044 8758 24164 8786
rect 23940 8424 23992 8430
rect 23940 8366 23992 8372
rect 24044 7954 24072 8758
rect 24124 8628 24176 8634
rect 24124 8570 24176 8576
rect 24032 7948 24084 7954
rect 24032 7890 24084 7896
rect 24136 7750 24164 8570
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 23848 7540 23900 7546
rect 23848 7482 23900 7488
rect 24228 7478 24256 9590
rect 24320 9466 24348 13767
rect 24412 12434 24440 14826
rect 24504 14396 24532 16000
rect 24596 15638 24624 16458
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 24584 15632 24636 15638
rect 24584 15574 24636 15580
rect 24780 15366 24808 15982
rect 24952 15428 25004 15434
rect 24952 15370 25004 15376
rect 24768 15360 24820 15366
rect 24768 15302 24820 15308
rect 24780 15094 24808 15302
rect 24964 15162 24992 15370
rect 25056 15314 25084 16594
rect 25148 15434 25176 18022
rect 25240 17610 25268 25094
rect 25884 21690 25912 37198
rect 27080 37126 27108 39200
rect 27436 37256 27488 37262
rect 27436 37198 27488 37204
rect 27068 37120 27120 37126
rect 27068 37062 27120 37068
rect 27448 30938 27476 37198
rect 28368 37126 28396 39200
rect 30300 37210 30328 39200
rect 30472 37256 30524 37262
rect 30300 37182 30420 37210
rect 30472 37198 30524 37204
rect 30840 37256 30892 37262
rect 30840 37198 30892 37204
rect 30392 37126 30420 37182
rect 28356 37120 28408 37126
rect 28356 37062 28408 37068
rect 30380 37120 30432 37126
rect 30380 37062 30432 37068
rect 30484 35290 30512 37198
rect 30472 35284 30524 35290
rect 30472 35226 30524 35232
rect 29644 35080 29696 35086
rect 29644 35022 29696 35028
rect 29656 32434 29684 35022
rect 29644 32428 29696 32434
rect 29644 32370 29696 32376
rect 27436 30932 27488 30938
rect 27436 30874 27488 30880
rect 29276 30592 29328 30598
rect 29276 30534 29328 30540
rect 26424 26784 26476 26790
rect 26424 26726 26476 26732
rect 25872 21684 25924 21690
rect 25872 21626 25924 21632
rect 25964 18624 26016 18630
rect 25964 18566 26016 18572
rect 25872 17808 25924 17814
rect 25872 17750 25924 17756
rect 25228 17604 25280 17610
rect 25228 17546 25280 17552
rect 25240 17116 25268 17546
rect 25412 17536 25464 17542
rect 25412 17478 25464 17484
rect 25424 17270 25452 17478
rect 25412 17264 25464 17270
rect 25412 17206 25464 17212
rect 25320 17128 25372 17134
rect 25240 17088 25320 17116
rect 25320 17070 25372 17076
rect 25780 16720 25832 16726
rect 25780 16662 25832 16668
rect 25792 16046 25820 16662
rect 25780 16040 25832 16046
rect 25780 15982 25832 15988
rect 25504 15972 25556 15978
rect 25504 15914 25556 15920
rect 25516 15502 25544 15914
rect 25504 15496 25556 15502
rect 25504 15438 25556 15444
rect 25136 15428 25188 15434
rect 25136 15370 25188 15376
rect 25056 15286 25268 15314
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 24676 15088 24728 15094
rect 24676 15030 24728 15036
rect 24768 15088 24820 15094
rect 24768 15030 24820 15036
rect 24688 14618 24716 15030
rect 24952 14952 25004 14958
rect 24952 14894 25004 14900
rect 25042 14920 25098 14929
rect 24676 14612 24728 14618
rect 24676 14554 24728 14560
rect 24964 14550 24992 14894
rect 25042 14855 25098 14864
rect 25056 14550 25084 14855
rect 24952 14544 25004 14550
rect 24952 14486 25004 14492
rect 25044 14544 25096 14550
rect 25044 14486 25096 14492
rect 24504 14368 24624 14396
rect 24412 12406 24532 12434
rect 24398 10296 24454 10305
rect 24398 10231 24454 10240
rect 24412 9654 24440 10231
rect 24400 9648 24452 9654
rect 24400 9590 24452 9596
rect 24320 9438 24440 9466
rect 24412 9042 24440 9438
rect 24308 9036 24360 9042
rect 24308 8978 24360 8984
rect 24400 9036 24452 9042
rect 24400 8978 24452 8984
rect 24320 8634 24348 8978
rect 24308 8628 24360 8634
rect 24308 8570 24360 8576
rect 24504 8430 24532 12406
rect 24596 11830 24624 14368
rect 24676 13728 24728 13734
rect 24676 13670 24728 13676
rect 24688 12918 24716 13670
rect 24964 13394 24992 14486
rect 25136 14476 25188 14482
rect 25136 14418 25188 14424
rect 25044 13864 25096 13870
rect 25044 13806 25096 13812
rect 24952 13388 25004 13394
rect 24952 13330 25004 13336
rect 24952 13252 25004 13258
rect 24952 13194 25004 13200
rect 24676 12912 24728 12918
rect 24676 12854 24728 12860
rect 24964 12434 24992 13194
rect 25056 12918 25084 13806
rect 25148 13258 25176 14418
rect 25240 13258 25268 15286
rect 25504 14952 25556 14958
rect 25504 14894 25556 14900
rect 25412 14816 25464 14822
rect 25412 14758 25464 14764
rect 25424 14006 25452 14758
rect 25516 14346 25544 14894
rect 25504 14340 25556 14346
rect 25504 14282 25556 14288
rect 25320 14000 25372 14006
rect 25320 13942 25372 13948
rect 25412 14000 25464 14006
rect 25412 13942 25464 13948
rect 25136 13252 25188 13258
rect 25136 13194 25188 13200
rect 25228 13252 25280 13258
rect 25228 13194 25280 13200
rect 25044 12912 25096 12918
rect 25044 12854 25096 12860
rect 24964 12406 25084 12434
rect 24860 12164 24912 12170
rect 24860 12106 24912 12112
rect 24872 11830 24900 12106
rect 24584 11824 24636 11830
rect 24584 11766 24636 11772
rect 24860 11824 24912 11830
rect 24860 11766 24912 11772
rect 24676 11280 24728 11286
rect 24676 11222 24728 11228
rect 24584 11212 24636 11218
rect 24584 11154 24636 11160
rect 24596 9178 24624 11154
rect 24688 9994 24716 11222
rect 24950 11112 25006 11121
rect 24950 11047 25006 11056
rect 24860 10736 24912 10742
rect 24860 10678 24912 10684
rect 24768 10056 24820 10062
rect 24768 9998 24820 10004
rect 24676 9988 24728 9994
rect 24676 9930 24728 9936
rect 24780 9722 24808 9998
rect 24768 9716 24820 9722
rect 24768 9658 24820 9664
rect 24872 9518 24900 10678
rect 24964 9654 24992 11047
rect 25056 10266 25084 12406
rect 25136 12300 25188 12306
rect 25136 12242 25188 12248
rect 25148 12170 25176 12242
rect 25136 12164 25188 12170
rect 25136 12106 25188 12112
rect 25228 12164 25280 12170
rect 25228 12106 25280 12112
rect 25240 11694 25268 12106
rect 25228 11688 25280 11694
rect 25228 11630 25280 11636
rect 25136 10600 25188 10606
rect 25134 10568 25136 10577
rect 25188 10568 25190 10577
rect 25134 10503 25190 10512
rect 25136 10464 25188 10470
rect 25136 10406 25188 10412
rect 25044 10260 25096 10266
rect 25044 10202 25096 10208
rect 25148 10198 25176 10406
rect 25136 10192 25188 10198
rect 25136 10134 25188 10140
rect 25044 9988 25096 9994
rect 25044 9930 25096 9936
rect 24952 9648 25004 9654
rect 24952 9590 25004 9596
rect 24860 9512 24912 9518
rect 24860 9454 24912 9460
rect 24952 9512 25004 9518
rect 24952 9454 25004 9460
rect 24584 9172 24636 9178
rect 24584 9114 24636 9120
rect 24768 9172 24820 9178
rect 24768 9114 24820 9120
rect 24780 8974 24808 9114
rect 24768 8968 24820 8974
rect 24768 8910 24820 8916
rect 24676 8560 24728 8566
rect 24676 8502 24728 8508
rect 24492 8424 24544 8430
rect 24492 8366 24544 8372
rect 24216 7472 24268 7478
rect 24216 7414 24268 7420
rect 24492 6792 24544 6798
rect 24492 6734 24544 6740
rect 23848 6248 23900 6254
rect 23848 6190 23900 6196
rect 23860 5386 23888 6190
rect 24032 5568 24084 5574
rect 24032 5510 24084 5516
rect 24044 5386 24072 5510
rect 23860 5358 24072 5386
rect 23756 5024 23808 5030
rect 23756 4966 23808 4972
rect 23768 3670 23796 4966
rect 23860 4826 23888 5358
rect 24400 5228 24452 5234
rect 24400 5170 24452 5176
rect 23848 4820 23900 4826
rect 23848 4762 23900 4768
rect 23860 4146 23888 4762
rect 24412 4214 24440 5170
rect 24504 4214 24532 6734
rect 24688 5710 24716 8502
rect 24780 8498 24808 8910
rect 24768 8492 24820 8498
rect 24768 8434 24820 8440
rect 24768 8356 24820 8362
rect 24768 8298 24820 8304
rect 24780 8090 24808 8298
rect 24768 8084 24820 8090
rect 24768 8026 24820 8032
rect 24768 6792 24820 6798
rect 24820 6740 24900 6746
rect 24768 6734 24900 6740
rect 24780 6718 24900 6734
rect 24768 6180 24820 6186
rect 24768 6122 24820 6128
rect 24584 5704 24636 5710
rect 24584 5646 24636 5652
rect 24676 5704 24728 5710
rect 24676 5646 24728 5652
rect 24400 4208 24452 4214
rect 24400 4150 24452 4156
rect 24492 4208 24544 4214
rect 24492 4150 24544 4156
rect 23848 4140 23900 4146
rect 23848 4082 23900 4088
rect 23756 3664 23808 3670
rect 23756 3606 23808 3612
rect 23860 3602 23888 4082
rect 23938 3632 23994 3641
rect 23848 3596 23900 3602
rect 23938 3567 23994 3576
rect 23848 3538 23900 3544
rect 23860 3126 23888 3538
rect 23952 3534 23980 3567
rect 23940 3528 23992 3534
rect 23940 3470 23992 3476
rect 23848 3120 23900 3126
rect 23848 3062 23900 3068
rect 23756 2984 23808 2990
rect 23952 2961 23980 3470
rect 24504 2990 24532 4150
rect 24596 3942 24624 5646
rect 24780 5302 24808 6122
rect 24768 5296 24820 5302
rect 24768 5238 24820 5244
rect 24768 5024 24820 5030
rect 24768 4966 24820 4972
rect 24780 4826 24808 4966
rect 24768 4820 24820 4826
rect 24768 4762 24820 4768
rect 24584 3936 24636 3942
rect 24584 3878 24636 3884
rect 24492 2984 24544 2990
rect 23756 2926 23808 2932
rect 23938 2952 23994 2961
rect 23492 2746 23704 2774
rect 23492 2582 23520 2746
rect 23480 2576 23532 2582
rect 23480 2518 23532 2524
rect 23768 2310 23796 2926
rect 24492 2926 24544 2932
rect 23938 2887 23994 2896
rect 24596 2774 24624 3878
rect 24872 2922 24900 6718
rect 24964 6118 24992 9454
rect 25056 8090 25084 9930
rect 25136 8900 25188 8906
rect 25136 8842 25188 8848
rect 25044 8084 25096 8090
rect 25044 8026 25096 8032
rect 25044 7200 25096 7206
rect 25044 7142 25096 7148
rect 25056 6934 25084 7142
rect 25044 6928 25096 6934
rect 25044 6870 25096 6876
rect 25148 6866 25176 8842
rect 25136 6860 25188 6866
rect 25136 6802 25188 6808
rect 25240 6322 25268 11630
rect 25332 10198 25360 13942
rect 25780 13864 25832 13870
rect 25516 13824 25780 13852
rect 25516 12170 25544 13824
rect 25780 13806 25832 13812
rect 25884 13716 25912 17750
rect 25976 17678 26004 18566
rect 25964 17672 26016 17678
rect 25962 17640 25964 17649
rect 26016 17640 26018 17649
rect 25962 17575 26018 17584
rect 26240 17128 26292 17134
rect 26240 17070 26292 17076
rect 26056 17060 26108 17066
rect 26056 17002 26108 17008
rect 26068 16658 26096 17002
rect 26148 16992 26200 16998
rect 26148 16934 26200 16940
rect 26056 16652 26108 16658
rect 26056 16594 26108 16600
rect 26160 16454 26188 16934
rect 26148 16448 26200 16454
rect 26148 16390 26200 16396
rect 26252 16250 26280 17070
rect 26436 16658 26464 26726
rect 28632 21548 28684 21554
rect 28632 21490 28684 21496
rect 26884 18896 26936 18902
rect 26884 18838 26936 18844
rect 26896 18426 26924 18838
rect 26884 18420 26936 18426
rect 26884 18362 26936 18368
rect 27068 17876 27120 17882
rect 27068 17818 27120 17824
rect 26884 17740 26936 17746
rect 26884 17682 26936 17688
rect 26424 16652 26476 16658
rect 26424 16594 26476 16600
rect 26792 16584 26844 16590
rect 26792 16526 26844 16532
rect 26332 16516 26384 16522
rect 26332 16458 26384 16464
rect 26424 16516 26476 16522
rect 26424 16458 26476 16464
rect 26344 16250 26372 16458
rect 26240 16244 26292 16250
rect 26240 16186 26292 16192
rect 26332 16244 26384 16250
rect 26332 16186 26384 16192
rect 25964 16040 26016 16046
rect 25964 15982 26016 15988
rect 25976 15094 26004 15982
rect 26332 15904 26384 15910
rect 26332 15846 26384 15852
rect 26344 15434 26372 15846
rect 26436 15745 26464 16458
rect 26608 16448 26660 16454
rect 26608 16390 26660 16396
rect 26516 16108 26568 16114
rect 26516 16050 26568 16056
rect 26422 15736 26478 15745
rect 26422 15671 26478 15680
rect 26332 15428 26384 15434
rect 26332 15370 26384 15376
rect 26424 15428 26476 15434
rect 26424 15370 26476 15376
rect 26436 15162 26464 15370
rect 26528 15337 26556 16050
rect 26514 15328 26570 15337
rect 26514 15263 26570 15272
rect 26424 15156 26476 15162
rect 26424 15098 26476 15104
rect 25964 15088 26016 15094
rect 25964 15030 26016 15036
rect 26436 14958 26464 15098
rect 26424 14952 26476 14958
rect 26424 14894 26476 14900
rect 26516 14816 26568 14822
rect 26514 14784 26516 14793
rect 26568 14784 26570 14793
rect 26514 14719 26570 14728
rect 26620 14346 26648 16390
rect 26804 16114 26832 16526
rect 26792 16108 26844 16114
rect 26792 16050 26844 16056
rect 26792 15428 26844 15434
rect 26792 15370 26844 15376
rect 26700 14816 26752 14822
rect 26700 14758 26752 14764
rect 25964 14340 26016 14346
rect 25964 14282 26016 14288
rect 26608 14340 26660 14346
rect 26608 14282 26660 14288
rect 25976 14006 26004 14282
rect 25964 14000 26016 14006
rect 25964 13942 26016 13948
rect 25608 13688 25912 13716
rect 25504 12164 25556 12170
rect 25504 12106 25556 12112
rect 25608 11744 25636 13688
rect 25962 13560 26018 13569
rect 25962 13495 26018 13504
rect 25976 13462 26004 13495
rect 25780 13456 25832 13462
rect 25780 13398 25832 13404
rect 25964 13456 26016 13462
rect 25964 13398 26016 13404
rect 25688 13252 25740 13258
rect 25688 13194 25740 13200
rect 25700 12850 25728 13194
rect 25792 12918 25820 13398
rect 26056 13388 26108 13394
rect 26056 13330 26108 13336
rect 25870 13016 25926 13025
rect 25870 12951 25872 12960
rect 25924 12951 25926 12960
rect 25872 12922 25924 12928
rect 25780 12912 25832 12918
rect 25780 12854 25832 12860
rect 26068 12850 26096 13330
rect 26712 13190 26740 14758
rect 26804 13326 26832 15370
rect 26896 13938 26924 17682
rect 27080 17542 27108 17818
rect 27068 17536 27120 17542
rect 27068 17478 27120 17484
rect 27080 17202 27108 17478
rect 27344 17332 27396 17338
rect 27344 17274 27396 17280
rect 27160 17264 27212 17270
rect 27160 17206 27212 17212
rect 27068 17196 27120 17202
rect 27068 17138 27120 17144
rect 26976 15564 27028 15570
rect 26976 15506 27028 15512
rect 26988 14414 27016 15506
rect 26976 14408 27028 14414
rect 26976 14350 27028 14356
rect 26884 13932 26936 13938
rect 26884 13874 26936 13880
rect 26988 13410 27016 14350
rect 27080 14278 27108 17138
rect 27172 16114 27200 17206
rect 27356 16658 27384 17274
rect 27804 17060 27856 17066
rect 27804 17002 27856 17008
rect 27344 16652 27396 16658
rect 27344 16594 27396 16600
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 27252 15496 27304 15502
rect 27252 15438 27304 15444
rect 27068 14272 27120 14278
rect 27068 14214 27120 14220
rect 27264 13870 27292 15438
rect 27356 15026 27384 16594
rect 27436 15700 27488 15706
rect 27436 15642 27488 15648
rect 27344 15020 27396 15026
rect 27344 14962 27396 14968
rect 27344 13932 27396 13938
rect 27344 13874 27396 13880
rect 27252 13864 27304 13870
rect 27252 13806 27304 13812
rect 27252 13728 27304 13734
rect 27066 13696 27122 13705
rect 27252 13670 27304 13676
rect 27066 13631 27122 13640
rect 27080 13530 27108 13631
rect 27068 13524 27120 13530
rect 27068 13466 27120 13472
rect 26988 13382 27108 13410
rect 26792 13320 26844 13326
rect 26792 13262 26844 13268
rect 26976 13320 27028 13326
rect 26976 13262 27028 13268
rect 26700 13184 26752 13190
rect 26700 13126 26752 13132
rect 25688 12844 25740 12850
rect 25688 12786 25740 12792
rect 26056 12844 26108 12850
rect 26056 12786 26108 12792
rect 25700 12753 25728 12786
rect 25686 12744 25742 12753
rect 25686 12679 25742 12688
rect 25780 12436 25832 12442
rect 25780 12378 25832 12384
rect 25608 11716 25728 11744
rect 25504 11688 25556 11694
rect 25504 11630 25556 11636
rect 25516 10588 25544 11630
rect 25700 10606 25728 11716
rect 25792 11218 25820 12378
rect 26068 11937 26096 12786
rect 26804 12434 26832 13262
rect 26988 12889 27016 13262
rect 27080 13190 27108 13382
rect 27068 13184 27120 13190
rect 27264 13161 27292 13670
rect 27356 13530 27384 13874
rect 27344 13524 27396 13530
rect 27344 13466 27396 13472
rect 27068 13126 27120 13132
rect 27250 13152 27306 13161
rect 27250 13087 27306 13096
rect 26974 12880 27030 12889
rect 26974 12815 27030 12824
rect 26620 12406 26832 12434
rect 26620 12238 26648 12406
rect 27448 12374 27476 15642
rect 27712 15360 27764 15366
rect 27712 15302 27764 15308
rect 27526 15056 27582 15065
rect 27526 14991 27528 15000
rect 27580 14991 27582 15000
rect 27528 14962 27580 14968
rect 27528 14408 27580 14414
rect 27526 14376 27528 14385
rect 27580 14376 27582 14385
rect 27526 14311 27582 14320
rect 27528 14272 27580 14278
rect 27528 14214 27580 14220
rect 27540 13938 27568 14214
rect 27724 14113 27752 15302
rect 27710 14104 27766 14113
rect 27710 14039 27766 14048
rect 27528 13932 27580 13938
rect 27528 13874 27580 13880
rect 27620 13796 27672 13802
rect 27620 13738 27672 13744
rect 27528 13252 27580 13258
rect 27528 13194 27580 13200
rect 27540 12986 27568 13194
rect 27528 12980 27580 12986
rect 27528 12922 27580 12928
rect 27526 12744 27582 12753
rect 27526 12679 27582 12688
rect 27540 12646 27568 12679
rect 27528 12640 27580 12646
rect 27528 12582 27580 12588
rect 27632 12442 27660 13738
rect 27816 13258 27844 17002
rect 28448 16448 28500 16454
rect 28448 16390 28500 16396
rect 27986 16280 28042 16289
rect 27986 16215 28042 16224
rect 28000 16114 28028 16215
rect 28460 16114 28488 16390
rect 27988 16108 28040 16114
rect 27988 16050 28040 16056
rect 28448 16108 28500 16114
rect 28448 16050 28500 16056
rect 28000 13920 28028 16050
rect 28172 15360 28224 15366
rect 28172 15302 28224 15308
rect 28080 13932 28132 13938
rect 28000 13892 28080 13920
rect 28080 13874 28132 13880
rect 27896 13864 27948 13870
rect 27896 13806 27948 13812
rect 27804 13252 27856 13258
rect 27804 13194 27856 13200
rect 27712 12708 27764 12714
rect 27712 12650 27764 12656
rect 27620 12436 27672 12442
rect 27620 12378 27672 12384
rect 27436 12368 27488 12374
rect 27436 12310 27488 12316
rect 27448 12238 27476 12310
rect 26608 12232 26660 12238
rect 26608 12174 26660 12180
rect 27436 12232 27488 12238
rect 27436 12174 27488 12180
rect 27620 12232 27672 12238
rect 27724 12209 27752 12650
rect 27620 12174 27672 12180
rect 27710 12200 27766 12209
rect 26054 11928 26110 11937
rect 26054 11863 26110 11872
rect 26332 11824 26384 11830
rect 26330 11792 26332 11801
rect 26384 11792 26386 11801
rect 26330 11727 26386 11736
rect 25872 11552 25924 11558
rect 25872 11494 25924 11500
rect 25780 11212 25832 11218
rect 25780 11154 25832 11160
rect 25780 10736 25832 10742
rect 25780 10678 25832 10684
rect 25596 10600 25648 10606
rect 25516 10560 25596 10588
rect 25596 10542 25648 10548
rect 25688 10600 25740 10606
rect 25688 10542 25740 10548
rect 25320 10192 25372 10198
rect 25320 10134 25372 10140
rect 25608 8090 25636 10542
rect 25792 10305 25820 10678
rect 25778 10296 25834 10305
rect 25778 10231 25834 10240
rect 25884 9874 25912 11494
rect 26620 11218 26648 12174
rect 27356 11886 27568 11914
rect 27356 11762 27384 11886
rect 27344 11756 27396 11762
rect 27344 11698 27396 11704
rect 27436 11756 27488 11762
rect 27436 11698 27488 11704
rect 27448 11642 27476 11698
rect 27172 11614 27476 11642
rect 27068 11552 27120 11558
rect 27172 11540 27200 11614
rect 27540 11558 27568 11886
rect 27120 11512 27200 11540
rect 27252 11552 27304 11558
rect 27068 11494 27120 11500
rect 27528 11552 27580 11558
rect 27252 11494 27304 11500
rect 27356 11512 27528 11540
rect 27264 11354 27292 11494
rect 27252 11348 27304 11354
rect 27252 11290 27304 11296
rect 26424 11212 26476 11218
rect 26608 11212 26660 11218
rect 26476 11172 26556 11200
rect 26424 11154 26476 11160
rect 26146 11112 26202 11121
rect 26146 11047 26148 11056
rect 26200 11047 26202 11056
rect 26332 11076 26384 11082
rect 26148 11018 26200 11024
rect 26384 11036 26464 11064
rect 26332 11018 26384 11024
rect 26054 10704 26110 10713
rect 26054 10639 26110 10648
rect 25964 10260 26016 10266
rect 25964 10202 26016 10208
rect 25976 9994 26004 10202
rect 25964 9988 26016 9994
rect 25964 9930 26016 9936
rect 25884 9846 26004 9874
rect 25872 9036 25924 9042
rect 25872 8978 25924 8984
rect 25884 8566 25912 8978
rect 25872 8560 25924 8566
rect 25872 8502 25924 8508
rect 25976 8498 26004 9846
rect 25780 8492 25832 8498
rect 25780 8434 25832 8440
rect 25964 8492 26016 8498
rect 25964 8434 26016 8440
rect 25596 8084 25648 8090
rect 25596 8026 25648 8032
rect 25686 7848 25742 7857
rect 25686 7783 25742 7792
rect 25700 7546 25728 7783
rect 25320 7540 25372 7546
rect 25320 7482 25372 7488
rect 25688 7540 25740 7546
rect 25688 7482 25740 7488
rect 25228 6316 25280 6322
rect 25228 6258 25280 6264
rect 24952 6112 25004 6118
rect 24952 6054 25004 6060
rect 25332 5794 25360 7482
rect 25596 7472 25648 7478
rect 25596 7414 25648 7420
rect 25608 6934 25636 7414
rect 25688 7336 25740 7342
rect 25688 7278 25740 7284
rect 25596 6928 25648 6934
rect 25410 6896 25466 6905
rect 25596 6870 25648 6876
rect 25410 6831 25466 6840
rect 25424 6118 25452 6831
rect 25700 6798 25728 7278
rect 25792 7041 25820 8434
rect 26068 8090 26096 10639
rect 26148 9988 26200 9994
rect 26148 9930 26200 9936
rect 26160 8650 26188 9930
rect 26240 9920 26292 9926
rect 26240 9862 26292 9868
rect 26252 9654 26280 9862
rect 26436 9654 26464 11036
rect 26528 10577 26556 11172
rect 26608 11154 26660 11160
rect 27068 10600 27120 10606
rect 26514 10568 26570 10577
rect 27068 10542 27120 10548
rect 26514 10503 26570 10512
rect 26528 10180 26556 10503
rect 26608 10192 26660 10198
rect 26528 10152 26608 10180
rect 26608 10134 26660 10140
rect 27080 9994 27108 10542
rect 27068 9988 27120 9994
rect 27068 9930 27120 9936
rect 26240 9648 26292 9654
rect 26240 9590 26292 9596
rect 26424 9648 26476 9654
rect 26424 9590 26476 9596
rect 26332 9580 26384 9586
rect 26332 9522 26384 9528
rect 26344 9217 26372 9522
rect 27080 9518 27108 9930
rect 27068 9512 27120 9518
rect 27068 9454 27120 9460
rect 27160 9512 27212 9518
rect 27160 9454 27212 9460
rect 26330 9208 26386 9217
rect 26330 9143 26386 9152
rect 26792 9104 26844 9110
rect 26792 9046 26844 9052
rect 26516 8900 26568 8906
rect 26516 8842 26568 8848
rect 26160 8622 26280 8650
rect 26252 8294 26280 8622
rect 26424 8492 26476 8498
rect 26424 8434 26476 8440
rect 26240 8288 26292 8294
rect 26240 8230 26292 8236
rect 26056 8084 26108 8090
rect 26056 8026 26108 8032
rect 26330 7984 26386 7993
rect 26330 7919 26386 7928
rect 26240 7880 26292 7886
rect 26240 7822 26292 7828
rect 26252 7410 26280 7822
rect 26344 7546 26372 7919
rect 26332 7540 26384 7546
rect 26332 7482 26384 7488
rect 26436 7410 26464 8434
rect 26240 7404 26292 7410
rect 26240 7346 26292 7352
rect 26424 7404 26476 7410
rect 26424 7346 26476 7352
rect 25962 7168 26018 7177
rect 25962 7103 26018 7112
rect 25778 7032 25834 7041
rect 25778 6967 25834 6976
rect 25596 6792 25648 6798
rect 25596 6734 25648 6740
rect 25688 6792 25740 6798
rect 25688 6734 25740 6740
rect 25412 6112 25464 6118
rect 25412 6054 25464 6060
rect 25240 5766 25360 5794
rect 25044 5228 25096 5234
rect 25044 5170 25096 5176
rect 24860 2916 24912 2922
rect 24860 2858 24912 2864
rect 24412 2746 24624 2774
rect 24412 2514 24440 2746
rect 25056 2514 25084 5170
rect 25240 2990 25268 5766
rect 25412 5636 25464 5642
rect 25412 5578 25464 5584
rect 25424 5166 25452 5578
rect 25504 5568 25556 5574
rect 25504 5510 25556 5516
rect 25412 5160 25464 5166
rect 25412 5102 25464 5108
rect 25516 4162 25544 5510
rect 25608 4554 25636 6734
rect 25700 6254 25728 6734
rect 25688 6248 25740 6254
rect 25688 6190 25740 6196
rect 25872 5908 25924 5914
rect 25872 5850 25924 5856
rect 25884 5710 25912 5850
rect 25872 5704 25924 5710
rect 25872 5646 25924 5652
rect 25976 5574 26004 7103
rect 26528 6662 26556 8842
rect 26608 8832 26660 8838
rect 26608 8774 26660 8780
rect 26516 6656 26568 6662
rect 26516 6598 26568 6604
rect 26514 6488 26570 6497
rect 26514 6423 26570 6432
rect 26528 5681 26556 6423
rect 26514 5672 26570 5681
rect 26514 5607 26570 5616
rect 25780 5568 25832 5574
rect 25780 5510 25832 5516
rect 25964 5568 26016 5574
rect 25964 5510 26016 5516
rect 25792 5370 25820 5510
rect 25780 5364 25832 5370
rect 25780 5306 25832 5312
rect 26424 5024 26476 5030
rect 26424 4966 26476 4972
rect 26240 4820 26292 4826
rect 26240 4762 26292 4768
rect 25596 4548 25648 4554
rect 25596 4490 25648 4496
rect 25516 4146 25820 4162
rect 25516 4140 25832 4146
rect 25516 4134 25780 4140
rect 25780 4082 25832 4088
rect 25504 3596 25556 3602
rect 25504 3538 25556 3544
rect 25516 3126 25544 3538
rect 25504 3120 25556 3126
rect 25504 3062 25556 3068
rect 26252 3058 26280 4762
rect 26332 4548 26384 4554
rect 26332 4490 26384 4496
rect 26344 4078 26372 4490
rect 26436 4282 26464 4966
rect 26424 4276 26476 4282
rect 26424 4218 26476 4224
rect 26332 4072 26384 4078
rect 26424 4072 26476 4078
rect 26332 4014 26384 4020
rect 26422 4040 26424 4049
rect 26476 4040 26478 4049
rect 26528 4010 26556 5607
rect 26422 3975 26478 3984
rect 26516 4004 26568 4010
rect 26516 3946 26568 3952
rect 26620 3670 26648 8774
rect 26804 8090 26832 9046
rect 27172 9042 27200 9454
rect 27160 9036 27212 9042
rect 27160 8978 27212 8984
rect 27252 8628 27304 8634
rect 27252 8570 27304 8576
rect 26884 8288 26936 8294
rect 26884 8230 26936 8236
rect 26792 8084 26844 8090
rect 26792 8026 26844 8032
rect 26896 7886 26924 8230
rect 27264 7886 27292 8570
rect 26884 7880 26936 7886
rect 26884 7822 26936 7828
rect 27252 7880 27304 7886
rect 27252 7822 27304 7828
rect 26896 6798 26924 7822
rect 27252 7744 27304 7750
rect 27252 7686 27304 7692
rect 27264 7546 27292 7686
rect 27252 7540 27304 7546
rect 27252 7482 27304 7488
rect 27252 7200 27304 7206
rect 27252 7142 27304 7148
rect 27264 7002 27292 7142
rect 27252 6996 27304 7002
rect 27252 6938 27304 6944
rect 26884 6792 26936 6798
rect 26884 6734 26936 6740
rect 27356 6746 27384 11512
rect 27528 11494 27580 11500
rect 27632 11257 27660 12174
rect 27710 12135 27766 12144
rect 27618 11248 27674 11257
rect 27618 11183 27674 11192
rect 27620 11008 27672 11014
rect 27620 10950 27672 10956
rect 27528 10056 27580 10062
rect 27528 9998 27580 10004
rect 27540 9897 27568 9998
rect 27526 9888 27582 9897
rect 27526 9823 27582 9832
rect 27436 9716 27488 9722
rect 27436 9658 27488 9664
rect 27448 7954 27476 9658
rect 27632 9654 27660 10950
rect 27712 10532 27764 10538
rect 27712 10474 27764 10480
rect 27528 9648 27580 9654
rect 27526 9616 27528 9625
rect 27620 9648 27672 9654
rect 27580 9616 27582 9625
rect 27620 9590 27672 9596
rect 27526 9551 27582 9560
rect 27528 9444 27580 9450
rect 27528 9386 27580 9392
rect 27620 9444 27672 9450
rect 27620 9386 27672 9392
rect 27540 8090 27568 9386
rect 27632 8498 27660 9386
rect 27724 9110 27752 10474
rect 27816 9518 27844 13194
rect 27908 12306 27936 13806
rect 28184 13258 28212 15302
rect 28460 14890 28488 16050
rect 28540 15564 28592 15570
rect 28540 15506 28592 15512
rect 28552 15366 28580 15506
rect 28540 15360 28592 15366
rect 28540 15302 28592 15308
rect 28644 15026 28672 21490
rect 29000 15496 29052 15502
rect 29000 15438 29052 15444
rect 28632 15020 28684 15026
rect 28632 14962 28684 14968
rect 28448 14884 28500 14890
rect 28448 14826 28500 14832
rect 29012 14822 29040 15438
rect 29000 14816 29052 14822
rect 29000 14758 29052 14764
rect 29012 14482 29040 14758
rect 29000 14476 29052 14482
rect 29000 14418 29052 14424
rect 28540 14408 28592 14414
rect 28540 14350 28592 14356
rect 28264 14068 28316 14074
rect 28264 14010 28316 14016
rect 28276 13258 28304 14010
rect 28552 13394 28580 14350
rect 29288 13938 29316 30534
rect 29656 25498 29684 32370
rect 30852 30938 30880 37198
rect 32232 37126 32260 39200
rect 33520 37126 33548 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35452 37330 35480 39200
rect 37186 38856 37242 38865
rect 37186 38791 37242 38800
rect 35440 37324 35492 37330
rect 35440 37266 35492 37272
rect 33600 37256 33652 37262
rect 33600 37198 33652 37204
rect 35808 37256 35860 37262
rect 35808 37198 35860 37204
rect 32220 37120 32272 37126
rect 32220 37062 32272 37068
rect 33508 37120 33560 37126
rect 33508 37062 33560 37068
rect 33612 36922 33640 37198
rect 33600 36916 33652 36922
rect 33600 36858 33652 36864
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35820 36378 35848 37198
rect 37200 36378 37228 38791
rect 37384 36922 37412 39200
rect 38290 37496 38346 37505
rect 38290 37431 38346 37440
rect 38304 37330 38332 37431
rect 38292 37324 38344 37330
rect 38292 37266 38344 37272
rect 37832 37256 37884 37262
rect 37832 37198 37884 37204
rect 37372 36916 37424 36922
rect 37372 36858 37424 36864
rect 37740 36780 37792 36786
rect 37740 36722 37792 36728
rect 35808 36372 35860 36378
rect 35808 36314 35860 36320
rect 37188 36372 37240 36378
rect 37188 36314 37240 36320
rect 36728 36032 36780 36038
rect 36728 35974 36780 35980
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 30840 30932 30892 30938
rect 30840 30874 30892 30880
rect 30564 30728 30616 30734
rect 30564 30670 30616 30676
rect 29644 25492 29696 25498
rect 29644 25434 29696 25440
rect 30576 24138 30604 30670
rect 36740 30054 36768 35974
rect 36728 30048 36780 30054
rect 36728 29990 36780 29996
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 30564 24132 30616 24138
rect 30564 24074 30616 24080
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 37464 21548 37516 21554
rect 37464 21490 37516 21496
rect 37476 21350 37504 21490
rect 37464 21344 37516 21350
rect 37464 21286 37516 21292
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 36636 19372 36688 19378
rect 36636 19314 36688 19320
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35900 17060 35952 17066
rect 35900 17002 35952 17008
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 30288 16516 30340 16522
rect 30288 16458 30340 16464
rect 30196 15972 30248 15978
rect 30196 15914 30248 15920
rect 29644 15020 29696 15026
rect 29644 14962 29696 14968
rect 28724 13932 28776 13938
rect 28724 13874 28776 13880
rect 29276 13932 29328 13938
rect 29276 13874 29328 13880
rect 29460 13932 29512 13938
rect 29460 13874 29512 13880
rect 28632 13456 28684 13462
rect 28632 13398 28684 13404
rect 28540 13388 28592 13394
rect 28540 13330 28592 13336
rect 28172 13252 28224 13258
rect 28172 13194 28224 13200
rect 28264 13252 28316 13258
rect 28264 13194 28316 13200
rect 28644 12850 28672 13398
rect 28736 13394 28764 13874
rect 28724 13388 28776 13394
rect 28724 13330 28776 13336
rect 28632 12844 28684 12850
rect 28632 12786 28684 12792
rect 28724 12776 28776 12782
rect 28724 12718 28776 12724
rect 27896 12300 27948 12306
rect 27896 12242 27948 12248
rect 27988 12232 28040 12238
rect 27988 12174 28040 12180
rect 27896 11824 27948 11830
rect 27896 11766 27948 11772
rect 27908 10606 27936 11766
rect 28000 11150 28028 12174
rect 28356 12096 28408 12102
rect 28356 12038 28408 12044
rect 28368 11286 28396 12038
rect 28448 11756 28500 11762
rect 28448 11698 28500 11704
rect 28460 11665 28488 11698
rect 28446 11656 28502 11665
rect 28446 11591 28502 11600
rect 28356 11280 28408 11286
rect 28356 11222 28408 11228
rect 27988 11144 28040 11150
rect 27988 11086 28040 11092
rect 27896 10600 27948 10606
rect 27896 10542 27948 10548
rect 27908 9518 27936 10542
rect 27804 9512 27856 9518
rect 27804 9454 27856 9460
rect 27896 9512 27948 9518
rect 27896 9454 27948 9460
rect 27712 9104 27764 9110
rect 27712 9046 27764 9052
rect 28000 8922 28028 11086
rect 28264 11008 28316 11014
rect 28264 10950 28316 10956
rect 28276 10742 28304 10950
rect 28264 10736 28316 10742
rect 28264 10678 28316 10684
rect 28356 10532 28408 10538
rect 28356 10474 28408 10480
rect 28264 10192 28316 10198
rect 28264 10134 28316 10140
rect 28172 9648 28224 9654
rect 28172 9590 28224 9596
rect 28184 8974 28212 9590
rect 27816 8894 28028 8922
rect 28172 8968 28224 8974
rect 28172 8910 28224 8916
rect 27620 8492 27672 8498
rect 27620 8434 27672 8440
rect 27528 8084 27580 8090
rect 27528 8026 27580 8032
rect 27436 7948 27488 7954
rect 27436 7890 27488 7896
rect 27436 7744 27488 7750
rect 27434 7712 27436 7721
rect 27488 7712 27490 7721
rect 27434 7647 27490 7656
rect 27528 7404 27580 7410
rect 27528 7346 27580 7352
rect 26698 5944 26754 5953
rect 26698 5879 26754 5888
rect 26712 5778 26740 5879
rect 26700 5772 26752 5778
rect 26700 5714 26752 5720
rect 26896 5234 26924 6734
rect 27252 6724 27304 6730
rect 27356 6718 27476 6746
rect 27252 6666 27304 6672
rect 27264 6322 27292 6666
rect 27344 6656 27396 6662
rect 27344 6598 27396 6604
rect 27252 6316 27304 6322
rect 27252 6258 27304 6264
rect 27356 6186 27384 6598
rect 27344 6180 27396 6186
rect 27344 6122 27396 6128
rect 27448 6118 27476 6718
rect 27436 6112 27488 6118
rect 27436 6054 27488 6060
rect 27066 5808 27122 5817
rect 27066 5743 27122 5752
rect 26884 5228 26936 5234
rect 26884 5170 26936 5176
rect 27080 4622 27108 5743
rect 27158 5536 27214 5545
rect 27158 5471 27214 5480
rect 27172 4758 27200 5471
rect 27250 5400 27306 5409
rect 27448 5386 27476 6054
rect 27540 5914 27568 7346
rect 27816 6497 27844 8894
rect 27988 8628 28040 8634
rect 27988 8570 28040 8576
rect 28172 8628 28224 8634
rect 28172 8570 28224 8576
rect 28000 8498 28028 8570
rect 27988 8492 28040 8498
rect 27988 8434 28040 8440
rect 28184 7886 28212 8570
rect 28080 7880 28132 7886
rect 28080 7822 28132 7828
rect 28172 7880 28224 7886
rect 28172 7822 28224 7828
rect 27894 7576 27950 7585
rect 27894 7511 27950 7520
rect 27908 7478 27936 7511
rect 27896 7472 27948 7478
rect 27896 7414 27948 7420
rect 28092 7410 28120 7822
rect 28080 7404 28132 7410
rect 28080 7346 28132 7352
rect 28092 6798 28120 7346
rect 28080 6792 28132 6798
rect 28080 6734 28132 6740
rect 27988 6656 28040 6662
rect 27988 6598 28040 6604
rect 27802 6488 27858 6497
rect 28000 6458 28028 6598
rect 27802 6423 27858 6432
rect 27988 6452 28040 6458
rect 27988 6394 28040 6400
rect 28092 6338 28120 6734
rect 27816 6322 28120 6338
rect 28184 6322 28212 7822
rect 27804 6316 28120 6322
rect 27856 6310 28120 6316
rect 27804 6258 27856 6264
rect 27896 6180 27948 6186
rect 27896 6122 27948 6128
rect 27908 5914 27936 6122
rect 27528 5908 27580 5914
rect 27528 5850 27580 5856
rect 27896 5908 27948 5914
rect 27896 5850 27948 5856
rect 27250 5335 27252 5344
rect 27304 5335 27306 5344
rect 27356 5358 27476 5386
rect 27252 5306 27304 5312
rect 27160 4752 27212 4758
rect 27160 4694 27212 4700
rect 27068 4616 27120 4622
rect 27068 4558 27120 4564
rect 26976 4480 27028 4486
rect 26976 4422 27028 4428
rect 27068 4480 27120 4486
rect 27068 4422 27120 4428
rect 26988 4282 27016 4422
rect 26976 4276 27028 4282
rect 26976 4218 27028 4224
rect 26424 3664 26476 3670
rect 26424 3606 26476 3612
rect 26608 3664 26660 3670
rect 26608 3606 26660 3612
rect 26240 3052 26292 3058
rect 26240 2994 26292 3000
rect 25228 2984 25280 2990
rect 25228 2926 25280 2932
rect 26252 2774 26280 2994
rect 26252 2746 26372 2774
rect 26344 2514 26372 2746
rect 24400 2508 24452 2514
rect 24400 2450 24452 2456
rect 25044 2508 25096 2514
rect 25044 2450 25096 2456
rect 26332 2508 26384 2514
rect 26332 2450 26384 2456
rect 26436 2378 26464 3606
rect 26792 3528 26844 3534
rect 26792 3470 26844 3476
rect 26514 2680 26570 2689
rect 26514 2615 26570 2624
rect 26528 2582 26556 2615
rect 26516 2576 26568 2582
rect 26516 2518 26568 2524
rect 25596 2372 25648 2378
rect 25596 2314 25648 2320
rect 26424 2372 26476 2378
rect 26424 2314 26476 2320
rect 23756 2304 23808 2310
rect 23756 2246 23808 2252
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 22192 2100 22244 2106
rect 22192 2042 22244 2048
rect 23860 800 23888 2246
rect 25608 1902 25636 2314
rect 25504 1896 25556 1902
rect 25504 1838 25556 1844
rect 25596 1896 25648 1902
rect 25596 1838 25648 1844
rect 25136 1760 25188 1766
rect 25136 1702 25188 1708
rect 25148 800 25176 1702
rect 25516 1630 25544 1838
rect 26804 1698 26832 3470
rect 27080 3097 27108 4422
rect 27356 3534 27384 5358
rect 27540 5234 27568 5850
rect 27908 5522 27936 5850
rect 27724 5494 27936 5522
rect 27528 5228 27580 5234
rect 27448 5188 27528 5216
rect 27448 4622 27476 5188
rect 27528 5170 27580 5176
rect 27526 5128 27582 5137
rect 27526 5063 27582 5072
rect 27436 4616 27488 4622
rect 27436 4558 27488 4564
rect 27436 4004 27488 4010
rect 27436 3946 27488 3952
rect 27344 3528 27396 3534
rect 27344 3470 27396 3476
rect 27066 3088 27122 3097
rect 27448 3058 27476 3946
rect 27540 3534 27568 5063
rect 27724 4826 27752 5494
rect 28092 5234 28120 6310
rect 28172 6316 28224 6322
rect 28172 6258 28224 6264
rect 28184 5710 28212 6258
rect 28172 5704 28224 5710
rect 28172 5646 28224 5652
rect 27988 5228 28040 5234
rect 27988 5170 28040 5176
rect 28080 5228 28132 5234
rect 28080 5170 28132 5176
rect 28000 5114 28028 5170
rect 28184 5114 28212 5646
rect 28000 5086 28212 5114
rect 27712 4820 27764 4826
rect 27712 4762 27764 4768
rect 28000 4146 28028 5086
rect 28172 4616 28224 4622
rect 28172 4558 28224 4564
rect 28184 4146 28212 4558
rect 27988 4140 28040 4146
rect 28172 4140 28224 4146
rect 27988 4082 28040 4088
rect 28092 4100 28172 4128
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 27066 3023 27122 3032
rect 27436 3052 27488 3058
rect 27436 2994 27488 3000
rect 27068 2848 27120 2854
rect 27068 2790 27120 2796
rect 27896 2848 27948 2854
rect 27896 2790 27948 2796
rect 26792 1692 26844 1698
rect 26792 1634 26844 1640
rect 25504 1624 25556 1630
rect 25504 1566 25556 1572
rect 27080 800 27108 2790
rect 27908 2446 27936 2790
rect 28000 2446 28028 4082
rect 28092 3534 28120 4100
rect 28172 4082 28224 4088
rect 28172 3936 28224 3942
rect 28172 3878 28224 3884
rect 28184 3738 28212 3878
rect 28172 3732 28224 3738
rect 28172 3674 28224 3680
rect 28080 3528 28132 3534
rect 28080 3470 28132 3476
rect 28276 3398 28304 10134
rect 28368 9722 28396 10474
rect 28632 9988 28684 9994
rect 28632 9930 28684 9936
rect 28356 9716 28408 9722
rect 28356 9658 28408 9664
rect 28540 9716 28592 9722
rect 28540 9658 28592 9664
rect 28368 3505 28396 9658
rect 28552 9217 28580 9658
rect 28538 9208 28594 9217
rect 28538 9143 28594 9152
rect 28448 7744 28500 7750
rect 28448 7686 28500 7692
rect 28460 4622 28488 7686
rect 28552 5370 28580 9143
rect 28644 8498 28672 9930
rect 28736 9353 28764 12718
rect 29472 12434 29500 13874
rect 29472 12406 29592 12434
rect 28908 12232 28960 12238
rect 28908 12174 28960 12180
rect 28816 10600 28868 10606
rect 28816 10542 28868 10548
rect 28828 9674 28856 10542
rect 28920 10470 28948 12174
rect 29000 10668 29052 10674
rect 29000 10610 29052 10616
rect 28908 10464 28960 10470
rect 28908 10406 28960 10412
rect 29012 10062 29040 10610
rect 29368 10464 29420 10470
rect 29368 10406 29420 10412
rect 29092 10260 29144 10266
rect 29092 10202 29144 10208
rect 29000 10056 29052 10062
rect 29000 9998 29052 10004
rect 28828 9646 28948 9674
rect 28722 9344 28778 9353
rect 28722 9279 28778 9288
rect 28816 8900 28868 8906
rect 28816 8842 28868 8848
rect 28632 8492 28684 8498
rect 28632 8434 28684 8440
rect 28644 7546 28672 8434
rect 28724 8424 28776 8430
rect 28722 8392 28724 8401
rect 28776 8392 28778 8401
rect 28722 8327 28778 8336
rect 28828 7886 28856 8842
rect 28920 8634 28948 9646
rect 29012 9450 29040 9998
rect 29104 9518 29132 10202
rect 29274 10160 29330 10169
rect 29380 10130 29408 10406
rect 29274 10095 29330 10104
rect 29368 10124 29420 10130
rect 29182 10024 29238 10033
rect 29182 9959 29238 9968
rect 29092 9512 29144 9518
rect 29092 9454 29144 9460
rect 29000 9444 29052 9450
rect 29000 9386 29052 9392
rect 29196 8634 29224 9959
rect 28908 8628 28960 8634
rect 28908 8570 28960 8576
rect 29184 8628 29236 8634
rect 29184 8570 29236 8576
rect 28920 8498 28948 8570
rect 28908 8492 28960 8498
rect 28908 8434 28960 8440
rect 29000 8356 29052 8362
rect 29000 8298 29052 8304
rect 29012 8265 29040 8298
rect 28998 8256 29054 8265
rect 28998 8191 29054 8200
rect 28816 7880 28868 7886
rect 28816 7822 28868 7828
rect 28632 7540 28684 7546
rect 28632 7482 28684 7488
rect 28828 7410 28856 7822
rect 29184 7472 29236 7478
rect 29182 7440 29184 7449
rect 29236 7440 29238 7449
rect 28816 7404 28868 7410
rect 29182 7375 29238 7384
rect 28816 7346 28868 7352
rect 29184 7336 29236 7342
rect 29184 7278 29236 7284
rect 29196 6798 29224 7278
rect 29288 6866 29316 10095
rect 29368 10066 29420 10072
rect 29368 9512 29420 9518
rect 29366 9480 29368 9489
rect 29420 9480 29422 9489
rect 29366 9415 29422 9424
rect 29276 6860 29328 6866
rect 29276 6802 29328 6808
rect 29184 6792 29236 6798
rect 29184 6734 29236 6740
rect 28630 6080 28686 6089
rect 28630 6015 28686 6024
rect 28540 5364 28592 5370
rect 28540 5306 28592 5312
rect 28448 4616 28500 4622
rect 28448 4558 28500 4564
rect 28460 4486 28488 4558
rect 28448 4480 28500 4486
rect 28448 4422 28500 4428
rect 28448 3936 28500 3942
rect 28448 3878 28500 3884
rect 28354 3496 28410 3505
rect 28460 3466 28488 3878
rect 28354 3431 28410 3440
rect 28448 3460 28500 3466
rect 28448 3402 28500 3408
rect 28264 3392 28316 3398
rect 28552 3346 28580 5306
rect 28644 4826 28672 6015
rect 29092 5840 29144 5846
rect 29092 5782 29144 5788
rect 28816 5024 28868 5030
rect 28816 4966 28868 4972
rect 28632 4820 28684 4826
rect 28632 4762 28684 4768
rect 28722 4584 28778 4593
rect 28722 4519 28778 4528
rect 28736 3738 28764 4519
rect 28828 4214 28856 4966
rect 28816 4208 28868 4214
rect 28816 4150 28868 4156
rect 29104 4146 29132 5782
rect 29196 5710 29224 6734
rect 29184 5704 29236 5710
rect 29184 5646 29236 5652
rect 29196 4622 29224 5646
rect 29184 4616 29236 4622
rect 29184 4558 29236 4564
rect 29000 4140 29052 4146
rect 29000 4082 29052 4088
rect 29092 4140 29144 4146
rect 29092 4082 29144 4088
rect 28724 3732 28776 3738
rect 28724 3674 28776 3680
rect 28816 3528 28868 3534
rect 28816 3470 28868 3476
rect 28264 3334 28316 3340
rect 28460 3318 28580 3346
rect 28630 3360 28686 3369
rect 28460 3126 28488 3318
rect 28630 3295 28686 3304
rect 28538 3224 28594 3233
rect 28538 3159 28594 3168
rect 28448 3120 28500 3126
rect 28448 3062 28500 3068
rect 28552 3058 28580 3159
rect 28644 3126 28672 3295
rect 28632 3120 28684 3126
rect 28632 3062 28684 3068
rect 28540 3052 28592 3058
rect 28540 2994 28592 3000
rect 28828 3040 28856 3470
rect 29012 3074 29040 4082
rect 29012 3058 29316 3074
rect 28908 3052 28960 3058
rect 28828 3012 28908 3040
rect 28632 2984 28684 2990
rect 28630 2952 28632 2961
rect 28684 2952 28686 2961
rect 28630 2887 28686 2896
rect 28828 2446 28856 3012
rect 29012 3052 29328 3058
rect 29012 3046 29276 3052
rect 28908 2994 28960 3000
rect 29276 2994 29328 3000
rect 28908 2848 28960 2854
rect 28908 2790 28960 2796
rect 29276 2848 29328 2854
rect 29276 2790 29328 2796
rect 27896 2440 27948 2446
rect 27896 2382 27948 2388
rect 27988 2440 28040 2446
rect 27988 2382 28040 2388
rect 28816 2440 28868 2446
rect 28816 2382 28868 2388
rect 28080 2372 28132 2378
rect 28080 2314 28132 2320
rect 28092 1766 28120 2314
rect 28724 2304 28776 2310
rect 28724 2246 28776 2252
rect 28736 2106 28764 2246
rect 28920 2106 28948 2790
rect 29288 2582 29316 2790
rect 29564 2650 29592 12406
rect 29656 6390 29684 14962
rect 29828 13864 29880 13870
rect 29828 13806 29880 13812
rect 29840 12442 29868 13806
rect 29828 12436 29880 12442
rect 29828 12378 29880 12384
rect 30208 11014 30236 15914
rect 30300 12442 30328 16458
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 30932 15360 30984 15366
rect 30932 15302 30984 15308
rect 30288 12436 30340 12442
rect 30288 12378 30340 12384
rect 30748 11620 30800 11626
rect 30748 11562 30800 11568
rect 30196 11008 30248 11014
rect 30196 10950 30248 10956
rect 30196 10056 30248 10062
rect 30196 9998 30248 10004
rect 29920 9988 29972 9994
rect 29920 9930 29972 9936
rect 29932 9586 29960 9930
rect 29920 9580 29972 9586
rect 29920 9522 29972 9528
rect 29828 8560 29880 8566
rect 29828 8502 29880 8508
rect 29840 7546 29868 8502
rect 29932 8294 29960 9522
rect 30208 8974 30236 9998
rect 30760 9178 30788 11562
rect 30748 9172 30800 9178
rect 30748 9114 30800 9120
rect 30564 9036 30616 9042
rect 30564 8978 30616 8984
rect 30196 8968 30248 8974
rect 30196 8910 30248 8916
rect 30286 8936 30342 8945
rect 30286 8871 30342 8880
rect 30012 8492 30064 8498
rect 30012 8434 30064 8440
rect 29920 8288 29972 8294
rect 29920 8230 29972 8236
rect 29828 7540 29880 7546
rect 29828 7482 29880 7488
rect 29644 6384 29696 6390
rect 29644 6326 29696 6332
rect 29932 5386 29960 8230
rect 30024 7886 30052 8434
rect 30300 8090 30328 8871
rect 30288 8084 30340 8090
rect 30288 8026 30340 8032
rect 30012 7880 30064 7886
rect 30012 7822 30064 7828
rect 30288 7880 30340 7886
rect 30288 7822 30340 7828
rect 30024 7410 30052 7822
rect 30012 7404 30064 7410
rect 30012 7346 30064 7352
rect 29840 5358 29960 5386
rect 29840 4146 29868 5358
rect 30024 5234 30052 7346
rect 30300 7342 30328 7822
rect 30288 7336 30340 7342
rect 30288 7278 30340 7284
rect 30470 7304 30526 7313
rect 30470 7239 30472 7248
rect 30524 7239 30526 7248
rect 30472 7210 30524 7216
rect 30380 6180 30432 6186
rect 30380 6122 30432 6128
rect 30392 5574 30420 6122
rect 30380 5568 30432 5574
rect 30380 5510 30432 5516
rect 29920 5228 29972 5234
rect 29920 5170 29972 5176
rect 30012 5228 30064 5234
rect 30012 5170 30064 5176
rect 29828 4140 29880 4146
rect 29828 4082 29880 4088
rect 29932 3534 29960 5170
rect 30024 4214 30052 5170
rect 30392 5098 30420 5510
rect 30380 5092 30432 5098
rect 30380 5034 30432 5040
rect 30380 4276 30432 4282
rect 30380 4218 30432 4224
rect 30012 4208 30064 4214
rect 30012 4150 30064 4156
rect 30024 3602 30052 4150
rect 30288 4140 30340 4146
rect 30288 4082 30340 4088
rect 30012 3596 30064 3602
rect 30012 3538 30064 3544
rect 30300 3534 30328 4082
rect 30392 3738 30420 4218
rect 30576 4146 30604 8978
rect 30840 5568 30892 5574
rect 30840 5510 30892 5516
rect 30564 4140 30616 4146
rect 30564 4082 30616 4088
rect 30380 3732 30432 3738
rect 30380 3674 30432 3680
rect 29920 3528 29972 3534
rect 29920 3470 29972 3476
rect 30288 3528 30340 3534
rect 30288 3470 30340 3476
rect 30300 3058 30328 3470
rect 30472 3392 30524 3398
rect 30472 3334 30524 3340
rect 29736 3052 29788 3058
rect 29736 2994 29788 3000
rect 30288 3052 30340 3058
rect 30288 2994 30340 3000
rect 29552 2644 29604 2650
rect 29552 2586 29604 2592
rect 29276 2576 29328 2582
rect 29276 2518 29328 2524
rect 29748 2446 29776 2994
rect 29920 2848 29972 2854
rect 29920 2790 29972 2796
rect 29826 2544 29882 2553
rect 29826 2479 29828 2488
rect 29880 2479 29882 2488
rect 29828 2450 29880 2456
rect 29736 2440 29788 2446
rect 29932 2417 29960 2790
rect 29736 2382 29788 2388
rect 29918 2408 29974 2417
rect 29918 2343 29974 2352
rect 30288 2304 30340 2310
rect 30288 2246 30340 2252
rect 28724 2100 28776 2106
rect 28724 2042 28776 2048
rect 28908 2100 28960 2106
rect 28908 2042 28960 2048
rect 28080 1760 28132 1766
rect 28080 1702 28132 1708
rect 29000 1760 29052 1766
rect 29000 1702 29052 1708
rect 29012 800 29040 1702
rect 30300 800 30328 2246
rect 30484 1630 30512 3334
rect 30852 2922 30880 5510
rect 30840 2916 30892 2922
rect 30840 2858 30892 2864
rect 30564 2848 30616 2854
rect 30564 2790 30616 2796
rect 30576 1902 30604 2790
rect 30944 2582 30972 15302
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35912 12986 35940 17002
rect 36648 15706 36676 19314
rect 37476 18698 37504 21286
rect 37464 18692 37516 18698
rect 37464 18634 37516 18640
rect 37752 18426 37780 36722
rect 37844 29646 37872 37198
rect 37924 36712 37976 36718
rect 37924 36654 37976 36660
rect 37936 35630 37964 36654
rect 38016 36576 38068 36582
rect 38016 36518 38068 36524
rect 38028 36174 38056 36518
rect 38672 36378 38700 39200
rect 38660 36372 38712 36378
rect 38660 36314 38712 36320
rect 38016 36168 38068 36174
rect 38016 36110 38068 36116
rect 37924 35624 37976 35630
rect 37924 35566 37976 35572
rect 38292 35624 38344 35630
rect 38292 35566 38344 35572
rect 37832 29640 37884 29646
rect 37832 29582 37884 29588
rect 37844 29306 37872 29582
rect 37832 29300 37884 29306
rect 37832 29242 37884 29248
rect 37936 26994 37964 35566
rect 38304 35465 38332 35566
rect 38290 35456 38346 35465
rect 38290 35391 38346 35400
rect 38304 35290 38332 35391
rect 38292 35284 38344 35290
rect 38292 35226 38344 35232
rect 38198 33416 38254 33425
rect 38198 33351 38200 33360
rect 38252 33351 38254 33360
rect 38200 33322 38252 33328
rect 38292 32360 38344 32366
rect 38292 32302 38344 32308
rect 38304 32065 38332 32302
rect 38290 32056 38346 32065
rect 38290 31991 38292 32000
rect 38344 31991 38346 32000
rect 38292 31962 38344 31968
rect 38016 30252 38068 30258
rect 38016 30194 38068 30200
rect 38028 29850 38056 30194
rect 38200 30048 38252 30054
rect 38198 30016 38200 30025
rect 38252 30016 38254 30025
rect 38198 29951 38254 29960
rect 38016 29844 38068 29850
rect 38016 29786 38068 29792
rect 38108 29300 38160 29306
rect 38108 29242 38160 29248
rect 37924 26988 37976 26994
rect 37924 26930 37976 26936
rect 38016 26920 38068 26926
rect 38016 26862 38068 26868
rect 38028 26586 38056 26862
rect 38016 26580 38068 26586
rect 38016 26522 38068 26528
rect 38016 24812 38068 24818
rect 38016 24754 38068 24760
rect 37924 22500 37976 22506
rect 37924 22442 37976 22448
rect 37740 18420 37792 18426
rect 37740 18362 37792 18368
rect 36636 15700 36688 15706
rect 36636 15642 36688 15648
rect 35900 12980 35952 12986
rect 35900 12922 35952 12928
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34796 11008 34848 11014
rect 34796 10950 34848 10956
rect 33692 9376 33744 9382
rect 33692 9318 33744 9324
rect 33048 8968 33100 8974
rect 33048 8910 33100 8916
rect 31022 6352 31078 6361
rect 31022 6287 31078 6296
rect 31036 3534 31064 6287
rect 31114 5264 31170 5273
rect 31114 5199 31170 5208
rect 31128 4010 31156 5199
rect 33060 4826 33088 8910
rect 33140 6248 33192 6254
rect 33140 6190 33192 6196
rect 33048 4820 33100 4826
rect 33048 4762 33100 4768
rect 33060 4622 33088 4762
rect 31208 4616 31260 4622
rect 31208 4558 31260 4564
rect 31852 4616 31904 4622
rect 31852 4558 31904 4564
rect 33048 4616 33100 4622
rect 33048 4558 33100 4564
rect 31220 4146 31248 4558
rect 31208 4140 31260 4146
rect 31208 4082 31260 4088
rect 31116 4004 31168 4010
rect 31116 3946 31168 3952
rect 31760 4004 31812 4010
rect 31760 3946 31812 3952
rect 31772 3670 31800 3946
rect 31760 3664 31812 3670
rect 31760 3606 31812 3612
rect 31864 3534 31892 4558
rect 33060 4146 33088 4558
rect 33048 4140 33100 4146
rect 33048 4082 33100 4088
rect 32496 4072 32548 4078
rect 32496 4014 32548 4020
rect 32508 3534 32536 4014
rect 32954 3632 33010 3641
rect 32954 3567 32956 3576
rect 33008 3567 33010 3576
rect 32956 3538 33008 3544
rect 31024 3528 31076 3534
rect 31024 3470 31076 3476
rect 31852 3528 31904 3534
rect 31852 3470 31904 3476
rect 32496 3528 32548 3534
rect 32496 3470 32548 3476
rect 31300 3460 31352 3466
rect 31300 3402 31352 3408
rect 31024 2984 31076 2990
rect 31022 2952 31024 2961
rect 31076 2952 31078 2961
rect 31022 2887 31078 2896
rect 31208 2848 31260 2854
rect 31208 2790 31260 2796
rect 30932 2576 30984 2582
rect 30932 2518 30984 2524
rect 31220 2038 31248 2790
rect 31312 2650 31340 3402
rect 31760 3392 31812 3398
rect 31760 3334 31812 3340
rect 31300 2644 31352 2650
rect 31300 2586 31352 2592
rect 31312 2446 31340 2586
rect 31300 2440 31352 2446
rect 31300 2382 31352 2388
rect 31208 2032 31260 2038
rect 31208 1974 31260 1980
rect 31772 1970 31800 3334
rect 32508 3058 32536 3470
rect 33152 3058 33180 6190
rect 33600 5092 33652 5098
rect 33600 5034 33652 5040
rect 33612 3398 33640 5034
rect 33600 3392 33652 3398
rect 33600 3334 33652 3340
rect 32496 3052 32548 3058
rect 32496 2994 32548 3000
rect 33140 3052 33192 3058
rect 33140 2994 33192 3000
rect 32312 2848 32364 2854
rect 32312 2790 32364 2796
rect 32324 2446 32352 2790
rect 32312 2440 32364 2446
rect 32312 2382 32364 2388
rect 32220 2372 32272 2378
rect 32220 2314 32272 2320
rect 31760 1964 31812 1970
rect 31760 1906 31812 1912
rect 30564 1896 30616 1902
rect 30564 1838 30616 1844
rect 30472 1624 30524 1630
rect 30472 1566 30524 1572
rect 32232 800 32260 2314
rect 32324 1766 32352 2382
rect 33152 2310 33180 2994
rect 33612 2650 33640 3334
rect 33600 2644 33652 2650
rect 33600 2586 33652 2592
rect 33704 2530 33732 9318
rect 34808 3738 34836 10950
rect 37004 10532 37056 10538
rect 37004 10474 37056 10480
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 37016 9654 37044 10474
rect 37004 9648 37056 9654
rect 37004 9590 37056 9596
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 37936 9178 37964 22442
rect 38028 16182 38056 24754
rect 38120 24410 38148 29242
rect 38198 27976 38254 27985
rect 38198 27911 38200 27920
rect 38252 27911 38254 27920
rect 38200 27882 38252 27888
rect 38292 26920 38344 26926
rect 38292 26862 38344 26868
rect 38304 26625 38332 26862
rect 38290 26616 38346 26625
rect 38290 26551 38292 26560
rect 38344 26551 38346 26560
rect 38292 26522 38344 26528
rect 38200 24608 38252 24614
rect 38198 24576 38200 24585
rect 38252 24576 38254 24585
rect 38198 24511 38254 24520
rect 38108 24404 38160 24410
rect 38108 24346 38160 24352
rect 38200 22636 38252 22642
rect 38200 22578 38252 22584
rect 38212 22545 38240 22578
rect 38198 22536 38254 22545
rect 38198 22471 38254 22480
rect 38200 21344 38252 21350
rect 38200 21286 38252 21292
rect 38212 21185 38240 21286
rect 38198 21176 38254 21185
rect 38198 21111 38254 21120
rect 38200 19168 38252 19174
rect 38198 19136 38200 19145
rect 38252 19136 38254 19145
rect 38198 19071 38254 19080
rect 38200 17196 38252 17202
rect 38200 17138 38252 17144
rect 38212 17105 38240 17138
rect 38198 17096 38254 17105
rect 38198 17031 38254 17040
rect 38016 16176 38068 16182
rect 38016 16118 38068 16124
rect 38200 16108 38252 16114
rect 38200 16050 38252 16056
rect 38014 16008 38070 16017
rect 38014 15943 38016 15952
rect 38068 15943 38070 15952
rect 38016 15914 38068 15920
rect 38212 15745 38240 16050
rect 38198 15736 38254 15745
rect 38198 15671 38254 15680
rect 38200 13932 38252 13938
rect 38200 13874 38252 13880
rect 38212 13705 38240 13874
rect 38198 13696 38254 13705
rect 38198 13631 38254 13640
rect 38016 12436 38068 12442
rect 38016 12378 38068 12384
rect 37924 9172 37976 9178
rect 37924 9114 37976 9120
rect 38028 8566 38056 12378
rect 38200 11756 38252 11762
rect 38200 11698 38252 11704
rect 38212 11665 38240 11698
rect 38198 11656 38254 11665
rect 38198 11591 38254 11600
rect 38200 10668 38252 10674
rect 38200 10610 38252 10616
rect 38212 10305 38240 10610
rect 38198 10296 38254 10305
rect 38198 10231 38254 10240
rect 38016 8560 38068 8566
rect 38016 8502 38068 8508
rect 38200 8492 38252 8498
rect 38200 8434 38252 8440
rect 38212 8265 38240 8434
rect 38198 8256 38254 8265
rect 34934 8188 35242 8197
rect 38198 8191 38254 8200
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 37922 6760 37978 6769
rect 37922 6695 37978 6704
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34796 3732 34848 3738
rect 34796 3674 34848 3680
rect 34060 3392 34112 3398
rect 34060 3334 34112 3340
rect 33612 2502 33732 2530
rect 34072 2514 34100 3334
rect 34336 2984 34388 2990
rect 34336 2926 34388 2932
rect 34060 2508 34112 2514
rect 33612 2310 33640 2502
rect 34060 2450 34112 2456
rect 34348 2446 34376 2926
rect 34808 2446 34836 3674
rect 37936 3670 37964 6695
rect 38200 6316 38252 6322
rect 38200 6258 38252 6264
rect 38212 6225 38240 6258
rect 38198 6216 38254 6225
rect 38198 6151 38254 6160
rect 38016 5160 38068 5166
rect 38016 5102 38068 5108
rect 38292 5160 38344 5166
rect 38292 5102 38344 5108
rect 38028 4690 38056 5102
rect 38304 4865 38332 5102
rect 38290 4856 38346 4865
rect 38290 4791 38292 4800
rect 38344 4791 38346 4800
rect 38292 4762 38344 4768
rect 38016 4684 38068 4690
rect 38016 4626 38068 4632
rect 38016 4004 38068 4010
rect 38016 3946 38068 3952
rect 37924 3664 37976 3670
rect 37924 3606 37976 3612
rect 38028 3058 38056 3946
rect 39304 3460 39356 3466
rect 39304 3402 39356 3408
rect 38016 3052 38068 3058
rect 38016 2994 38068 3000
rect 36636 2916 36688 2922
rect 36636 2858 36688 2864
rect 35440 2848 35492 2854
rect 35440 2790 35492 2796
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34336 2440 34388 2446
rect 34336 2382 34388 2388
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 35452 2378 35480 2790
rect 36648 2446 36676 2858
rect 38200 2848 38252 2854
rect 38198 2816 38200 2825
rect 38252 2816 38254 2825
rect 38198 2751 38254 2760
rect 36636 2440 36688 2446
rect 36636 2382 36688 2388
rect 37464 2440 37516 2446
rect 37464 2382 37516 2388
rect 35440 2372 35492 2378
rect 35440 2314 35492 2320
rect 33140 2304 33192 2310
rect 33140 2246 33192 2252
rect 33600 2304 33652 2310
rect 33600 2246 33652 2252
rect 34152 2304 34204 2310
rect 34152 2246 34204 2252
rect 33612 1834 33640 2246
rect 33600 1828 33652 1834
rect 33600 1770 33652 1776
rect 32312 1760 32364 1766
rect 32312 1702 32364 1708
rect 34164 800 34192 2246
rect 35452 800 35480 2314
rect 37188 2304 37240 2310
rect 37188 2246 37240 2252
rect 37372 2304 37424 2310
rect 37372 2246 37424 2252
rect 37200 1465 37228 2246
rect 37186 1456 37242 1465
rect 37186 1391 37242 1400
rect 37384 800 37412 2246
rect 37476 2106 37504 2382
rect 37464 2100 37516 2106
rect 37464 2042 37516 2048
rect 39316 800 39344 3402
rect 16868 734 17264 762
rect 18694 200 18750 800
rect 19982 200 20038 800
rect 21914 200 21970 800
rect 23846 200 23902 800
rect 25134 200 25190 800
rect 27066 200 27122 800
rect 28998 200 29054 800
rect 30286 200 30342 800
rect 32218 200 32274 800
rect 34150 200 34206 800
rect 35438 200 35494 800
rect 37370 200 37426 800
rect 39302 200 39358 800
<< via2 >>
rect 2962 39480 3018 39536
rect 2870 37440 2926 37496
rect 1674 36080 1730 36136
rect 1674 34040 1730 34096
rect 1582 32020 1638 32056
rect 1582 32000 1584 32020
rect 1584 32000 1636 32020
rect 1636 32000 1638 32020
rect 1674 30660 1730 30696
rect 1674 30640 1676 30660
rect 1676 30640 1728 30660
rect 1728 30640 1730 30660
rect 1582 28636 1584 28656
rect 1584 28636 1636 28656
rect 1636 28636 1638 28656
rect 1582 28600 1638 28636
rect 1674 26560 1730 26616
rect 1582 25236 1584 25256
rect 1584 25236 1636 25256
rect 1636 25236 1638 25256
rect 1582 25200 1638 25236
rect 1674 23160 1730 23216
rect 1674 21120 1730 21176
rect 1674 19760 1730 19816
rect 1582 17756 1584 17776
rect 1584 17756 1636 17776
rect 1636 17756 1638 17776
rect 1582 17720 1638 17756
rect 1674 15680 1730 15736
rect 1674 14320 1730 14376
rect 1674 12280 1730 12336
rect 1582 10260 1638 10296
rect 1582 10240 1584 10260
rect 1584 10240 1636 10260
rect 1636 10240 1638 10260
rect 1582 8916 1584 8936
rect 1584 8916 1636 8936
rect 1636 8916 1638 8936
rect 1582 8880 1638 8916
rect 1582 6840 1638 6896
rect 1674 4800 1730 4856
rect 1582 3476 1584 3496
rect 1584 3476 1636 3496
rect 1636 3476 1638 3496
rect 1582 3440 1638 3476
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4618 2896 4674 2952
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 1674 1400 1730 1456
rect 9586 12280 9642 12336
rect 9770 12144 9826 12200
rect 9862 11192 9918 11248
rect 9310 9152 9366 9208
rect 10782 15000 10838 15056
rect 11150 15444 11152 15464
rect 11152 15444 11204 15464
rect 11204 15444 11206 15464
rect 11150 15408 11206 15444
rect 10138 10920 10194 10976
rect 10322 13776 10378 13832
rect 10506 14356 10508 14376
rect 10508 14356 10560 14376
rect 10560 14356 10562 14376
rect 10506 14320 10562 14356
rect 10690 12688 10746 12744
rect 10782 12436 10838 12472
rect 10782 12416 10784 12436
rect 10784 12416 10836 12436
rect 10836 12416 10838 12436
rect 10506 9968 10562 10024
rect 10046 4276 10102 4312
rect 10046 4256 10048 4276
rect 10048 4256 10100 4276
rect 10100 4256 10102 4276
rect 11058 13388 11114 13424
rect 11058 13368 11060 13388
rect 11060 13368 11112 13388
rect 11112 13368 11114 13388
rect 11242 12824 11298 12880
rect 12070 16088 12126 16144
rect 12530 15816 12586 15872
rect 11978 14456 12034 14512
rect 11426 12280 11482 12336
rect 10874 9016 10930 9072
rect 10690 6024 10746 6080
rect 11610 11056 11666 11112
rect 11242 10104 11298 10160
rect 11242 9868 11244 9888
rect 11244 9868 11296 9888
rect 11296 9868 11298 9888
rect 11242 9832 11298 9868
rect 11242 8508 11244 8528
rect 11244 8508 11296 8528
rect 11296 8508 11298 8528
rect 11242 8472 11298 8508
rect 11150 6976 11206 7032
rect 10874 2796 10876 2816
rect 10876 2796 10928 2816
rect 10928 2796 10930 2816
rect 10874 2760 10930 2796
rect 11518 10512 11574 10568
rect 12438 14068 12494 14104
rect 12438 14048 12440 14068
rect 12440 14048 12492 14068
rect 12492 14048 12494 14068
rect 12346 13796 12402 13832
rect 12346 13776 12348 13796
rect 12348 13776 12400 13796
rect 12400 13776 12402 13796
rect 12346 13096 12402 13152
rect 12530 13676 12532 13696
rect 12532 13676 12584 13696
rect 12584 13676 12586 13696
rect 12530 13640 12586 13676
rect 12622 12960 12678 13016
rect 12346 11056 12402 11112
rect 11886 6196 11888 6216
rect 11888 6196 11940 6216
rect 11940 6196 11942 6216
rect 11886 6160 11942 6196
rect 11978 3712 12034 3768
rect 11886 3032 11942 3088
rect 12806 12688 12862 12744
rect 12346 5752 12402 5808
rect 12254 5480 12310 5536
rect 12254 4392 12310 4448
rect 13174 14340 13230 14376
rect 13174 14320 13176 14340
rect 13176 14320 13228 14340
rect 13228 14320 13230 14340
rect 14922 17040 14978 17096
rect 14922 15272 14978 15328
rect 14002 14456 14058 14512
rect 14462 14456 14518 14512
rect 13174 12688 13230 12744
rect 13266 10920 13322 10976
rect 13266 10548 13268 10568
rect 13268 10548 13320 10568
rect 13320 10548 13322 10568
rect 13266 10512 13322 10548
rect 13818 14048 13874 14104
rect 13910 13948 13912 13968
rect 13912 13948 13964 13968
rect 13964 13948 13966 13968
rect 13910 13912 13966 13948
rect 13910 13796 13966 13832
rect 13910 13776 13912 13796
rect 13912 13776 13964 13796
rect 13964 13776 13966 13796
rect 13726 12552 13782 12608
rect 13450 11076 13506 11112
rect 13450 11056 13452 11076
rect 13452 11056 13504 11076
rect 13504 11056 13506 11076
rect 14186 13096 14242 13152
rect 14094 12960 14150 13016
rect 13634 10104 13690 10160
rect 12622 5480 12678 5536
rect 12346 4120 12402 4176
rect 12438 3984 12494 4040
rect 12622 3732 12678 3768
rect 12622 3712 12624 3732
rect 12624 3712 12676 3732
rect 12676 3712 12678 3732
rect 13358 4392 13414 4448
rect 12806 2760 12862 2816
rect 12346 2388 12348 2408
rect 12348 2388 12400 2408
rect 12400 2388 12402 2408
rect 12346 2352 12402 2388
rect 14094 7928 14150 7984
rect 14646 13676 14648 13696
rect 14648 13676 14700 13696
rect 14700 13676 14702 13696
rect 14462 13404 14464 13424
rect 14464 13404 14516 13424
rect 14516 13404 14518 13424
rect 14462 13368 14518 13404
rect 14646 13640 14702 13676
rect 15014 13368 15070 13424
rect 15106 12688 15162 12744
rect 15014 12552 15070 12608
rect 15198 9968 15254 10024
rect 14922 9832 14978 9888
rect 13726 5072 13782 5128
rect 13634 4564 13636 4584
rect 13636 4564 13688 4584
rect 13688 4564 13690 4584
rect 13634 4528 13690 4564
rect 13910 3068 13912 3088
rect 13912 3068 13964 3088
rect 13964 3068 13966 3088
rect 13910 3032 13966 3068
rect 15750 15852 15752 15872
rect 15752 15852 15804 15872
rect 15804 15852 15806 15872
rect 15750 15816 15806 15852
rect 15566 12164 15622 12200
rect 15566 12144 15568 12164
rect 15568 12144 15620 12164
rect 15620 12144 15622 12164
rect 15014 7112 15070 7168
rect 15106 6432 15162 6488
rect 14554 4936 14610 4992
rect 14646 4428 14648 4448
rect 14648 4428 14700 4448
rect 14700 4428 14702 4448
rect 14646 4392 14702 4428
rect 14554 4120 14610 4176
rect 14646 3984 14702 4040
rect 14922 4256 14978 4312
rect 13726 2488 13782 2544
rect 16026 12416 16082 12472
rect 16302 15000 16358 15056
rect 16394 13640 16450 13696
rect 16118 6160 16174 6216
rect 16578 11056 16634 11112
rect 16486 9988 16542 10024
rect 16486 9968 16488 9988
rect 16488 9968 16540 9988
rect 16540 9968 16542 9988
rect 16394 9036 16450 9072
rect 16394 9016 16396 9036
rect 16396 9016 16448 9036
rect 16448 9016 16450 9036
rect 16486 6568 16542 6624
rect 16670 6024 16726 6080
rect 16486 5244 16488 5264
rect 16488 5244 16540 5264
rect 16540 5244 16542 5264
rect 16486 5208 16542 5244
rect 16854 4256 16910 4312
rect 17590 14900 17592 14920
rect 17592 14900 17644 14920
rect 17644 14900 17646 14920
rect 17590 14864 17646 14900
rect 17314 11192 17370 11248
rect 17590 12280 17646 12336
rect 17406 9696 17462 9752
rect 17314 8492 17370 8528
rect 17314 8472 17316 8492
rect 17316 8472 17368 8492
rect 17368 8472 17370 8492
rect 17314 3848 17370 3904
rect 17314 3440 17370 3496
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 18142 15308 18144 15328
rect 18144 15308 18196 15328
rect 18196 15308 18198 15328
rect 18142 15272 18198 15308
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19890 18808 19946 18864
rect 17866 13912 17922 13968
rect 17866 11056 17922 11112
rect 18326 12860 18328 12880
rect 18328 12860 18380 12880
rect 18380 12860 18382 12880
rect 18326 12824 18382 12860
rect 18050 7792 18106 7848
rect 18326 10104 18382 10160
rect 18510 7384 18566 7440
rect 17682 6976 17738 7032
rect 17958 6860 18014 6896
rect 17958 6840 17960 6860
rect 17960 6840 18012 6860
rect 18012 6840 18014 6860
rect 17590 6604 17592 6624
rect 17592 6604 17644 6624
rect 17644 6604 17646 6624
rect 17590 6568 17646 6604
rect 18970 14864 19026 14920
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19890 17740 19946 17776
rect 19890 17720 19892 17740
rect 19892 17720 19944 17740
rect 19944 17720 19946 17740
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19890 15680 19946 15736
rect 19522 15580 19524 15600
rect 19524 15580 19576 15600
rect 19576 15580 19578 15600
rect 19522 15544 19578 15580
rect 20074 15428 20130 15464
rect 20074 15408 20076 15428
rect 20076 15408 20128 15428
rect 20128 15408 20130 15428
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19154 13812 19156 13832
rect 19156 13812 19208 13832
rect 19208 13812 19210 13832
rect 19154 13776 19210 13812
rect 19798 14728 19854 14784
rect 19246 13368 19302 13424
rect 19246 13232 19302 13288
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19614 13504 19670 13560
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 18786 8900 18842 8936
rect 18786 8880 18788 8900
rect 18788 8880 18840 8900
rect 18840 8880 18842 8900
rect 18050 4936 18106 4992
rect 19430 12180 19432 12200
rect 19432 12180 19484 12200
rect 19484 12180 19486 12200
rect 19430 12144 19486 12180
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19430 11228 19432 11248
rect 19432 11228 19484 11248
rect 19484 11228 19486 11248
rect 19430 11192 19486 11228
rect 20626 17740 20682 17776
rect 20626 17720 20628 17740
rect 20628 17720 20680 17740
rect 20680 17720 20682 17740
rect 20534 15544 20590 15600
rect 20718 15272 20774 15328
rect 20534 14864 20590 14920
rect 20626 13368 20682 13424
rect 20258 11328 20314 11384
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19522 10668 19578 10704
rect 19522 10648 19524 10668
rect 19524 10648 19576 10668
rect 19576 10648 19578 10668
rect 19338 10240 19394 10296
rect 19706 10240 19762 10296
rect 19246 9832 19302 9888
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19430 9696 19486 9752
rect 20166 9696 20222 9752
rect 19614 9016 19670 9072
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19430 8472 19486 8528
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19614 6976 19670 7032
rect 19430 6840 19486 6896
rect 20074 7248 20130 7304
rect 20350 9832 20406 9888
rect 20258 8744 20314 8800
rect 19154 6316 19210 6352
rect 19154 6296 19156 6316
rect 19156 6296 19208 6316
rect 19208 6296 19210 6316
rect 19338 6432 19394 6488
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 18970 4020 18972 4040
rect 18972 4020 19024 4040
rect 19024 4020 19026 4040
rect 18970 3984 19026 4020
rect 19154 3848 19210 3904
rect 20258 5908 20314 5944
rect 20258 5888 20260 5908
rect 20260 5888 20312 5908
rect 20312 5888 20314 5908
rect 20626 12960 20682 13016
rect 20810 13932 20866 13968
rect 20810 13912 20812 13932
rect 20812 13912 20864 13932
rect 20864 13912 20866 13932
rect 21270 15020 21326 15056
rect 21270 15000 21272 15020
rect 21272 15000 21324 15020
rect 21324 15000 21326 15020
rect 20718 12316 20720 12336
rect 20720 12316 20772 12336
rect 20772 12316 20774 12336
rect 20718 12280 20774 12316
rect 20902 11328 20958 11384
rect 20442 7112 20498 7168
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 20074 4800 20130 4856
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 20718 8200 20774 8256
rect 20534 4664 20590 4720
rect 21178 8492 21234 8528
rect 21178 8472 21180 8492
rect 21180 8472 21232 8492
rect 21232 8472 21234 8492
rect 21270 7520 21326 7576
rect 21270 5480 21326 5536
rect 21546 11872 21602 11928
rect 22006 16108 22062 16144
rect 22006 16088 22008 16108
rect 22008 16088 22060 16108
rect 22060 16088 22062 16108
rect 21914 15544 21970 15600
rect 21730 13640 21786 13696
rect 21730 13524 21786 13560
rect 21730 13504 21732 13524
rect 21732 13504 21784 13524
rect 21784 13504 21786 13524
rect 22374 13640 22430 13696
rect 22282 12724 22284 12744
rect 22284 12724 22336 12744
rect 22336 12724 22338 12744
rect 22282 12688 22338 12724
rect 21638 9696 21694 9752
rect 21730 9288 21786 9344
rect 21546 7656 21602 7712
rect 21822 8084 21878 8120
rect 21822 8064 21824 8084
rect 21824 8064 21876 8084
rect 21876 8064 21878 8084
rect 22190 9596 22192 9616
rect 22192 9596 22244 9616
rect 22244 9596 22246 9616
rect 22834 14320 22890 14376
rect 23202 15408 23258 15464
rect 22190 9560 22246 9596
rect 22190 9424 22246 9480
rect 22282 8780 22284 8800
rect 22284 8780 22336 8800
rect 22336 8780 22338 8800
rect 22282 8744 22338 8780
rect 22650 9560 22706 9616
rect 23018 13388 23074 13424
rect 23018 13368 23020 13388
rect 23020 13368 23072 13388
rect 23072 13368 23074 13388
rect 22926 13096 22982 13152
rect 23110 12824 23166 12880
rect 22282 8064 22338 8120
rect 22558 8336 22614 8392
rect 22190 7692 22192 7712
rect 22192 7692 22244 7712
rect 22244 7692 22246 7712
rect 22190 7656 22246 7692
rect 22374 7112 22430 7168
rect 22098 6840 22154 6896
rect 22282 6840 22338 6896
rect 22190 5616 22246 5672
rect 22282 5344 22338 5400
rect 22558 6024 22614 6080
rect 22834 7112 22890 7168
rect 21178 3168 21234 3224
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 22006 2644 22062 2680
rect 22006 2624 22008 2644
rect 22008 2624 22060 2644
rect 22060 2624 22062 2644
rect 23386 15272 23442 15328
rect 23386 14048 23442 14104
rect 23754 15272 23810 15328
rect 23294 12144 23350 12200
rect 23478 12164 23534 12200
rect 23478 12144 23480 12164
rect 23480 12144 23532 12164
rect 23532 12144 23534 12164
rect 23202 11756 23258 11792
rect 23202 11736 23204 11756
rect 23204 11736 23256 11756
rect 23256 11736 23258 11756
rect 23570 11192 23626 11248
rect 23294 9444 23350 9480
rect 23294 9424 23296 9444
rect 23296 9424 23348 9444
rect 23348 9424 23350 9444
rect 23202 4664 23258 4720
rect 22926 4120 22982 4176
rect 23386 7656 23442 7712
rect 24398 17584 24454 17640
rect 24214 15272 24270 15328
rect 24306 13776 24362 13832
rect 24030 11600 24086 11656
rect 23478 4020 23480 4040
rect 23480 4020 23532 4040
rect 23532 4020 23534 4040
rect 23478 3984 23534 4020
rect 22466 3304 22522 3360
rect 23386 3032 23442 3088
rect 25042 14864 25098 14920
rect 24398 10240 24454 10296
rect 24950 11056 25006 11112
rect 25134 10548 25136 10568
rect 25136 10548 25188 10568
rect 25188 10548 25190 10568
rect 25134 10512 25190 10548
rect 23938 3576 23994 3632
rect 23938 2896 23994 2952
rect 25962 17620 25964 17640
rect 25964 17620 26016 17640
rect 26016 17620 26018 17640
rect 25962 17584 26018 17620
rect 26422 15680 26478 15736
rect 26514 15272 26570 15328
rect 26514 14764 26516 14784
rect 26516 14764 26568 14784
rect 26568 14764 26570 14784
rect 26514 14728 26570 14764
rect 25962 13504 26018 13560
rect 25870 12980 25926 13016
rect 25870 12960 25872 12980
rect 25872 12960 25924 12980
rect 25924 12960 25926 12980
rect 27066 13640 27122 13696
rect 25686 12688 25742 12744
rect 27250 13096 27306 13152
rect 26974 12824 27030 12880
rect 27526 15020 27582 15056
rect 27526 15000 27528 15020
rect 27528 15000 27580 15020
rect 27580 15000 27582 15020
rect 27526 14356 27528 14376
rect 27528 14356 27580 14376
rect 27580 14356 27582 14376
rect 27526 14320 27582 14356
rect 27710 14048 27766 14104
rect 27526 12688 27582 12744
rect 27986 16224 28042 16280
rect 26054 11872 26110 11928
rect 26330 11772 26332 11792
rect 26332 11772 26384 11792
rect 26384 11772 26386 11792
rect 26330 11736 26386 11772
rect 25778 10240 25834 10296
rect 26146 11076 26202 11112
rect 26146 11056 26148 11076
rect 26148 11056 26200 11076
rect 26200 11056 26202 11076
rect 26054 10648 26110 10704
rect 25686 7792 25742 7848
rect 25410 6840 25466 6896
rect 26514 10512 26570 10568
rect 26330 9152 26386 9208
rect 26330 7928 26386 7984
rect 25962 7112 26018 7168
rect 25778 6976 25834 7032
rect 26514 6432 26570 6488
rect 26514 5616 26570 5672
rect 26422 4020 26424 4040
rect 26424 4020 26476 4040
rect 26476 4020 26478 4040
rect 26422 3984 26478 4020
rect 27710 12144 27766 12200
rect 27618 11192 27674 11248
rect 27526 9832 27582 9888
rect 27526 9596 27528 9616
rect 27528 9596 27580 9616
rect 27580 9596 27582 9616
rect 27526 9560 27582 9596
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 37186 38800 37242 38856
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 38290 37440 38346 37496
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 28446 11600 28502 11656
rect 27434 7692 27436 7712
rect 27436 7692 27488 7712
rect 27488 7692 27490 7712
rect 27434 7656 27490 7692
rect 26698 5888 26754 5944
rect 27066 5752 27122 5808
rect 27158 5480 27214 5536
rect 27250 5364 27306 5400
rect 27894 7520 27950 7576
rect 27802 6432 27858 6488
rect 27250 5344 27252 5364
rect 27252 5344 27304 5364
rect 27304 5344 27306 5364
rect 26514 2624 26570 2680
rect 27526 5072 27582 5128
rect 27066 3032 27122 3088
rect 28538 9152 28594 9208
rect 28722 9288 28778 9344
rect 28722 8372 28724 8392
rect 28724 8372 28776 8392
rect 28776 8372 28778 8392
rect 28722 8336 28778 8372
rect 29274 10104 29330 10160
rect 29182 9968 29238 10024
rect 28998 8200 29054 8256
rect 29182 7420 29184 7440
rect 29184 7420 29236 7440
rect 29236 7420 29238 7440
rect 29182 7384 29238 7420
rect 29366 9460 29368 9480
rect 29368 9460 29420 9480
rect 29420 9460 29422 9480
rect 29366 9424 29422 9460
rect 28630 6024 28686 6080
rect 28354 3440 28410 3496
rect 28722 4528 28778 4584
rect 28630 3304 28686 3360
rect 28538 3168 28594 3224
rect 28630 2932 28632 2952
rect 28632 2932 28684 2952
rect 28684 2932 28686 2952
rect 28630 2896 28686 2932
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 30286 8880 30342 8936
rect 30470 7268 30526 7304
rect 30470 7248 30472 7268
rect 30472 7248 30524 7268
rect 30524 7248 30526 7268
rect 29826 2508 29882 2544
rect 29826 2488 29828 2508
rect 29828 2488 29880 2508
rect 29880 2488 29882 2508
rect 29918 2352 29974 2408
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 38290 35400 38346 35456
rect 38198 33380 38254 33416
rect 38198 33360 38200 33380
rect 38200 33360 38252 33380
rect 38252 33360 38254 33380
rect 38290 32020 38346 32056
rect 38290 32000 38292 32020
rect 38292 32000 38344 32020
rect 38344 32000 38346 32020
rect 38198 29996 38200 30016
rect 38200 29996 38252 30016
rect 38252 29996 38254 30016
rect 38198 29960 38254 29996
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 31022 6296 31078 6352
rect 31114 5208 31170 5264
rect 32954 3596 33010 3632
rect 32954 3576 32956 3596
rect 32956 3576 33008 3596
rect 33008 3576 33010 3596
rect 31022 2932 31024 2952
rect 31024 2932 31076 2952
rect 31076 2932 31078 2952
rect 31022 2896 31078 2932
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 38198 27940 38254 27976
rect 38198 27920 38200 27940
rect 38200 27920 38252 27940
rect 38252 27920 38254 27940
rect 38290 26580 38346 26616
rect 38290 26560 38292 26580
rect 38292 26560 38344 26580
rect 38344 26560 38346 26580
rect 38198 24556 38200 24576
rect 38200 24556 38252 24576
rect 38252 24556 38254 24576
rect 38198 24520 38254 24556
rect 38198 22480 38254 22536
rect 38198 21120 38254 21176
rect 38198 19116 38200 19136
rect 38200 19116 38252 19136
rect 38252 19116 38254 19136
rect 38198 19080 38254 19116
rect 38198 17040 38254 17096
rect 38014 15972 38070 16008
rect 38014 15952 38016 15972
rect 38016 15952 38068 15972
rect 38068 15952 38070 15972
rect 38198 15680 38254 15736
rect 38198 13640 38254 13696
rect 38198 11600 38254 11656
rect 38198 10240 38254 10296
rect 38198 8200 38254 8256
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 37922 6704 37978 6760
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 38198 6160 38254 6216
rect 38290 4820 38346 4856
rect 38290 4800 38292 4820
rect 38292 4800 38344 4820
rect 38344 4800 38346 4820
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 38198 2796 38200 2816
rect 38200 2796 38252 2816
rect 38252 2796 38254 2816
rect 38198 2760 38254 2796
rect 37186 1400 37242 1456
<< metal3 >>
rect 200 39538 800 39568
rect 2957 39538 3023 39541
rect 200 39536 3023 39538
rect 200 39480 2962 39536
rect 3018 39480 3023 39536
rect 200 39478 3023 39480
rect 200 39448 800 39478
rect 2957 39475 3023 39478
rect 37181 38858 37247 38861
rect 39200 38858 39800 38888
rect 37181 38856 39800 38858
rect 37181 38800 37186 38856
rect 37242 38800 39800 38856
rect 37181 38798 39800 38800
rect 37181 38795 37247 38798
rect 39200 38768 39800 38798
rect 4210 37568 4526 37569
rect 200 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 2865 37498 2931 37501
rect 200 37496 2931 37498
rect 200 37440 2870 37496
rect 2926 37440 2931 37496
rect 200 37438 2931 37440
rect 200 37408 800 37438
rect 2865 37435 2931 37438
rect 38285 37498 38351 37501
rect 39200 37498 39800 37528
rect 38285 37496 39800 37498
rect 38285 37440 38290 37496
rect 38346 37440 39800 37496
rect 38285 37438 39800 37440
rect 38285 37435 38351 37438
rect 39200 37408 39800 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 200 36138 800 36168
rect 1669 36138 1735 36141
rect 200 36136 1735 36138
rect 200 36080 1674 36136
rect 1730 36080 1735 36136
rect 200 36078 1735 36080
rect 200 36048 800 36078
rect 1669 36075 1735 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 38285 35458 38351 35461
rect 39200 35458 39800 35488
rect 38285 35456 39800 35458
rect 38285 35400 38290 35456
rect 38346 35400 39800 35456
rect 38285 35398 39800 35400
rect 38285 35395 38351 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 39200 35368 39800 35398
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 200 34098 800 34128
rect 1669 34098 1735 34101
rect 200 34096 1735 34098
rect 200 34040 1674 34096
rect 1730 34040 1735 34096
rect 200 34038 1735 34040
rect 200 34008 800 34038
rect 1669 34035 1735 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 38193 33418 38259 33421
rect 39200 33418 39800 33448
rect 38193 33416 39800 33418
rect 38193 33360 38198 33416
rect 38254 33360 39800 33416
rect 38193 33358 39800 33360
rect 38193 33355 38259 33358
rect 39200 33328 39800 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 200 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1577 32058 1643 32061
rect 200 32056 1643 32058
rect 200 32000 1582 32056
rect 1638 32000 1643 32056
rect 200 31998 1643 32000
rect 200 31968 800 31998
rect 1577 31995 1643 31998
rect 38285 32058 38351 32061
rect 39200 32058 39800 32088
rect 38285 32056 39800 32058
rect 38285 32000 38290 32056
rect 38346 32000 39800 32056
rect 38285 31998 39800 32000
rect 38285 31995 38351 31998
rect 39200 31968 39800 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30698 800 30728
rect 1669 30698 1735 30701
rect 200 30696 1735 30698
rect 200 30640 1674 30696
rect 1730 30640 1735 30696
rect 200 30638 1735 30640
rect 200 30608 800 30638
rect 1669 30635 1735 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 38193 30018 38259 30021
rect 39200 30018 39800 30048
rect 38193 30016 39800 30018
rect 38193 29960 38198 30016
rect 38254 29960 39800 30016
rect 38193 29958 39800 29960
rect 38193 29955 38259 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 39200 29928 39800 29958
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 200 28658 800 28688
rect 1577 28658 1643 28661
rect 200 28656 1643 28658
rect 200 28600 1582 28656
rect 1638 28600 1643 28656
rect 200 28598 1643 28600
rect 200 28568 800 28598
rect 1577 28595 1643 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 38193 27978 38259 27981
rect 39200 27978 39800 28008
rect 38193 27976 39800 27978
rect 38193 27920 38198 27976
rect 38254 27920 39800 27976
rect 38193 27918 39800 27920
rect 38193 27915 38259 27918
rect 39200 27888 39800 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 200 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 1669 26618 1735 26621
rect 200 26616 1735 26618
rect 200 26560 1674 26616
rect 1730 26560 1735 26616
rect 200 26558 1735 26560
rect 200 26528 800 26558
rect 1669 26555 1735 26558
rect 38285 26618 38351 26621
rect 39200 26618 39800 26648
rect 38285 26616 39800 26618
rect 38285 26560 38290 26616
rect 38346 26560 39800 26616
rect 38285 26558 39800 26560
rect 38285 26555 38351 26558
rect 39200 26528 39800 26558
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 200 25258 800 25288
rect 1577 25258 1643 25261
rect 200 25256 1643 25258
rect 200 25200 1582 25256
rect 1638 25200 1643 25256
rect 200 25198 1643 25200
rect 200 25168 800 25198
rect 1577 25195 1643 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 38193 24578 38259 24581
rect 39200 24578 39800 24608
rect 38193 24576 39800 24578
rect 38193 24520 38198 24576
rect 38254 24520 39800 24576
rect 38193 24518 39800 24520
rect 38193 24515 38259 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 39200 24488 39800 24518
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 200 23218 800 23248
rect 1669 23218 1735 23221
rect 200 23216 1735 23218
rect 200 23160 1674 23216
rect 1730 23160 1735 23216
rect 200 23158 1735 23160
rect 200 23128 800 23158
rect 1669 23155 1735 23158
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 38193 22538 38259 22541
rect 39200 22538 39800 22568
rect 38193 22536 39800 22538
rect 38193 22480 38198 22536
rect 38254 22480 39800 22536
rect 38193 22478 39800 22480
rect 38193 22475 38259 22478
rect 39200 22448 39800 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 200 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 1669 21178 1735 21181
rect 200 21176 1735 21178
rect 200 21120 1674 21176
rect 1730 21120 1735 21176
rect 200 21118 1735 21120
rect 200 21088 800 21118
rect 1669 21115 1735 21118
rect 38193 21178 38259 21181
rect 39200 21178 39800 21208
rect 38193 21176 39800 21178
rect 38193 21120 38198 21176
rect 38254 21120 39800 21176
rect 38193 21118 39800 21120
rect 38193 21115 38259 21118
rect 39200 21088 39800 21118
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 200 19818 800 19848
rect 1669 19818 1735 19821
rect 200 19816 1735 19818
rect 200 19760 1674 19816
rect 1730 19760 1735 19816
rect 200 19758 1735 19760
rect 200 19728 800 19758
rect 1669 19755 1735 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 38193 19138 38259 19141
rect 39200 19138 39800 19168
rect 38193 19136 39800 19138
rect 38193 19080 38198 19136
rect 38254 19080 39800 19136
rect 38193 19078 39800 19080
rect 38193 19075 38259 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 39800 19078
rect 34930 19007 35246 19008
rect 19885 18866 19951 18869
rect 20110 18866 20116 18868
rect 19885 18864 20116 18866
rect 19885 18808 19890 18864
rect 19946 18808 20116 18864
rect 19885 18806 20116 18808
rect 19885 18803 19951 18806
rect 20110 18804 20116 18806
rect 20180 18804 20186 18868
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 200 17778 800 17808
rect 1577 17778 1643 17781
rect 200 17776 1643 17778
rect 200 17720 1582 17776
rect 1638 17720 1643 17776
rect 200 17718 1643 17720
rect 200 17688 800 17718
rect 1577 17715 1643 17718
rect 19885 17778 19951 17781
rect 20621 17778 20687 17781
rect 19885 17776 20687 17778
rect 19885 17720 19890 17776
rect 19946 17720 20626 17776
rect 20682 17720 20687 17776
rect 19885 17718 20687 17720
rect 19885 17715 19951 17718
rect 20621 17715 20687 17718
rect 24393 17642 24459 17645
rect 25957 17642 26023 17645
rect 24393 17640 26023 17642
rect 24393 17584 24398 17640
rect 24454 17584 25962 17640
rect 26018 17584 26023 17640
rect 24393 17582 26023 17584
rect 24393 17579 24459 17582
rect 25957 17579 26023 17582
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 14590 17036 14596 17100
rect 14660 17098 14666 17100
rect 14917 17098 14983 17101
rect 14660 17096 14983 17098
rect 14660 17040 14922 17096
rect 14978 17040 14983 17096
rect 14660 17038 14983 17040
rect 14660 17036 14666 17038
rect 14917 17035 14983 17038
rect 38193 17098 38259 17101
rect 39200 17098 39800 17128
rect 38193 17096 39800 17098
rect 38193 17040 38198 17096
rect 38254 17040 39800 17096
rect 38193 17038 39800 17040
rect 38193 17035 38259 17038
rect 39200 17008 39800 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 20110 16220 20116 16284
rect 20180 16282 20186 16284
rect 27981 16282 28047 16285
rect 20180 16280 28047 16282
rect 20180 16224 27986 16280
rect 28042 16224 28047 16280
rect 20180 16222 28047 16224
rect 20180 16220 20186 16222
rect 27981 16219 28047 16222
rect 12065 16146 12131 16149
rect 22001 16146 22067 16149
rect 12065 16144 22067 16146
rect 12065 16088 12070 16144
rect 12126 16088 22006 16144
rect 22062 16088 22067 16144
rect 12065 16086 22067 16088
rect 12065 16083 12131 16086
rect 22001 16083 22067 16086
rect 20662 15948 20668 16012
rect 20732 16010 20738 16012
rect 38009 16010 38075 16013
rect 20732 16008 38075 16010
rect 20732 15952 38014 16008
rect 38070 15952 38075 16008
rect 20732 15950 38075 15952
rect 20732 15948 20738 15950
rect 38009 15947 38075 15950
rect 12525 15874 12591 15877
rect 15745 15874 15811 15877
rect 12525 15872 15811 15874
rect 12525 15816 12530 15872
rect 12586 15816 15750 15872
rect 15806 15816 15811 15872
rect 12525 15814 15811 15816
rect 12525 15811 12591 15814
rect 15745 15811 15811 15814
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1669 15738 1735 15741
rect 200 15736 1735 15738
rect 200 15680 1674 15736
rect 1730 15680 1735 15736
rect 200 15678 1735 15680
rect 200 15648 800 15678
rect 1669 15675 1735 15678
rect 19885 15738 19951 15741
rect 26417 15738 26483 15741
rect 19885 15736 26483 15738
rect 19885 15680 19890 15736
rect 19946 15680 26422 15736
rect 26478 15680 26483 15736
rect 19885 15678 26483 15680
rect 19885 15675 19951 15678
rect 26417 15675 26483 15678
rect 38193 15738 38259 15741
rect 39200 15738 39800 15768
rect 38193 15736 39800 15738
rect 38193 15680 38198 15736
rect 38254 15680 39800 15736
rect 38193 15678 39800 15680
rect 38193 15675 38259 15678
rect 39200 15648 39800 15678
rect 19374 15540 19380 15604
rect 19444 15602 19450 15604
rect 19517 15602 19583 15605
rect 19444 15600 19583 15602
rect 19444 15544 19522 15600
rect 19578 15544 19583 15600
rect 19444 15542 19583 15544
rect 19444 15540 19450 15542
rect 19517 15539 19583 15542
rect 20529 15602 20595 15605
rect 21909 15602 21975 15605
rect 20529 15600 21975 15602
rect 20529 15544 20534 15600
rect 20590 15544 21914 15600
rect 21970 15544 21975 15600
rect 20529 15542 21975 15544
rect 20529 15539 20595 15542
rect 21909 15539 21975 15542
rect 11145 15466 11211 15469
rect 11278 15466 11284 15468
rect 11145 15464 11284 15466
rect 11145 15408 11150 15464
rect 11206 15408 11284 15464
rect 11145 15406 11284 15408
rect 11145 15403 11211 15406
rect 11278 15404 11284 15406
rect 11348 15404 11354 15468
rect 20069 15466 20135 15469
rect 23197 15466 23263 15469
rect 20069 15464 23263 15466
rect 20069 15408 20074 15464
rect 20130 15408 23202 15464
rect 23258 15408 23263 15464
rect 20069 15406 23263 15408
rect 20069 15403 20135 15406
rect 23197 15403 23263 15406
rect 14917 15330 14983 15333
rect 18137 15330 18203 15333
rect 14917 15328 18203 15330
rect 14917 15272 14922 15328
rect 14978 15272 18142 15328
rect 18198 15272 18203 15328
rect 14917 15270 18203 15272
rect 14917 15267 14983 15270
rect 18137 15267 18203 15270
rect 20713 15330 20779 15333
rect 23381 15330 23447 15333
rect 20713 15328 23447 15330
rect 20713 15272 20718 15328
rect 20774 15272 23386 15328
rect 23442 15272 23447 15328
rect 20713 15270 23447 15272
rect 20713 15267 20779 15270
rect 23381 15267 23447 15270
rect 23749 15330 23815 15333
rect 24209 15330 24275 15333
rect 26509 15330 26575 15333
rect 23749 15328 26575 15330
rect 23749 15272 23754 15328
rect 23810 15272 24214 15328
rect 24270 15272 26514 15328
rect 26570 15272 26575 15328
rect 23749 15270 26575 15272
rect 23749 15267 23815 15270
rect 24209 15267 24275 15270
rect 26509 15267 26575 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 10777 15058 10843 15061
rect 16297 15058 16363 15061
rect 10777 15056 16363 15058
rect 10777 15000 10782 15056
rect 10838 15000 16302 15056
rect 16358 15000 16363 15056
rect 10777 14998 16363 15000
rect 10777 14995 10843 14998
rect 16297 14995 16363 14998
rect 21265 15058 21331 15061
rect 27521 15058 27587 15061
rect 21265 15056 27587 15058
rect 21265 15000 21270 15056
rect 21326 15000 27526 15056
rect 27582 15000 27587 15056
rect 21265 14998 27587 15000
rect 21265 14995 21331 14998
rect 27521 14995 27587 14998
rect 17585 14922 17651 14925
rect 18965 14922 19031 14925
rect 17585 14920 19031 14922
rect 17585 14864 17590 14920
rect 17646 14864 18970 14920
rect 19026 14864 19031 14920
rect 17585 14862 19031 14864
rect 17585 14859 17651 14862
rect 18965 14859 19031 14862
rect 20529 14922 20595 14925
rect 25037 14922 25103 14925
rect 20529 14920 25103 14922
rect 20529 14864 20534 14920
rect 20590 14864 25042 14920
rect 25098 14864 25103 14920
rect 20529 14862 25103 14864
rect 20529 14859 20595 14862
rect 25037 14859 25103 14862
rect 19793 14786 19859 14789
rect 26509 14786 26575 14789
rect 19793 14784 26575 14786
rect 19793 14728 19798 14784
rect 19854 14728 26514 14784
rect 26570 14728 26575 14784
rect 19793 14726 26575 14728
rect 19793 14723 19859 14726
rect 26509 14723 26575 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 11973 14514 12039 14517
rect 13997 14514 14063 14517
rect 14457 14514 14523 14517
rect 11973 14512 14523 14514
rect 11973 14456 11978 14512
rect 12034 14456 14002 14512
rect 14058 14456 14462 14512
rect 14518 14456 14523 14512
rect 11973 14454 14523 14456
rect 11973 14451 12039 14454
rect 13997 14451 14063 14454
rect 14457 14451 14523 14454
rect 200 14378 800 14408
rect 1669 14378 1735 14381
rect 200 14376 1735 14378
rect 200 14320 1674 14376
rect 1730 14320 1735 14376
rect 200 14318 1735 14320
rect 200 14288 800 14318
rect 1669 14315 1735 14318
rect 10501 14378 10567 14381
rect 13169 14378 13235 14381
rect 10501 14376 13235 14378
rect 10501 14320 10506 14376
rect 10562 14320 13174 14376
rect 13230 14320 13235 14376
rect 10501 14318 13235 14320
rect 10501 14315 10567 14318
rect 13169 14315 13235 14318
rect 22829 14378 22895 14381
rect 27521 14378 27587 14381
rect 22829 14376 27587 14378
rect 22829 14320 22834 14376
rect 22890 14320 27526 14376
rect 27582 14320 27587 14376
rect 22829 14318 27587 14320
rect 22829 14315 22895 14318
rect 27521 14315 27587 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 12433 14106 12499 14109
rect 13813 14106 13879 14109
rect 12433 14104 13879 14106
rect 12433 14048 12438 14104
rect 12494 14048 13818 14104
rect 13874 14048 13879 14104
rect 12433 14046 13879 14048
rect 12433 14043 12499 14046
rect 13813 14043 13879 14046
rect 23381 14106 23447 14109
rect 27705 14106 27771 14109
rect 23381 14104 27771 14106
rect 23381 14048 23386 14104
rect 23442 14048 27710 14104
rect 27766 14048 27771 14104
rect 23381 14046 27771 14048
rect 23381 14043 23447 14046
rect 27705 14043 27771 14046
rect 13905 13970 13971 13973
rect 10366 13968 13971 13970
rect 10366 13912 13910 13968
rect 13966 13912 13971 13968
rect 10366 13910 13971 13912
rect 10366 13837 10426 13910
rect 13905 13907 13971 13910
rect 17861 13970 17927 13973
rect 20805 13970 20871 13973
rect 17861 13968 20871 13970
rect 17861 13912 17866 13968
rect 17922 13912 20810 13968
rect 20866 13912 20871 13968
rect 17861 13910 20871 13912
rect 17861 13907 17927 13910
rect 20805 13907 20871 13910
rect 10317 13832 10426 13837
rect 10317 13776 10322 13832
rect 10378 13776 10426 13832
rect 10317 13774 10426 13776
rect 12341 13834 12407 13837
rect 13905 13834 13971 13837
rect 12341 13832 13971 13834
rect 12341 13776 12346 13832
rect 12402 13776 13910 13832
rect 13966 13776 13971 13832
rect 12341 13774 13971 13776
rect 10317 13771 10383 13774
rect 12341 13771 12407 13774
rect 13905 13771 13971 13774
rect 19149 13834 19215 13837
rect 24301 13834 24367 13837
rect 19149 13832 24367 13834
rect 19149 13776 19154 13832
rect 19210 13776 24306 13832
rect 24362 13776 24367 13832
rect 19149 13774 24367 13776
rect 19149 13771 19215 13774
rect 24301 13771 24367 13774
rect 12525 13698 12591 13701
rect 14641 13698 14707 13701
rect 12525 13696 14707 13698
rect 12525 13640 12530 13696
rect 12586 13640 14646 13696
rect 14702 13640 14707 13696
rect 12525 13638 14707 13640
rect 12525 13635 12591 13638
rect 14641 13635 14707 13638
rect 16389 13698 16455 13701
rect 21725 13698 21791 13701
rect 16389 13696 21791 13698
rect 16389 13640 16394 13696
rect 16450 13640 21730 13696
rect 21786 13640 21791 13696
rect 16389 13638 21791 13640
rect 16389 13635 16455 13638
rect 21725 13635 21791 13638
rect 22369 13698 22435 13701
rect 27061 13698 27127 13701
rect 22369 13696 27127 13698
rect 22369 13640 22374 13696
rect 22430 13640 27066 13696
rect 27122 13640 27127 13696
rect 22369 13638 27127 13640
rect 22369 13635 22435 13638
rect 27061 13635 27127 13638
rect 38193 13698 38259 13701
rect 39200 13698 39800 13728
rect 38193 13696 39800 13698
rect 38193 13640 38198 13696
rect 38254 13640 39800 13696
rect 38193 13638 39800 13640
rect 38193 13635 38259 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 39200 13608 39800 13638
rect 34930 13567 35246 13568
rect 19374 13500 19380 13564
rect 19444 13562 19450 13564
rect 19609 13562 19675 13565
rect 19444 13560 19675 13562
rect 19444 13504 19614 13560
rect 19670 13504 19675 13560
rect 19444 13502 19675 13504
rect 19444 13500 19450 13502
rect 19609 13499 19675 13502
rect 21725 13562 21791 13565
rect 25957 13562 26023 13565
rect 21725 13560 26023 13562
rect 21725 13504 21730 13560
rect 21786 13504 25962 13560
rect 26018 13504 26023 13560
rect 21725 13502 26023 13504
rect 21725 13499 21791 13502
rect 25957 13499 26023 13502
rect 11053 13426 11119 13429
rect 14457 13426 14523 13429
rect 11053 13424 14523 13426
rect 11053 13368 11058 13424
rect 11114 13368 14462 13424
rect 14518 13368 14523 13424
rect 11053 13366 14523 13368
rect 11053 13363 11119 13366
rect 14457 13363 14523 13366
rect 15009 13426 15075 13429
rect 19241 13426 19307 13429
rect 15009 13424 19307 13426
rect 15009 13368 15014 13424
rect 15070 13368 19246 13424
rect 19302 13368 19307 13424
rect 15009 13366 19307 13368
rect 15009 13363 15075 13366
rect 19241 13363 19307 13366
rect 20621 13426 20687 13429
rect 23013 13426 23079 13429
rect 20621 13424 23079 13426
rect 20621 13368 20626 13424
rect 20682 13368 23018 13424
rect 23074 13368 23079 13424
rect 20621 13366 23079 13368
rect 20621 13363 20687 13366
rect 23013 13363 23079 13366
rect 19241 13290 19307 13293
rect 20110 13290 20116 13292
rect 19241 13288 20116 13290
rect 19241 13232 19246 13288
rect 19302 13232 20116 13288
rect 19241 13230 20116 13232
rect 19241 13227 19307 13230
rect 20110 13228 20116 13230
rect 20180 13228 20186 13292
rect 12341 13154 12407 13157
rect 14181 13154 14247 13157
rect 12341 13152 14247 13154
rect 12341 13096 12346 13152
rect 12402 13096 14186 13152
rect 14242 13096 14247 13152
rect 12341 13094 14247 13096
rect 12341 13091 12407 13094
rect 14181 13091 14247 13094
rect 22921 13154 22987 13157
rect 27245 13154 27311 13157
rect 22921 13152 27311 13154
rect 22921 13096 22926 13152
rect 22982 13096 27250 13152
rect 27306 13096 27311 13152
rect 22921 13094 27311 13096
rect 22921 13091 22987 13094
rect 27245 13091 27311 13094
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 12617 13018 12683 13021
rect 14089 13018 14155 13021
rect 12617 13016 14155 13018
rect 12617 12960 12622 13016
rect 12678 12960 14094 13016
rect 14150 12960 14155 13016
rect 12617 12958 14155 12960
rect 12617 12955 12683 12958
rect 14089 12955 14155 12958
rect 20621 13018 20687 13021
rect 25865 13018 25931 13021
rect 20621 13016 25931 13018
rect 20621 12960 20626 13016
rect 20682 12960 25870 13016
rect 25926 12960 25931 13016
rect 20621 12958 25931 12960
rect 20621 12955 20687 12958
rect 25865 12955 25931 12958
rect 11237 12882 11303 12885
rect 18321 12882 18387 12885
rect 11237 12880 18387 12882
rect 11237 12824 11242 12880
rect 11298 12824 18326 12880
rect 18382 12824 18387 12880
rect 11237 12822 18387 12824
rect 11237 12819 11303 12822
rect 18321 12819 18387 12822
rect 23105 12882 23171 12885
rect 26969 12882 27035 12885
rect 23105 12880 27035 12882
rect 23105 12824 23110 12880
rect 23166 12824 26974 12880
rect 27030 12824 27035 12880
rect 23105 12822 27035 12824
rect 23105 12819 23171 12822
rect 26969 12819 27035 12822
rect 10685 12746 10751 12749
rect 12801 12746 12867 12749
rect 10685 12744 12867 12746
rect 10685 12688 10690 12744
rect 10746 12688 12806 12744
rect 12862 12688 12867 12744
rect 10685 12686 12867 12688
rect 10685 12683 10751 12686
rect 12801 12683 12867 12686
rect 13169 12746 13235 12749
rect 15101 12746 15167 12749
rect 22277 12746 22343 12749
rect 13169 12744 22343 12746
rect 13169 12688 13174 12744
rect 13230 12688 15106 12744
rect 15162 12688 22282 12744
rect 22338 12688 22343 12744
rect 13169 12686 22343 12688
rect 13169 12683 13235 12686
rect 15101 12683 15167 12686
rect 22277 12683 22343 12686
rect 25681 12746 25747 12749
rect 27521 12746 27587 12749
rect 25681 12744 27587 12746
rect 25681 12688 25686 12744
rect 25742 12688 27526 12744
rect 27582 12688 27587 12744
rect 25681 12686 27587 12688
rect 25681 12683 25747 12686
rect 27521 12683 27587 12686
rect 13721 12610 13787 12613
rect 15009 12610 15075 12613
rect 13721 12608 15075 12610
rect 13721 12552 13726 12608
rect 13782 12552 15014 12608
rect 15070 12552 15075 12608
rect 13721 12550 15075 12552
rect 13721 12547 13787 12550
rect 15009 12547 15075 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 10777 12474 10843 12477
rect 16021 12474 16087 12477
rect 10777 12472 16087 12474
rect 10777 12416 10782 12472
rect 10838 12416 16026 12472
rect 16082 12416 16087 12472
rect 10777 12414 16087 12416
rect 10777 12411 10843 12414
rect 16021 12411 16087 12414
rect 200 12338 800 12368
rect 1669 12338 1735 12341
rect 200 12336 1735 12338
rect 200 12280 1674 12336
rect 1730 12280 1735 12336
rect 200 12278 1735 12280
rect 200 12248 800 12278
rect 1669 12275 1735 12278
rect 9581 12338 9647 12341
rect 11421 12338 11487 12341
rect 9581 12336 11487 12338
rect 9581 12280 9586 12336
rect 9642 12280 11426 12336
rect 11482 12280 11487 12336
rect 9581 12278 11487 12280
rect 9581 12275 9647 12278
rect 11421 12275 11487 12278
rect 17585 12338 17651 12341
rect 20713 12338 20779 12341
rect 17585 12336 20779 12338
rect 17585 12280 17590 12336
rect 17646 12280 20718 12336
rect 20774 12280 20779 12336
rect 17585 12278 20779 12280
rect 17585 12275 17651 12278
rect 20713 12275 20779 12278
rect 9765 12202 9831 12205
rect 15561 12202 15627 12205
rect 9765 12200 15627 12202
rect 9765 12144 9770 12200
rect 9826 12144 15566 12200
rect 15622 12144 15627 12200
rect 9765 12142 15627 12144
rect 9765 12139 9831 12142
rect 15561 12139 15627 12142
rect 19425 12202 19491 12205
rect 23289 12202 23355 12205
rect 19425 12200 23355 12202
rect 19425 12144 19430 12200
rect 19486 12144 23294 12200
rect 23350 12144 23355 12200
rect 19425 12142 23355 12144
rect 19425 12139 19491 12142
rect 23289 12139 23355 12142
rect 23473 12202 23539 12205
rect 27705 12202 27771 12205
rect 23473 12200 27771 12202
rect 23473 12144 23478 12200
rect 23534 12144 27710 12200
rect 27766 12144 27771 12200
rect 23473 12142 27771 12144
rect 23473 12139 23539 12142
rect 27705 12139 27771 12142
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 21541 11930 21607 11933
rect 26049 11930 26115 11933
rect 21541 11928 26115 11930
rect 21541 11872 21546 11928
rect 21602 11872 26054 11928
rect 26110 11872 26115 11928
rect 21541 11870 26115 11872
rect 21541 11867 21607 11870
rect 26049 11867 26115 11870
rect 23197 11794 23263 11797
rect 26325 11794 26391 11797
rect 23197 11792 26391 11794
rect 23197 11736 23202 11792
rect 23258 11736 26330 11792
rect 26386 11736 26391 11792
rect 23197 11734 26391 11736
rect 23197 11731 23263 11734
rect 26325 11731 26391 11734
rect 24025 11658 24091 11661
rect 28441 11658 28507 11661
rect 24025 11656 28507 11658
rect 24025 11600 24030 11656
rect 24086 11600 28446 11656
rect 28502 11600 28507 11656
rect 24025 11598 28507 11600
rect 24025 11595 24091 11598
rect 28441 11595 28507 11598
rect 38193 11658 38259 11661
rect 39200 11658 39800 11688
rect 38193 11656 39800 11658
rect 38193 11600 38198 11656
rect 38254 11600 39800 11656
rect 38193 11598 39800 11600
rect 38193 11595 38259 11598
rect 39200 11568 39800 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 20253 11386 20319 11389
rect 20897 11386 20963 11389
rect 20253 11384 20963 11386
rect 20253 11328 20258 11384
rect 20314 11328 20902 11384
rect 20958 11328 20963 11384
rect 20253 11326 20963 11328
rect 20253 11323 20319 11326
rect 20897 11323 20963 11326
rect 9857 11250 9923 11253
rect 17309 11250 17375 11253
rect 19425 11252 19491 11253
rect 9857 11248 17375 11250
rect 9857 11192 9862 11248
rect 9918 11192 17314 11248
rect 17370 11192 17375 11248
rect 9857 11190 17375 11192
rect 9857 11187 9923 11190
rect 17309 11187 17375 11190
rect 19374 11188 19380 11252
rect 19444 11250 19491 11252
rect 23565 11250 23631 11253
rect 27613 11250 27679 11253
rect 19444 11248 19536 11250
rect 19486 11192 19536 11248
rect 19444 11190 19536 11192
rect 23565 11248 27679 11250
rect 23565 11192 23570 11248
rect 23626 11192 27618 11248
rect 27674 11192 27679 11248
rect 23565 11190 27679 11192
rect 19444 11188 19491 11190
rect 19425 11187 19491 11188
rect 23565 11187 23631 11190
rect 27613 11187 27679 11190
rect 11605 11114 11671 11117
rect 12341 11114 12407 11117
rect 13445 11114 13511 11117
rect 11605 11112 13511 11114
rect 11605 11056 11610 11112
rect 11666 11056 12346 11112
rect 12402 11056 13450 11112
rect 13506 11056 13511 11112
rect 11605 11054 13511 11056
rect 11605 11051 11671 11054
rect 12341 11051 12407 11054
rect 13445 11051 13511 11054
rect 16573 11114 16639 11117
rect 17861 11114 17927 11117
rect 24945 11114 25011 11117
rect 26141 11114 26207 11117
rect 16573 11112 26207 11114
rect 16573 11056 16578 11112
rect 16634 11056 17866 11112
rect 17922 11056 24950 11112
rect 25006 11056 26146 11112
rect 26202 11056 26207 11112
rect 16573 11054 26207 11056
rect 16573 11051 16639 11054
rect 17861 11051 17927 11054
rect 24945 11051 25011 11054
rect 26141 11051 26207 11054
rect 10133 10978 10199 10981
rect 13261 10978 13327 10981
rect 10133 10976 13327 10978
rect 10133 10920 10138 10976
rect 10194 10920 13266 10976
rect 13322 10920 13327 10976
rect 10133 10918 13327 10920
rect 10133 10915 10199 10918
rect 13261 10915 13327 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 19517 10706 19583 10709
rect 26049 10706 26115 10709
rect 19517 10704 26115 10706
rect 19517 10648 19522 10704
rect 19578 10648 26054 10704
rect 26110 10648 26115 10704
rect 19517 10646 26115 10648
rect 19517 10643 19583 10646
rect 26049 10643 26115 10646
rect 11513 10570 11579 10573
rect 13261 10570 13327 10573
rect 11513 10568 13327 10570
rect 11513 10512 11518 10568
rect 11574 10512 13266 10568
rect 13322 10512 13327 10568
rect 11513 10510 13327 10512
rect 11513 10507 11579 10510
rect 13261 10507 13327 10510
rect 25129 10570 25195 10573
rect 26509 10570 26575 10573
rect 25129 10568 26575 10570
rect 25129 10512 25134 10568
rect 25190 10512 26514 10568
rect 26570 10512 26575 10568
rect 25129 10510 26575 10512
rect 25129 10507 25195 10510
rect 26509 10507 26575 10510
rect 4210 10368 4526 10369
rect 200 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 1577 10298 1643 10301
rect 200 10296 1643 10298
rect 200 10240 1582 10296
rect 1638 10240 1643 10296
rect 200 10238 1643 10240
rect 200 10208 800 10238
rect 1577 10235 1643 10238
rect 19333 10298 19399 10301
rect 19701 10298 19767 10301
rect 19333 10296 19767 10298
rect 19333 10240 19338 10296
rect 19394 10240 19706 10296
rect 19762 10240 19767 10296
rect 19333 10238 19767 10240
rect 19333 10235 19399 10238
rect 19701 10235 19767 10238
rect 24393 10298 24459 10301
rect 25773 10298 25839 10301
rect 24393 10296 25839 10298
rect 24393 10240 24398 10296
rect 24454 10240 25778 10296
rect 25834 10240 25839 10296
rect 24393 10238 25839 10240
rect 24393 10235 24459 10238
rect 25773 10235 25839 10238
rect 38193 10298 38259 10301
rect 39200 10298 39800 10328
rect 38193 10296 39800 10298
rect 38193 10240 38198 10296
rect 38254 10240 39800 10296
rect 38193 10238 39800 10240
rect 38193 10235 38259 10238
rect 39200 10208 39800 10238
rect 11237 10162 11303 10165
rect 13629 10162 13695 10165
rect 11237 10160 13695 10162
rect 11237 10104 11242 10160
rect 11298 10104 13634 10160
rect 13690 10104 13695 10160
rect 11237 10102 13695 10104
rect 11237 10099 11303 10102
rect 13629 10099 13695 10102
rect 18321 10162 18387 10165
rect 29269 10162 29335 10165
rect 18321 10160 29335 10162
rect 18321 10104 18326 10160
rect 18382 10104 29274 10160
rect 29330 10104 29335 10160
rect 18321 10102 29335 10104
rect 18321 10099 18387 10102
rect 29269 10099 29335 10102
rect 10501 10026 10567 10029
rect 15193 10026 15259 10029
rect 10501 10024 15259 10026
rect 10501 9968 10506 10024
rect 10562 9968 15198 10024
rect 15254 9968 15259 10024
rect 10501 9966 15259 9968
rect 10501 9963 10567 9966
rect 15193 9963 15259 9966
rect 16481 10026 16547 10029
rect 29177 10026 29243 10029
rect 16481 10024 29243 10026
rect 16481 9968 16486 10024
rect 16542 9968 29182 10024
rect 29238 9968 29243 10024
rect 16481 9966 29243 9968
rect 16481 9963 16547 9966
rect 29177 9963 29243 9966
rect 11237 9890 11303 9893
rect 14917 9890 14983 9893
rect 19241 9890 19307 9893
rect 11237 9888 19307 9890
rect 11237 9832 11242 9888
rect 11298 9832 14922 9888
rect 14978 9832 19246 9888
rect 19302 9832 19307 9888
rect 11237 9830 19307 9832
rect 11237 9827 11303 9830
rect 14917 9827 14983 9830
rect 19241 9827 19307 9830
rect 20345 9890 20411 9893
rect 27521 9890 27587 9893
rect 20345 9888 27587 9890
rect 20345 9832 20350 9888
rect 20406 9832 27526 9888
rect 27582 9832 27587 9888
rect 20345 9830 27587 9832
rect 20345 9827 20411 9830
rect 27521 9827 27587 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 17401 9754 17467 9757
rect 19425 9756 19491 9757
rect 17902 9754 17908 9756
rect 17401 9752 17908 9754
rect 17401 9696 17406 9752
rect 17462 9696 17908 9752
rect 17401 9694 17908 9696
rect 17401 9691 17467 9694
rect 17902 9692 17908 9694
rect 17972 9692 17978 9756
rect 19374 9754 19380 9756
rect 19334 9694 19380 9754
rect 19444 9752 19491 9756
rect 19486 9696 19491 9752
rect 19374 9692 19380 9694
rect 19444 9692 19491 9696
rect 19425 9691 19491 9692
rect 20161 9754 20227 9757
rect 21633 9754 21699 9757
rect 20161 9752 21699 9754
rect 20161 9696 20166 9752
rect 20222 9696 21638 9752
rect 21694 9696 21699 9752
rect 20161 9694 21699 9696
rect 20161 9691 20227 9694
rect 21633 9691 21699 9694
rect 22185 9618 22251 9621
rect 22645 9618 22711 9621
rect 22185 9616 22711 9618
rect 22185 9560 22190 9616
rect 22246 9560 22650 9616
rect 22706 9560 22711 9616
rect 22185 9558 22711 9560
rect 22185 9555 22251 9558
rect 22645 9555 22711 9558
rect 27521 9616 27587 9621
rect 27521 9560 27526 9616
rect 27582 9560 27587 9616
rect 27521 9555 27587 9560
rect 22185 9482 22251 9485
rect 23289 9482 23355 9485
rect 22185 9480 23355 9482
rect 22185 9424 22190 9480
rect 22246 9424 23294 9480
rect 23350 9424 23355 9480
rect 22185 9422 23355 9424
rect 22185 9419 22251 9422
rect 23289 9419 23355 9422
rect 21725 9346 21791 9349
rect 27524 9346 27584 9555
rect 29361 9482 29427 9485
rect 28950 9480 29427 9482
rect 28950 9424 29366 9480
rect 29422 9424 29427 9480
rect 28950 9422 29427 9424
rect 28717 9346 28783 9349
rect 28950 9346 29010 9422
rect 29361 9419 29427 9422
rect 21725 9344 29010 9346
rect 21725 9288 21730 9344
rect 21786 9288 28722 9344
rect 28778 9288 29010 9344
rect 21725 9286 29010 9288
rect 21725 9283 21791 9286
rect 28717 9283 28783 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 9305 9210 9371 9213
rect 26325 9210 26391 9213
rect 28533 9210 28599 9213
rect 9305 9208 18154 9210
rect 9305 9152 9310 9208
rect 9366 9152 18154 9208
rect 9305 9150 18154 9152
rect 9305 9147 9371 9150
rect 10869 9074 10935 9077
rect 16389 9074 16455 9077
rect 10869 9072 16455 9074
rect 10869 9016 10874 9072
rect 10930 9016 16394 9072
rect 16450 9016 16455 9072
rect 10869 9014 16455 9016
rect 18094 9074 18154 9150
rect 26325 9208 28599 9210
rect 26325 9152 26330 9208
rect 26386 9152 28538 9208
rect 28594 9152 28599 9208
rect 26325 9150 28599 9152
rect 26325 9147 26391 9150
rect 28533 9147 28599 9150
rect 19609 9074 19675 9077
rect 20662 9074 20668 9076
rect 18094 9072 20668 9074
rect 18094 9016 19614 9072
rect 19670 9016 20668 9072
rect 18094 9014 20668 9016
rect 10869 9011 10935 9014
rect 16389 9011 16455 9014
rect 19609 9011 19675 9014
rect 20662 9012 20668 9014
rect 20732 9012 20738 9076
rect 200 8938 800 8968
rect 1577 8938 1643 8941
rect 200 8936 1643 8938
rect 200 8880 1582 8936
rect 1638 8880 1643 8936
rect 200 8878 1643 8880
rect 200 8848 800 8878
rect 1577 8875 1643 8878
rect 18781 8938 18847 8941
rect 30281 8938 30347 8941
rect 18781 8936 30347 8938
rect 18781 8880 18786 8936
rect 18842 8880 30286 8936
rect 30342 8880 30347 8936
rect 18781 8878 30347 8880
rect 18781 8875 18847 8878
rect 30281 8875 30347 8878
rect 20253 8802 20319 8805
rect 22277 8802 22343 8805
rect 20253 8800 22343 8802
rect 20253 8744 20258 8800
rect 20314 8744 22282 8800
rect 22338 8744 22343 8800
rect 20253 8742 22343 8744
rect 20253 8739 20319 8742
rect 22277 8739 22343 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 11237 8532 11303 8533
rect 11237 8530 11284 8532
rect 11156 8528 11284 8530
rect 11348 8530 11354 8532
rect 17309 8530 17375 8533
rect 11348 8528 17375 8530
rect 11156 8472 11242 8528
rect 11348 8472 17314 8528
rect 17370 8472 17375 8528
rect 11156 8470 11284 8472
rect 11237 8468 11284 8470
rect 11348 8470 17375 8472
rect 11348 8468 11354 8470
rect 11237 8467 11303 8468
rect 17309 8467 17375 8470
rect 19425 8530 19491 8533
rect 21173 8530 21239 8533
rect 19425 8528 21239 8530
rect 19425 8472 19430 8528
rect 19486 8472 21178 8528
rect 21234 8472 21239 8528
rect 19425 8470 21239 8472
rect 19425 8467 19491 8470
rect 21173 8467 21239 8470
rect 22553 8394 22619 8397
rect 28717 8394 28783 8397
rect 22553 8392 28783 8394
rect 22553 8336 22558 8392
rect 22614 8336 28722 8392
rect 28778 8336 28783 8392
rect 22553 8334 28783 8336
rect 22553 8331 22619 8334
rect 28717 8331 28783 8334
rect 20713 8258 20779 8261
rect 28993 8258 29059 8261
rect 20713 8256 29059 8258
rect 20713 8200 20718 8256
rect 20774 8200 28998 8256
rect 29054 8200 29059 8256
rect 20713 8198 29059 8200
rect 20713 8195 20779 8198
rect 28993 8195 29059 8198
rect 38193 8258 38259 8261
rect 39200 8258 39800 8288
rect 38193 8256 39800 8258
rect 38193 8200 38198 8256
rect 38254 8200 39800 8256
rect 38193 8198 39800 8200
rect 38193 8195 38259 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 39200 8168 39800 8198
rect 34930 8127 35246 8128
rect 21817 8122 21883 8125
rect 22277 8122 22343 8125
rect 21817 8120 22343 8122
rect 21817 8064 21822 8120
rect 21878 8064 22282 8120
rect 22338 8064 22343 8120
rect 21817 8062 22343 8064
rect 21817 8059 21883 8062
rect 22277 8059 22343 8062
rect 14089 7986 14155 7989
rect 26325 7986 26391 7989
rect 14089 7984 26391 7986
rect 14089 7928 14094 7984
rect 14150 7928 26330 7984
rect 26386 7928 26391 7984
rect 14089 7926 26391 7928
rect 14089 7923 14155 7926
rect 26325 7923 26391 7926
rect 18045 7850 18111 7853
rect 25681 7850 25747 7853
rect 18045 7848 25747 7850
rect 18045 7792 18050 7848
rect 18106 7792 25686 7848
rect 25742 7792 25747 7848
rect 18045 7790 25747 7792
rect 18045 7787 18111 7790
rect 25681 7787 25747 7790
rect 21541 7714 21607 7717
rect 22185 7714 22251 7717
rect 21541 7712 22251 7714
rect 21541 7656 21546 7712
rect 21602 7656 22190 7712
rect 22246 7656 22251 7712
rect 21541 7654 22251 7656
rect 21541 7651 21607 7654
rect 22185 7651 22251 7654
rect 23381 7714 23447 7717
rect 27429 7714 27495 7717
rect 23381 7712 27495 7714
rect 23381 7656 23386 7712
rect 23442 7656 27434 7712
rect 27490 7656 27495 7712
rect 23381 7654 27495 7656
rect 23381 7651 23447 7654
rect 27429 7651 27495 7654
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 21265 7578 21331 7581
rect 27889 7578 27955 7581
rect 21265 7576 27955 7578
rect 21265 7520 21270 7576
rect 21326 7520 27894 7576
rect 27950 7520 27955 7576
rect 21265 7518 27955 7520
rect 21265 7515 21331 7518
rect 27889 7515 27955 7518
rect 18505 7442 18571 7445
rect 29177 7442 29243 7445
rect 18505 7440 29243 7442
rect 18505 7384 18510 7440
rect 18566 7384 29182 7440
rect 29238 7384 29243 7440
rect 18505 7382 29243 7384
rect 18505 7379 18571 7382
rect 29177 7379 29243 7382
rect 20069 7306 20135 7309
rect 30465 7306 30531 7309
rect 20069 7304 30531 7306
rect 20069 7248 20074 7304
rect 20130 7248 30470 7304
rect 30526 7248 30531 7304
rect 20069 7246 30531 7248
rect 20069 7243 20135 7246
rect 30465 7243 30531 7246
rect 15009 7170 15075 7173
rect 20437 7170 20503 7173
rect 15009 7168 20503 7170
rect 15009 7112 15014 7168
rect 15070 7112 20442 7168
rect 20498 7112 20503 7168
rect 15009 7110 20503 7112
rect 15009 7107 15075 7110
rect 20437 7107 20503 7110
rect 22369 7170 22435 7173
rect 22829 7170 22895 7173
rect 25957 7170 26023 7173
rect 22369 7168 26023 7170
rect 22369 7112 22374 7168
rect 22430 7112 22834 7168
rect 22890 7112 25962 7168
rect 26018 7112 26023 7168
rect 22369 7110 26023 7112
rect 22369 7107 22435 7110
rect 22829 7107 22895 7110
rect 25957 7107 26023 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 11145 7034 11211 7037
rect 17677 7034 17743 7037
rect 11145 7032 17743 7034
rect 11145 6976 11150 7032
rect 11206 6976 17682 7032
rect 17738 6976 17743 7032
rect 11145 6974 17743 6976
rect 11145 6971 11211 6974
rect 17677 6971 17743 6974
rect 19609 7034 19675 7037
rect 25773 7034 25839 7037
rect 19609 7032 25839 7034
rect 19609 6976 19614 7032
rect 19670 6976 25778 7032
rect 25834 6976 25839 7032
rect 19609 6974 25839 6976
rect 19609 6971 19675 6974
rect 25773 6971 25839 6974
rect 200 6898 800 6928
rect 1577 6898 1643 6901
rect 17953 6900 18019 6901
rect 200 6896 1643 6898
rect 200 6840 1582 6896
rect 1638 6840 1643 6896
rect 200 6838 1643 6840
rect 200 6808 800 6838
rect 1577 6835 1643 6838
rect 17902 6836 17908 6900
rect 17972 6898 18019 6900
rect 19425 6898 19491 6901
rect 22093 6898 22159 6901
rect 17972 6896 19258 6898
rect 18014 6840 19258 6896
rect 17972 6838 19258 6840
rect 17972 6836 18019 6838
rect 17953 6835 18019 6836
rect 19198 6762 19258 6838
rect 19425 6896 22159 6898
rect 19425 6840 19430 6896
rect 19486 6840 22098 6896
rect 22154 6840 22159 6896
rect 19425 6838 22159 6840
rect 19425 6835 19491 6838
rect 22093 6835 22159 6838
rect 22277 6898 22343 6901
rect 25405 6898 25471 6901
rect 22277 6896 25471 6898
rect 22277 6840 22282 6896
rect 22338 6840 25410 6896
rect 25466 6840 25471 6896
rect 22277 6838 25471 6840
rect 22277 6835 22343 6838
rect 25405 6835 25471 6838
rect 37917 6762 37983 6765
rect 19198 6760 37983 6762
rect 19198 6704 37922 6760
rect 37978 6704 37983 6760
rect 19198 6702 37983 6704
rect 37917 6699 37983 6702
rect 16481 6626 16547 6629
rect 17585 6626 17651 6629
rect 16481 6624 17651 6626
rect 16481 6568 16486 6624
rect 16542 6568 17590 6624
rect 17646 6568 17651 6624
rect 16481 6566 17651 6568
rect 16481 6563 16547 6566
rect 17585 6563 17651 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 15101 6490 15167 6493
rect 19333 6490 19399 6493
rect 15101 6488 19399 6490
rect 15101 6432 15106 6488
rect 15162 6432 19338 6488
rect 19394 6432 19399 6488
rect 15101 6430 19399 6432
rect 15101 6427 15167 6430
rect 19333 6427 19399 6430
rect 26509 6490 26575 6493
rect 27797 6490 27863 6493
rect 26509 6488 27863 6490
rect 26509 6432 26514 6488
rect 26570 6432 27802 6488
rect 27858 6432 27863 6488
rect 26509 6430 27863 6432
rect 26509 6427 26575 6430
rect 27797 6427 27863 6430
rect 19149 6354 19215 6357
rect 31017 6354 31083 6357
rect 19149 6352 31083 6354
rect 19149 6296 19154 6352
rect 19210 6296 31022 6352
rect 31078 6296 31083 6352
rect 19149 6294 31083 6296
rect 19149 6291 19215 6294
rect 31017 6291 31083 6294
rect 11881 6218 11947 6221
rect 16113 6218 16179 6221
rect 11881 6216 16179 6218
rect 11881 6160 11886 6216
rect 11942 6160 16118 6216
rect 16174 6160 16179 6216
rect 11881 6158 16179 6160
rect 11881 6155 11947 6158
rect 16113 6155 16179 6158
rect 38193 6218 38259 6221
rect 39200 6218 39800 6248
rect 38193 6216 39800 6218
rect 38193 6160 38198 6216
rect 38254 6160 39800 6216
rect 38193 6158 39800 6160
rect 38193 6155 38259 6158
rect 39200 6128 39800 6158
rect 10685 6082 10751 6085
rect 16665 6082 16731 6085
rect 10685 6080 16731 6082
rect 10685 6024 10690 6080
rect 10746 6024 16670 6080
rect 16726 6024 16731 6080
rect 10685 6022 16731 6024
rect 10685 6019 10751 6022
rect 16665 6019 16731 6022
rect 22553 6082 22619 6085
rect 28625 6082 28691 6085
rect 22553 6080 28691 6082
rect 22553 6024 22558 6080
rect 22614 6024 28630 6080
rect 28686 6024 28691 6080
rect 22553 6022 28691 6024
rect 22553 6019 22619 6022
rect 28625 6019 28691 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 20253 5946 20319 5949
rect 26693 5946 26759 5949
rect 20253 5944 26759 5946
rect 20253 5888 20258 5944
rect 20314 5888 26698 5944
rect 26754 5888 26759 5944
rect 20253 5886 26759 5888
rect 20253 5883 20319 5886
rect 26693 5883 26759 5886
rect 12341 5810 12407 5813
rect 27061 5810 27127 5813
rect 12341 5808 27127 5810
rect 12341 5752 12346 5808
rect 12402 5752 27066 5808
rect 27122 5752 27127 5808
rect 12341 5750 27127 5752
rect 12341 5747 12407 5750
rect 27061 5747 27127 5750
rect 22185 5674 22251 5677
rect 26509 5674 26575 5677
rect 22185 5672 26575 5674
rect 22185 5616 22190 5672
rect 22246 5616 26514 5672
rect 26570 5616 26575 5672
rect 22185 5614 26575 5616
rect 22185 5611 22251 5614
rect 26509 5611 26575 5614
rect 12249 5538 12315 5541
rect 12617 5538 12683 5541
rect 12249 5536 12683 5538
rect 12249 5480 12254 5536
rect 12310 5480 12622 5536
rect 12678 5480 12683 5536
rect 12249 5478 12683 5480
rect 12249 5475 12315 5478
rect 12617 5475 12683 5478
rect 21265 5538 21331 5541
rect 27153 5538 27219 5541
rect 21265 5536 27219 5538
rect 21265 5480 21270 5536
rect 21326 5480 27158 5536
rect 27214 5480 27219 5536
rect 21265 5478 27219 5480
rect 21265 5475 21331 5478
rect 27153 5475 27219 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 22277 5402 22343 5405
rect 27245 5402 27311 5405
rect 22277 5400 27311 5402
rect 22277 5344 22282 5400
rect 22338 5344 27250 5400
rect 27306 5344 27311 5400
rect 22277 5342 27311 5344
rect 22277 5339 22343 5342
rect 27245 5339 27311 5342
rect 16481 5266 16547 5269
rect 31109 5266 31175 5269
rect 16481 5264 31175 5266
rect 16481 5208 16486 5264
rect 16542 5208 31114 5264
rect 31170 5208 31175 5264
rect 16481 5206 31175 5208
rect 16481 5203 16547 5206
rect 31109 5203 31175 5206
rect 13721 5130 13787 5133
rect 27521 5130 27587 5133
rect 13721 5128 27587 5130
rect 13721 5072 13726 5128
rect 13782 5072 27526 5128
rect 27582 5072 27587 5128
rect 13721 5070 27587 5072
rect 13721 5067 13787 5070
rect 27521 5067 27587 5070
rect 14549 4994 14615 4997
rect 18045 4994 18111 4997
rect 14549 4992 18111 4994
rect 14549 4936 14554 4992
rect 14610 4936 18050 4992
rect 18106 4936 18111 4992
rect 14549 4934 18111 4936
rect 14549 4931 14615 4934
rect 18045 4931 18111 4934
rect 4210 4928 4526 4929
rect 200 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 1669 4858 1735 4861
rect 200 4856 1735 4858
rect 200 4800 1674 4856
rect 1730 4800 1735 4856
rect 200 4798 1735 4800
rect 200 4768 800 4798
rect 1669 4795 1735 4798
rect 20069 4858 20135 4861
rect 20662 4858 20668 4860
rect 20069 4856 20668 4858
rect 20069 4800 20074 4856
rect 20130 4800 20668 4856
rect 20069 4798 20668 4800
rect 20069 4795 20135 4798
rect 20662 4796 20668 4798
rect 20732 4796 20738 4860
rect 38285 4858 38351 4861
rect 39200 4858 39800 4888
rect 38285 4856 39800 4858
rect 38285 4800 38290 4856
rect 38346 4800 39800 4856
rect 38285 4798 39800 4800
rect 38285 4795 38351 4798
rect 39200 4768 39800 4798
rect 20529 4722 20595 4725
rect 23197 4722 23263 4725
rect 20529 4720 23263 4722
rect 20529 4664 20534 4720
rect 20590 4664 23202 4720
rect 23258 4664 23263 4720
rect 20529 4662 23263 4664
rect 20529 4659 20595 4662
rect 23197 4659 23263 4662
rect 13629 4586 13695 4589
rect 28717 4586 28783 4589
rect 13629 4584 28783 4586
rect 13629 4528 13634 4584
rect 13690 4528 28722 4584
rect 28778 4528 28783 4584
rect 13629 4526 28783 4528
rect 13629 4523 13695 4526
rect 28717 4523 28783 4526
rect 12249 4450 12315 4453
rect 13353 4450 13419 4453
rect 14641 4450 14707 4453
rect 12249 4448 14707 4450
rect 12249 4392 12254 4448
rect 12310 4392 13358 4448
rect 13414 4392 14646 4448
rect 14702 4392 14707 4448
rect 12249 4390 14707 4392
rect 12249 4387 12315 4390
rect 13353 4387 13419 4390
rect 14641 4387 14707 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 10041 4314 10107 4317
rect 14917 4314 14983 4317
rect 16849 4314 16915 4317
rect 10041 4312 16915 4314
rect 10041 4256 10046 4312
rect 10102 4256 14922 4312
rect 14978 4256 16854 4312
rect 16910 4256 16915 4312
rect 10041 4254 16915 4256
rect 10041 4251 10107 4254
rect 14917 4251 14983 4254
rect 16849 4251 16915 4254
rect 12341 4178 12407 4181
rect 14549 4180 14615 4181
rect 14549 4178 14596 4180
rect 12341 4176 14596 4178
rect 14660 4178 14666 4180
rect 22921 4178 22987 4181
rect 14660 4176 22987 4178
rect 12341 4120 12346 4176
rect 12402 4120 14554 4176
rect 14660 4120 22926 4176
rect 22982 4120 22987 4176
rect 12341 4118 14596 4120
rect 12341 4115 12407 4118
rect 14549 4116 14596 4118
rect 14660 4118 22987 4120
rect 14660 4116 14666 4118
rect 14549 4115 14615 4116
rect 22921 4115 22987 4118
rect 12433 4042 12499 4045
rect 14641 4042 14707 4045
rect 18965 4042 19031 4045
rect 12433 4040 19031 4042
rect 12433 3984 12438 4040
rect 12494 3984 14646 4040
rect 14702 3984 18970 4040
rect 19026 3984 19031 4040
rect 12433 3982 19031 3984
rect 12433 3979 12499 3982
rect 14641 3979 14707 3982
rect 18965 3979 19031 3982
rect 23473 4042 23539 4045
rect 26417 4042 26483 4045
rect 23473 4040 26483 4042
rect 23473 3984 23478 4040
rect 23534 3984 26422 4040
rect 26478 3984 26483 4040
rect 23473 3982 26483 3984
rect 23473 3979 23539 3982
rect 26417 3979 26483 3982
rect 17309 3906 17375 3909
rect 19149 3906 19215 3909
rect 17309 3904 19215 3906
rect 17309 3848 17314 3904
rect 17370 3848 19154 3904
rect 19210 3848 19215 3904
rect 17309 3846 19215 3848
rect 17309 3843 17375 3846
rect 19149 3843 19215 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 11973 3770 12039 3773
rect 12617 3770 12683 3773
rect 11973 3768 12683 3770
rect 11973 3712 11978 3768
rect 12034 3712 12622 3768
rect 12678 3712 12683 3768
rect 11973 3710 12683 3712
rect 11973 3707 12039 3710
rect 12617 3707 12683 3710
rect 23933 3634 23999 3637
rect 32949 3634 33015 3637
rect 23933 3632 33015 3634
rect 23933 3576 23938 3632
rect 23994 3576 32954 3632
rect 33010 3576 33015 3632
rect 23933 3574 33015 3576
rect 23933 3571 23999 3574
rect 32949 3571 33015 3574
rect 200 3498 800 3528
rect 1577 3498 1643 3501
rect 200 3496 1643 3498
rect 200 3440 1582 3496
rect 1638 3440 1643 3496
rect 200 3438 1643 3440
rect 200 3408 800 3438
rect 1577 3435 1643 3438
rect 17309 3498 17375 3501
rect 28349 3498 28415 3501
rect 17309 3496 28415 3498
rect 17309 3440 17314 3496
rect 17370 3440 28354 3496
rect 28410 3440 28415 3496
rect 17309 3438 28415 3440
rect 17309 3435 17375 3438
rect 28349 3435 28415 3438
rect 22461 3362 22527 3365
rect 28625 3362 28691 3365
rect 22461 3360 28691 3362
rect 22461 3304 22466 3360
rect 22522 3304 28630 3360
rect 28686 3304 28691 3360
rect 22461 3302 28691 3304
rect 22461 3299 22527 3302
rect 28625 3299 28691 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 21173 3226 21239 3229
rect 28533 3226 28599 3229
rect 21173 3224 28599 3226
rect 21173 3168 21178 3224
rect 21234 3168 28538 3224
rect 28594 3168 28599 3224
rect 21173 3166 28599 3168
rect 21173 3163 21239 3166
rect 28533 3163 28599 3166
rect 11881 3090 11947 3093
rect 13905 3090 13971 3093
rect 11881 3088 13971 3090
rect 11881 3032 11886 3088
rect 11942 3032 13910 3088
rect 13966 3032 13971 3088
rect 11881 3030 13971 3032
rect 11881 3027 11947 3030
rect 13905 3027 13971 3030
rect 23381 3090 23447 3093
rect 27061 3090 27127 3093
rect 23381 3088 27127 3090
rect 23381 3032 23386 3088
rect 23442 3032 27066 3088
rect 27122 3032 27127 3088
rect 23381 3030 27127 3032
rect 23381 3027 23447 3030
rect 27061 3027 27127 3030
rect 4613 2954 4679 2957
rect 23933 2954 23999 2957
rect 4613 2952 23999 2954
rect 4613 2896 4618 2952
rect 4674 2896 23938 2952
rect 23994 2896 23999 2952
rect 4613 2894 23999 2896
rect 4613 2891 4679 2894
rect 23933 2891 23999 2894
rect 28625 2954 28691 2957
rect 31017 2954 31083 2957
rect 28625 2952 31083 2954
rect 28625 2896 28630 2952
rect 28686 2896 31022 2952
rect 31078 2896 31083 2952
rect 28625 2894 31083 2896
rect 28625 2891 28691 2894
rect 31017 2891 31083 2894
rect 10869 2818 10935 2821
rect 12801 2818 12867 2821
rect 10869 2816 12867 2818
rect 10869 2760 10874 2816
rect 10930 2760 12806 2816
rect 12862 2760 12867 2816
rect 10869 2758 12867 2760
rect 10869 2755 10935 2758
rect 12801 2755 12867 2758
rect 38193 2818 38259 2821
rect 39200 2818 39800 2848
rect 38193 2816 39800 2818
rect 38193 2760 38198 2816
rect 38254 2760 39800 2816
rect 38193 2758 39800 2760
rect 38193 2755 38259 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 39200 2728 39800 2758
rect 34930 2687 35246 2688
rect 22001 2682 22067 2685
rect 26509 2682 26575 2685
rect 22001 2680 26575 2682
rect 22001 2624 22006 2680
rect 22062 2624 26514 2680
rect 26570 2624 26575 2680
rect 22001 2622 26575 2624
rect 22001 2619 22067 2622
rect 26509 2619 26575 2622
rect 13721 2546 13787 2549
rect 29821 2546 29887 2549
rect 13721 2544 29887 2546
rect 13721 2488 13726 2544
rect 13782 2488 29826 2544
rect 29882 2488 29887 2544
rect 13721 2486 29887 2488
rect 13721 2483 13787 2486
rect 29821 2483 29887 2486
rect 12341 2410 12407 2413
rect 29913 2410 29979 2413
rect 12341 2408 29979 2410
rect 12341 2352 12346 2408
rect 12402 2352 29918 2408
rect 29974 2352 29979 2408
rect 12341 2350 29979 2352
rect 12341 2347 12407 2350
rect 29913 2347 29979 2350
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 200 1458 800 1488
rect 1669 1458 1735 1461
rect 200 1456 1735 1458
rect 200 1400 1674 1456
rect 1730 1400 1735 1456
rect 200 1398 1735 1400
rect 200 1368 800 1398
rect 1669 1395 1735 1398
rect 37181 1458 37247 1461
rect 37181 1456 39314 1458
rect 37181 1400 37186 1456
rect 37242 1400 39314 1456
rect 37181 1398 39314 1400
rect 37181 1395 37247 1398
rect 39254 1050 39314 1398
rect 39070 990 39314 1050
rect 39070 778 39130 990
rect 39200 778 39800 808
rect 39070 718 39800 778
rect 39200 688 39800 718
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 20116 18804 20180 18868
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 14596 17036 14660 17100
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 20116 16220 20180 16284
rect 20668 15948 20732 16012
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19380 15540 19444 15604
rect 11284 15404 11348 15468
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19380 13500 19444 13564
rect 20116 13228 20180 13292
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19380 11248 19444 11252
rect 19380 11192 19430 11248
rect 19430 11192 19444 11248
rect 19380 11188 19444 11192
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 17908 9692 17972 9756
rect 19380 9752 19444 9756
rect 19380 9696 19430 9752
rect 19430 9696 19444 9752
rect 19380 9692 19444 9696
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 20668 9012 20732 9076
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 11284 8528 11348 8532
rect 11284 8472 11298 8528
rect 11298 8472 11348 8528
rect 11284 8468 11348 8472
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 17908 6896 17972 6900
rect 17908 6840 17958 6896
rect 17958 6840 17972 6896
rect 17908 6836 17972 6840
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 20668 4796 20732 4860
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 14596 4176 14660 4180
rect 14596 4120 14610 4176
rect 14610 4120 14660 4176
rect 14596 4116 14660 4120
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 20115 18868 20181 18869
rect 20115 18804 20116 18868
rect 20180 18804 20181 18868
rect 20115 18803 20181 18804
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 14595 17100 14661 17101
rect 14595 17036 14596 17100
rect 14660 17036 14661 17100
rect 14595 17035 14661 17036
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 11283 15468 11349 15469
rect 11283 15404 11284 15468
rect 11348 15404 11349 15468
rect 11283 15403 11349 15404
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 11286 8533 11346 15403
rect 11283 8532 11349 8533
rect 11283 8468 11284 8532
rect 11348 8468 11349 8532
rect 11283 8467 11349 8468
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 14598 4181 14658 17035
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19379 15604 19445 15605
rect 19379 15540 19380 15604
rect 19444 15540 19445 15604
rect 19379 15539 19445 15540
rect 19382 13565 19442 15539
rect 19568 15264 19888 16288
rect 20118 16285 20178 18803
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 20115 16284 20181 16285
rect 20115 16220 20116 16284
rect 20180 16220 20181 16284
rect 20115 16219 20181 16220
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19379 13564 19445 13565
rect 19379 13500 19380 13564
rect 19444 13500 19445 13564
rect 19379 13499 19445 13500
rect 19568 13088 19888 14112
rect 20118 13293 20178 16219
rect 20667 16012 20733 16013
rect 20667 15948 20668 16012
rect 20732 15948 20733 16012
rect 20667 15947 20733 15948
rect 20115 13292 20181 13293
rect 20115 13228 20116 13292
rect 20180 13228 20181 13292
rect 20115 13227 20181 13228
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19379 11252 19445 11253
rect 19379 11188 19380 11252
rect 19444 11188 19445 11252
rect 19379 11187 19445 11188
rect 19382 9757 19442 11187
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 17907 9756 17973 9757
rect 17907 9692 17908 9756
rect 17972 9692 17973 9756
rect 17907 9691 17973 9692
rect 19379 9756 19445 9757
rect 19379 9692 19380 9756
rect 19444 9692 19445 9756
rect 19379 9691 19445 9692
rect 17910 6901 17970 9691
rect 19568 8736 19888 9760
rect 20670 9077 20730 15947
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 20667 9076 20733 9077
rect 20667 9012 20668 9076
rect 20732 9012 20733 9076
rect 20667 9011 20733 9012
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 17907 6900 17973 6901
rect 17907 6836 17908 6900
rect 17972 6836 17973 6900
rect 17907 6835 17973 6836
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 20670 4861 20730 9011
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 20667 4860 20733 4861
rect 20667 4796 20668 4860
rect 20732 4796 20733 4860
rect 20667 4795 20733 4796
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 14595 4180 14661 4181
rect 14595 4116 14596 4180
rect 14660 4116 14661 4180
rect 14595 4115 14661 4116
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 26956 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A
timestamp 1667941163
transform 1 0 18124 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__A
timestamp 1667941163
transform -1 0 25852 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A
timestamp 1667941163
transform 1 0 17388 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__A
timestamp 1667941163
transform -1 0 23368 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A
timestamp 1667941163
transform -1 0 20148 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A
timestamp 1667941163
transform 1 0 14352 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__A
timestamp 1667941163
transform 1 0 29716 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A
timestamp 1667941163
transform 1 0 15548 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A
timestamp 1667941163
transform -1 0 24748 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__A
timestamp 1667941163
transform -1 0 29900 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__A
timestamp 1667941163
transform -1 0 28428 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__A
timestamp 1667941163
transform 1 0 18124 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A
timestamp 1667941163
transform -1 0 16284 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1667941163
transform -1 0 8096 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A
timestamp 1667941163
transform -1 0 13892 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A
timestamp 1667941163
transform -1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1667941163
transform -1 0 6992 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1667941163
transform -1 0 7544 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A
timestamp 1667941163
transform 1 0 19688 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__A
timestamp 1667941163
transform -1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A
timestamp 1667941163
transform -1 0 30452 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__A
timestamp 1667941163
transform 1 0 18124 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A
timestamp 1667941163
transform -1 0 30912 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A
timestamp 1667941163
transform -1 0 16928 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A
timestamp 1667941163
transform -1 0 30084 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__A
timestamp 1667941163
transform -1 0 29532 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A
timestamp 1667941163
transform -1 0 29256 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__A
timestamp 1667941163
transform 1 0 30176 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__A
timestamp 1667941163
transform 1 0 7820 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A
timestamp 1667941163
transform -1 0 31556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__A
timestamp 1667941163
transform -1 0 7360 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A
timestamp 1667941163
transform -1 0 9384 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__A
timestamp 1667941163
transform -1 0 23736 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A
timestamp 1667941163
transform -1 0 30452 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__A
timestamp 1667941163
transform 1 0 17756 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__A
timestamp 1667941163
transform -1 0 6808 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__A
timestamp 1667941163
transform -1 0 28980 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A
timestamp 1667941163
transform 1 0 9752 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__A
timestamp 1667941163
transform 1 0 26404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__A
timestamp 1667941163
transform -1 0 29900 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__A
timestamp 1667941163
transform 1 0 25116 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A
timestamp 1667941163
transform -1 0 9936 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__298__A
timestamp 1667941163
transform -1 0 22172 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__A
timestamp 1667941163
transform 1 0 29072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__302__A
timestamp 1667941163
transform 1 0 29072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__A
timestamp 1667941163
transform 1 0 19044 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__310__A
timestamp 1667941163
transform -1 0 29900 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__A
timestamp 1667941163
transform -1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__318__A
timestamp 1667941163
transform 1 0 22724 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__A
timestamp 1667941163
transform -1 0 15088 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__A
timestamp 1667941163
transform 1 0 22724 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__A
timestamp 1667941163
transform 1 0 28796 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__329__A
timestamp 1667941163
transform -1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__A
timestamp 1667941163
transform -1 0 29900 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__333__A
timestamp 1667941163
transform -1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__A
timestamp 1667941163
transform -1 0 8648 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__A
timestamp 1667941163
transform 1 0 11684 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__A
timestamp 1667941163
transform 1 0 8648 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__A
timestamp 1667941163
transform 1 0 8464 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A
timestamp 1667941163
transform -1 0 8096 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__A
timestamp 1667941163
transform -1 0 13340 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__A
timestamp 1667941163
transform 1 0 12328 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A
timestamp 1667941163
transform 1 0 11408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A
timestamp 1667941163
transform 1 0 12972 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__A
timestamp 1667941163
transform 1 0 9660 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A
timestamp 1667941163
transform -1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__A
timestamp 1667941163
transform -1 0 20148 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__A
timestamp 1667941163
transform -1 0 15456 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__A
timestamp 1667941163
transform 1 0 7268 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__A
timestamp 1667941163
transform -1 0 31556 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__358__A
timestamp 1667941163
transform 1 0 30820 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__A
timestamp 1667941163
transform 1 0 29624 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__A
timestamp 1667941163
transform 1 0 10028 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__A
timestamp 1667941163
transform 1 0 29716 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__362__A
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__A
timestamp 1667941163
transform 1 0 6624 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__A
timestamp 1667941163
transform -1 0 7728 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__365__A
timestamp 1667941163
transform 1 0 8096 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__A
timestamp 1667941163
transform 1 0 23644 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__A
timestamp 1667941163
transform 1 0 29624 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__A
timestamp 1667941163
transform -1 0 29808 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1667941163
transform 1 0 31188 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__371__A
timestamp 1667941163
transform 1 0 14996 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__A
timestamp 1667941163
transform -1 0 18400 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A
timestamp 1667941163
transform 1 0 20700 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__375__A
timestamp 1667941163
transform -1 0 30452 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__377__A
timestamp 1667941163
transform -1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__379__A
timestamp 1667941163
transform 1 0 22264 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__A
timestamp 1667941163
transform -1 0 16928 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__381__A
timestamp 1667941163
transform 1 0 28888 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__A
timestamp 1667941163
transform 1 0 20884 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__383__A
timestamp 1667941163
transform 1 0 28336 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1667941163
transform 1 0 9660 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__387__A
timestamp 1667941163
transform 1 0 8648 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__389__A
timestamp 1667941163
transform 1 0 17848 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__392__A
timestamp 1667941163
transform 1 0 2668 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__395__A
timestamp 1667941163
transform -1 0 7544 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__A
timestamp 1667941163
transform 1 0 33396 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__442__A
timestamp 1667941163
transform 1 0 32936 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__453__A
timestamp 1667941163
transform -1 0 33396 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__CLK
timestamp 1667941163
transform 1 0 7360 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__471__CLK
timestamp 1667941163
transform 1 0 7912 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__472__CLK
timestamp 1667941163
transform 1 0 10304 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__472__D
timestamp 1667941163
transform -1 0 10672 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__473__CLK
timestamp 1667941163
transform 1 0 17204 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__CLK
timestamp 1667941163
transform 1 0 20056 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__D
timestamp 1667941163
transform 1 0 18768 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__CLK
timestamp 1667941163
transform 1 0 34132 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__D
timestamp 1667941163
transform -1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__RESET_B
timestamp 1667941163
transform 1 0 33580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__476__CLK
timestamp 1667941163
transform 1 0 30268 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__477__CLK
timestamp 1667941163
transform 1 0 33488 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__CLK
timestamp 1667941163
transform 1 0 25668 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__D
timestamp 1667941163
transform -1 0 26588 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__479__CLK
timestamp 1667941163
transform 1 0 10212 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__CLK
timestamp 1667941163
transform 1 0 11684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__D
timestamp 1667941163
transform 1 0 9200 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__481__CLK
timestamp 1667941163
transform 1 0 27600 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__CLK
timestamp 1667941163
transform 1 0 11408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__483__CLK
timestamp 1667941163
transform 1 0 10856 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__CLK
timestamp 1667941163
transform 1 0 9936 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__D
timestamp 1667941163
transform -1 0 10488 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__485__CLK
timestamp 1667941163
transform 1 0 20240 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__CLK
timestamp 1667941163
transform 1 0 20792 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__487__CLK
timestamp 1667941163
transform 1 0 25300 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__488__CLK
timestamp 1667941163
transform 1 0 9200 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__489__CLK
timestamp 1667941163
transform 1 0 7912 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__CLK
timestamp 1667941163
transform 1 0 11040 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__D
timestamp 1667941163
transform -1 0 10672 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__491__CLK
timestamp 1667941163
transform 1 0 14996 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__CLK
timestamp 1667941163
transform 1 0 20608 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__CLK
timestamp 1667941163
transform 1 0 23552 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__CLK
timestamp 1667941163
transform 1 0 29716 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__495__CLK
timestamp 1667941163
transform 1 0 30636 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__CLK
timestamp 1667941163
transform 1 0 29532 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__D
timestamp 1667941163
transform -1 0 34408 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__CLK
timestamp 1667941163
transform 1 0 24748 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__D
timestamp 1667941163
transform -1 0 27416 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__CLK
timestamp 1667941163
transform 1 0 24288 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__499__CLK
timestamp 1667941163
transform 1 0 20516 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__500__CLK
timestamp 1667941163
transform 1 0 7636 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__501__CLK
timestamp 1667941163
transform 1 0 8280 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__502__CLK
timestamp 1667941163
transform 1 0 10856 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__502__D
timestamp 1667941163
transform -1 0 10488 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__503__CLK
timestamp 1667941163
transform 1 0 21344 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__504__CLK
timestamp 1667941163
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__504__D
timestamp 1667941163
transform -1 0 10672 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__505__CLK
timestamp 1667941163
transform 1 0 28980 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__506__CLK
timestamp 1667941163
transform 1 0 9936 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__507__CLK
timestamp 1667941163
transform 1 0 9752 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__508__CLK
timestamp 1667941163
transform 1 0 11040 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__509__CLK
timestamp 1667941163
transform 1 0 11408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__509__D
timestamp 1667941163
transform -1 0 11040 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__510__CLK
timestamp 1667941163
transform 1 0 13892 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__510__D
timestamp 1667941163
transform 1 0 14444 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__511__CLK
timestamp 1667941163
transform 1 0 11408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__512__CLK
timestamp 1667941163
transform 1 0 10488 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__512__D
timestamp 1667941163
transform -1 0 11040 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__513__CLK
timestamp 1667941163
transform 1 0 9660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__513__D
timestamp 1667941163
transform -1 0 9292 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__514__CLK
timestamp 1667941163
transform 1 0 25116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__514__D
timestamp 1667941163
transform -1 0 11960 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__515__CLK
timestamp 1667941163
transform 1 0 19412 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__516__CLK
timestamp 1667941163
transform 1 0 11960 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__517__CLK
timestamp 1667941163
transform 1 0 12052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__518__CLK
timestamp 1667941163
transform 1 0 11408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__519__CLK
timestamp 1667941163
transform 1 0 10212 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__519__D
timestamp 1667941163
transform 1 0 8740 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__520__CLK
timestamp 1667941163
transform 1 0 8188 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__520__D
timestamp 1667941163
transform -1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__521__CLK
timestamp 1667941163
transform 1 0 20976 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__522__CLK
timestamp 1667941163
transform 1 0 24196 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__523__CLK
timestamp 1667941163
transform 1 0 14352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__523__D
timestamp 1667941163
transform -1 0 11960 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__524__CLK
timestamp 1667941163
transform 1 0 27784 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__524__D
timestamp 1667941163
transform -1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__525__CLK
timestamp 1667941163
transform 1 0 26220 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__CLK
timestamp 1667941163
transform 1 0 24564 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__527__CLK
timestamp 1667941163
transform 1 0 23736 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__527__D
timestamp 1667941163
transform -1 0 25576 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__528__CLK
timestamp 1667941163
transform 1 0 16836 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__528__D
timestamp 1667941163
transform -1 0 12788 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__529__CLK
timestamp 1667941163
transform 1 0 28428 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__529__D
timestamp 1667941163
transform 1 0 10304 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__530__CLK
timestamp 1667941163
transform 1 0 11040 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__531__CLK
timestamp 1667941163
transform 1 0 10488 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__532__CLK
timestamp 1667941163
transform 1 0 8832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__532__D
timestamp 1667941163
transform -1 0 9568 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__533__CLK
timestamp 1667941163
transform 1 0 9384 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__533__D
timestamp 1667941163
transform -1 0 9936 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__534__CLK
timestamp 1667941163
transform 1 0 10764 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__534__D
timestamp 1667941163
transform -1 0 31188 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__535__CLK
timestamp 1667941163
transform 1 0 21344 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__547__A
timestamp 1667941163
transform -1 0 18216 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__548__A
timestamp 1667941163
transform -1 0 8832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__549__A
timestamp 1667941163
transform 1 0 7176 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__551__A
timestamp 1667941163
transform 1 0 22632 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__552__A
timestamp 1667941163
transform 1 0 19504 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__553__A
timestamp 1667941163
transform 1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__554__A
timestamp 1667941163
transform -1 0 8096 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__555__A
timestamp 1667941163
transform -1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__557__A
timestamp 1667941163
transform 1 0 23552 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__558__A
timestamp 1667941163
transform -1 0 22908 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__559__A
timestamp 1667941163
transform 1 0 22816 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__560__A
timestamp 1667941163
transform -1 0 30268 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__561__A
timestamp 1667941163
transform 1 0 14720 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__563__A
timestamp 1667941163
transform -1 0 30544 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__565__A
timestamp 1667941163
transform -1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__566__A
timestamp 1667941163
transform -1 0 9384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__567__A
timestamp 1667941163
transform -1 0 28980 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__570__A
timestamp 1667941163
transform 1 0 2576 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__571__A
timestamp 1667941163
transform 1 0 5244 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__572__A
timestamp 1667941163
transform -1 0 38272 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__573__A
timestamp 1667941163
transform -1 0 3128 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__574__A
timestamp 1667941163
transform -1 0 20884 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__575__A
timestamp 1667941163
transform -1 0 31004 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__576__A
timestamp 1667941163
transform 1 0 15640 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__579__A
timestamp 1667941163
transform 1 0 31188 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__580__A
timestamp 1667941163
transform 1 0 11960 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__581__A
timestamp 1667941163
transform 1 0 20424 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__582__A
timestamp 1667941163
transform -1 0 27324 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__583__A
timestamp 1667941163
transform -1 0 28060 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__584__A
timestamp 1667941163
transform 1 0 26312 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__611__A
timestamp 1667941163
transform 1 0 23000 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__653__A
timestamp 1667941163
transform -1 0 7360 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__683__A
timestamp 1667941163
transform -1 0 29256 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1667941163
transform -1 0 2392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1667941163
transform -1 0 1748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1667941163
transform -1 0 36064 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1667941163
transform -1 0 14536 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1667941163
transform -1 0 16376 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1667941163
transform -1 0 17756 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1667941163
transform -1 0 10120 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1667941163
transform -1 0 37628 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1667941163
transform -1 0 35144 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1667941163
transform -1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1667941163
transform -1 0 7268 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1667941163
transform -1 0 37628 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1667941163
transform -1 0 37628 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1667941163
transform -1 0 38364 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1667941163
transform -1 0 38364 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1667941163
transform -1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1667941163
transform -1 0 1748 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1667941163
transform -1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1667941163
transform -1 0 38364 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1667941163
transform -1 0 1748 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1667941163
transform -1 0 37628 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1667941163
transform -1 0 3220 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1667941163
transform -1 0 1748 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1667941163
transform -1 0 1748 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1667941163
transform -1 0 1748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1667941163
transform -1 0 36984 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1667941163
transform -1 0 7452 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1667941163
transform -1 0 4140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1667941163
transform -1 0 6716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1667941163
transform -1 0 35512 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1667941163
transform -1 0 37628 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1667941163
transform -1 0 37628 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1667941163
transform -1 0 34224 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1667941163
transform -1 0 2484 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1667941163
transform -1 0 37628 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1667941163
transform -1 0 1748 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1667941163
transform -1 0 37628 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1667941163
transform -1 0 1748 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1667941163
transform -1 0 34960 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1667941163
transform -1 0 37628 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output41_A
timestamp 1667941163
transform -1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output43_A
timestamp 1667941163
transform 1 0 37444 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output52_A
timestamp 1667941163
transform 1 0 2300 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output55_A
timestamp 1667941163
transform -1 0 35052 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output57_A
timestamp 1667941163
transform 1 0 37444 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output61_A
timestamp 1667941163
transform 1 0 37444 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output62_A
timestamp 1667941163
transform -1 0 12604 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output65_A
timestamp 1667941163
transform 1 0 2668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output66_A
timestamp 1667941163
transform -1 0 33120 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output72_A
timestamp 1667941163
transform 1 0 3220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output76_A
timestamp 1667941163
transform -1 0 36892 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output78_A
timestamp 1667941163
transform -1 0 5520 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output79_A
timestamp 1667941163
transform 1 0 37444 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17
timestamp 1667941163
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3036 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33
timestamp 1667941163
transform 1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37
timestamp 1667941163
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4968 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50
timestamp 1667941163
transform 1 0 5704 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1667941163
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1667941163
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67
timestamp 1667941163
transform 1 0 7268 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70
timestamp 1667941163
transform 1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76
timestamp 1667941163
transform 1 0 8096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91
timestamp 1667941163
transform 1 0 9476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_98
timestamp 1667941163
transform 1 0 10120 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1667941163
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117
timestamp 1667941163
transform 1 0 11868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp 1667941163
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1667941163
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_173
timestamp 1667941163
transform 1 0 17020 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1667941163
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1667941163
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1667941163
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1667941163
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_275
timestamp 1667941163
transform 1 0 26404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1667941163
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_287
timestamp 1667941163
transform 1 0 27508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_295
timestamp 1667941163
transform 1 0 28244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_302 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 28888 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_314
timestamp 1667941163
transform 1 0 29992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_322
timestamp 1667941163
transform 1 0 30728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_329
timestamp 1667941163
transform 1 0 31372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1667941163
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_342
timestamp 1667941163
transform 1 0 32568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1667941163
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_355
timestamp 1667941163
transform 1 0 33764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_371
timestamp 1667941163
transform 1 0 35236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_379
timestamp 1667941163
transform 1 0 35972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_385
timestamp 1667941163
transform 1 0 36524 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1667941163
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_399
timestamp 1667941163
transform 1 0 37812 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_19
timestamp 1667941163
transform 1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_25
timestamp 1667941163
transform 1 0 3404 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_33
timestamp 1667941163
transform 1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_39
timestamp 1667941163
transform 1 0 4692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_46
timestamp 1667941163
transform 1 0 5336 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_61
timestamp 1667941163
transform 1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_67
timestamp 1667941163
transform 1 0 7268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_73
timestamp 1667941163
transform 1 0 7820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_79
timestamp 1667941163
transform 1 0 8372 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_85
timestamp 1667941163
transform 1 0 8924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_92
timestamp 1667941163
transform 1 0 9568 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_102
timestamp 1667941163
transform 1 0 10488 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1667941163
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_118
timestamp 1667941163
transform 1 0 11960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_142
timestamp 1667941163
transform 1 0 14168 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1667941163
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1667941163
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1667941163
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_250
timestamp 1667941163
transform 1 0 24104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_274
timestamp 1667941163
transform 1 0 26312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_287
timestamp 1667941163
transform 1 0 27508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_294
timestamp 1667941163
transform 1 0 28152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_301
timestamp 1667941163
transform 1 0 28796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_308
timestamp 1667941163
transform 1 0 29440 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_315
timestamp 1667941163
transform 1 0 30084 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_322
timestamp 1667941163
transform 1 0 30728 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1667941163
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_342
timestamp 1667941163
transform 1 0 32568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_356
timestamp 1667941163
transform 1 0 33856 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_362
timestamp 1667941163
transform 1 0 34408 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_368
timestamp 1667941163
transform 1 0 34960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_374
timestamp 1667941163
transform 1 0 35512 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_380 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 36064 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_8
timestamp 1667941163
transform 1 0 1840 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_14
timestamp 1667941163
transform 1 0 2392 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1667941163
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_37
timestamp 1667941163
transform 1 0 4508 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_65
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_70
timestamp 1667941163
transform 1 0 7544 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_76
timestamp 1667941163
transform 1 0 8096 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1667941163
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_89
timestamp 1667941163
transform 1 0 9292 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_95
timestamp 1667941163
transform 1 0 9844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_101
timestamp 1667941163
transform 1 0 10396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_107
timestamp 1667941163
transform 1 0 10948 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_114
timestamp 1667941163
transform 1 0 11592 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1667941163
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_167
timestamp 1667941163
transform 1 0 16468 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1667941163
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_203
timestamp 1667941163
transform 1 0 19780 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_211
timestamp 1667941163
transform 1 0 20516 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_215
timestamp 1667941163
transform 1 0 20884 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_239
timestamp 1667941163
transform 1 0 23092 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp 1667941163
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1667941163
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_275
timestamp 1667941163
transform 1 0 26404 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_282
timestamp 1667941163
transform 1 0 27048 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_296
timestamp 1667941163
transform 1 0 28336 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_303
timestamp 1667941163
transform 1 0 28980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_314
timestamp 1667941163
transform 1 0 29992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_328
timestamp 1667941163
transform 1 0 31280 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_335
timestamp 1667941163
transform 1 0 31924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_342
timestamp 1667941163
transform 1 0 32568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_348
timestamp 1667941163
transform 1 0 33120 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_354
timestamp 1667941163
transform 1 0 33672 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1667941163
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_369
timestamp 1667941163
transform 1 0 35052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_381
timestamp 1667941163
transform 1 0 36156 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_393
timestamp 1667941163
transform 1 0 37260 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_397
timestamp 1667941163
transform 1 0 37628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1667941163
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1667941163
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1667941163
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1667941163
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_77
timestamp 1667941163
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_80
timestamp 1667941163
transform 1 0 8464 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_86
timestamp 1667941163
transform 1 0 9016 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_92
timestamp 1667941163
transform 1 0 9568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_98
timestamp 1667941163
transform 1 0 10120 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_104
timestamp 1667941163
transform 1 0 10672 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1667941163
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_139
timestamp 1667941163
transform 1 0 13892 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1667941163
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1667941163
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_213
timestamp 1667941163
transform 1 0 20700 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_219
timestamp 1667941163
transform 1 0 21252 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1667941163
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_247
timestamp 1667941163
transform 1 0 23828 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_271
timestamp 1667941163
transform 1 0 26036 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_277
timestamp 1667941163
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_285
timestamp 1667941163
transform 1 0 27324 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_289
timestamp 1667941163
transform 1 0 27692 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_296
timestamp 1667941163
transform 1 0 28336 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_307
timestamp 1667941163
transform 1 0 29348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_314
timestamp 1667941163
transform 1 0 29992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_321
timestamp 1667941163
transform 1 0 30636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_328
timestamp 1667941163
transform 1 0 31280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1667941163
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_345
timestamp 1667941163
transform 1 0 32844 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_351
timestamp 1667941163
transform 1 0 33396 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_363
timestamp 1667941163
transform 1 0 34500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_375
timestamp 1667941163
transform 1 0 35604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_387
timestamp 1667941163
transform 1 0 36708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1667941163
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_90
timestamp 1667941163
transform 1 0 9384 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_96
timestamp 1667941163
transform 1 0 9936 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_102
timestamp 1667941163
transform 1 0 10488 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_108
timestamp 1667941163
transform 1 0 11040 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_114
timestamp 1667941163
transform 1 0 11592 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1667941163
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_167
timestamp 1667941163
transform 1 0 16468 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_173
timestamp 1667941163
transform 1 0 17020 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1667941163
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_201
timestamp 1667941163
transform 1 0 19596 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_207
timestamp 1667941163
transform 1 0 20148 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1667941163
transform 1 0 20700 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_216
timestamp 1667941163
transform 1 0 20976 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_240
timestamp 1667941163
transform 1 0 23184 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_246
timestamp 1667941163
transform 1 0 23736 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_257
timestamp 1667941163
transform 1 0 24748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_263
timestamp 1667941163
transform 1 0 25300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_269
timestamp 1667941163
transform 1 0 25852 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_275
timestamp 1667941163
transform 1 0 26404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_284
timestamp 1667941163
transform 1 0 27232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_290
timestamp 1667941163
transform 1 0 27784 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_294
timestamp 1667941163
transform 1 0 28152 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_298
timestamp 1667941163
transform 1 0 28520 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_302
timestamp 1667941163
transform 1 0 28888 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1667941163
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_314
timestamp 1667941163
transform 1 0 29992 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_327
timestamp 1667941163
transform 1 0 31188 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_335
timestamp 1667941163
transform 1 0 31924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_342
timestamp 1667941163
transform 1 0 32568 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_348
timestamp 1667941163
transform 1 0 33120 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_360
timestamp 1667941163
transform 1 0 34224 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_401
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1667941163
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_9
timestamp 1667941163
transform 1 0 1932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_21
timestamp 1667941163
transform 1 0 3036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_33
timestamp 1667941163
transform 1 0 4140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_45
timestamp 1667941163
transform 1 0 5244 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1667941163
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_89
timestamp 1667941163
transform 1 0 9292 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_92
timestamp 1667941163
transform 1 0 9568 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_98
timestamp 1667941163
transform 1 0 10120 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_104
timestamp 1667941163
transform 1 0 10672 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1667941163
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1667941163
transform 1 0 11960 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_142
timestamp 1667941163
transform 1 0 14168 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1667941163
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_173
timestamp 1667941163
transform 1 0 17020 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_197
timestamp 1667941163
transform 1 0 19228 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_221
timestamp 1667941163
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_247
timestamp 1667941163
transform 1 0 23828 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_253
timestamp 1667941163
transform 1 0 24380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_259
timestamp 1667941163
transform 1 0 24932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_265
timestamp 1667941163
transform 1 0 25484 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_277
timestamp 1667941163
transform 1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_286
timestamp 1667941163
transform 1 0 27416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_299
timestamp 1667941163
transform 1 0 28612 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_303
timestamp 1667941163
transform 1 0 28980 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_310
timestamp 1667941163
transform 1 0 29624 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_323
timestamp 1667941163
transform 1 0 30820 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1667941163
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1667941163
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1667941163
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1667941163
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_93
timestamp 1667941163
transform 1 0 9660 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_96
timestamp 1667941163
transform 1 0 9936 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_102
timestamp 1667941163
transform 1 0 10488 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_108
timestamp 1667941163
transform 1 0 11040 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_114
timestamp 1667941163
transform 1 0 11592 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1667941163
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_146
timestamp 1667941163
transform 1 0 14536 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_170
timestamp 1667941163
transform 1 0 16744 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1667941163
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_201
timestamp 1667941163
transform 1 0 19596 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_204
timestamp 1667941163
transform 1 0 19872 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_210
timestamp 1667941163
transform 1 0 20424 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_218
timestamp 1667941163
transform 1 0 21160 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_242
timestamp 1667941163
transform 1 0 23368 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_248
timestamp 1667941163
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_258
timestamp 1667941163
transform 1 0 24840 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_266
timestamp 1667941163
transform 1 0 25576 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_270
timestamp 1667941163
transform 1 0 25944 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1667941163
transform 1 0 26496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_280
timestamp 1667941163
transform 1 0 26864 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_286
timestamp 1667941163
transform 1 0 27416 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_292
timestamp 1667941163
transform 1 0 27968 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_303
timestamp 1667941163
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_313
timestamp 1667941163
transform 1 0 29900 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_319
timestamp 1667941163
transform 1 0 30452 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_325
timestamp 1667941163
transform 1 0 31004 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_337
timestamp 1667941163
transform 1 0 32108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_349
timestamp 1667941163
transform 1 0 33212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_361
timestamp 1667941163
transform 1 0 34316 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_401
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1667941163
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1667941163
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_98
timestamp 1667941163
transform 1 0 10120 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_104
timestamp 1667941163
transform 1 0 10672 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1667941163
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1667941163
transform 1 0 11960 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_142
timestamp 1667941163
transform 1 0 14168 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1667941163
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_177
timestamp 1667941163
transform 1 0 17388 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_202
timestamp 1667941163
transform 1 0 19688 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_210
timestamp 1667941163
transform 1 0 20424 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_213
timestamp 1667941163
transform 1 0 20700 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp 1667941163
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_248
timestamp 1667941163
transform 1 0 23920 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_256
timestamp 1667941163
transform 1 0 24656 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_260
timestamp 1667941163
transform 1 0 25024 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_266
timestamp 1667941163
transform 1 0 25576 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_270
timestamp 1667941163
transform 1 0 25944 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_274
timestamp 1667941163
transform 1 0 26312 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_286
timestamp 1667941163
transform 1 0 27416 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_299
timestamp 1667941163
transform 1 0 28612 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_311
timestamp 1667941163
transform 1 0 29716 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_397
timestamp 1667941163
transform 1 0 37628 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7
timestamp 1667941163
transform 1 0 1748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_19
timestamp 1667941163
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1667941163
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_102
timestamp 1667941163
transform 1 0 10488 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_108
timestamp 1667941163
transform 1 0 11040 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_114
timestamp 1667941163
transform 1 0 11592 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1667941163
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_147
timestamp 1667941163
transform 1 0 14628 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_178
timestamp 1667941163
transform 1 0 17480 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_184
timestamp 1667941163
transform 1 0 18032 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1667941163
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_202
timestamp 1667941163
transform 1 0 19688 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_208
timestamp 1667941163
transform 1 0 20240 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_214
timestamp 1667941163
transform 1 0 20792 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_239
timestamp 1667941163
transform 1 0 23092 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1667941163
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_257
timestamp 1667941163
transform 1 0 24748 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_261
timestamp 1667941163
transform 1 0 25116 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_268
timestamp 1667941163
transform 1 0 25760 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1667941163
transform 1 0 26496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_280
timestamp 1667941163
transform 1 0 26864 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_287
timestamp 1667941163
transform 1 0 27508 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_294
timestamp 1667941163
transform 1 0 28152 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_302
timestamp 1667941163
transform 1 0 28888 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1667941163
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_9
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_21
timestamp 1667941163
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_33
timestamp 1667941163
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_45
timestamp 1667941163
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1667941163
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_101
timestamp 1667941163
transform 1 0 10396 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_104
timestamp 1667941163
transform 1 0 10672 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1667941163
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_121
timestamp 1667941163
transform 1 0 12236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_127
timestamp 1667941163
transform 1 0 12788 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_134
timestamp 1667941163
transform 1 0 13432 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_138
timestamp 1667941163
transform 1 0 13800 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_141
timestamp 1667941163
transform 1 0 14076 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1667941163
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_174
timestamp 1667941163
transform 1 0 17112 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_188
timestamp 1667941163
transform 1 0 18400 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_213
timestamp 1667941163
transform 1 0 20700 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_219
timestamp 1667941163
transform 1 0 21252 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1667941163
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_248
timestamp 1667941163
transform 1 0 23920 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_255
timestamp 1667941163
transform 1 0 24564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_262
timestamp 1667941163
transform 1 0 25208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_269
timestamp 1667941163
transform 1 0 25852 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1667941163
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_286
timestamp 1667941163
transform 1 0 27416 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_300
timestamp 1667941163
transform 1 0 28704 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_307
timestamp 1667941163
transform 1 0 29348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_314
timestamp 1667941163
transform 1 0 29992 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_321
timestamp 1667941163
transform 1 0 30636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp 1667941163
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1667941163
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1667941163
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1667941163
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1667941163
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_105
timestamp 1667941163
transform 1 0 10764 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_108
timestamp 1667941163
transform 1 0 11040 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_114
timestamp 1667941163
transform 1 0 11592 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_120
timestamp 1667941163
transform 1 0 12144 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_127
timestamp 1667941163
transform 1 0 12788 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_134
timestamp 1667941163
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_145
timestamp 1667941163
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_167
timestamp 1667941163
transform 1 0 16468 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1667941163
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_220
timestamp 1667941163
transform 1 0 21344 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_260
timestamp 1667941163
transform 1 0 25024 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_267
timestamp 1667941163
transform 1 0 25668 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_274
timestamp 1667941163
transform 1 0 26312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_281
timestamp 1667941163
transform 1 0 26956 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_288
timestamp 1667941163
transform 1 0 27600 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_295
timestamp 1667941163
transform 1 0 28244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_302
timestamp 1667941163
transform 1 0 28888 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_314
timestamp 1667941163
transform 1 0 29992 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_401
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_7
timestamp 1667941163
transform 1 0 1748 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_15
timestamp 1667941163
transform 1 0 2484 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_20
timestamp 1667941163
transform 1 0 2944 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_32
timestamp 1667941163
transform 1 0 4048 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_44
timestamp 1667941163
transform 1 0 5152 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_101
timestamp 1667941163
transform 1 0 10396 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_104
timestamp 1667941163
transform 1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1667941163
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_117
timestamp 1667941163
transform 1 0 11868 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_141
timestamp 1667941163
transform 1 0 14076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1667941163
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_175
timestamp 1667941163
transform 1 0 17204 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_179
timestamp 1667941163
transform 1 0 17572 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_206
timestamp 1667941163
transform 1 0 20056 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_213
timestamp 1667941163
transform 1 0 20700 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp 1667941163
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_248
timestamp 1667941163
transform 1 0 23920 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_254
timestamp 1667941163
transform 1 0 24472 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_267
timestamp 1667941163
transform 1 0 25668 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_274
timestamp 1667941163
transform 1 0 26312 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_286
timestamp 1667941163
transform 1 0 27416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_300
timestamp 1667941163
transform 1 0 28704 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_307
timestamp 1667941163
transform 1 0 29348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_314
timestamp 1667941163
transform 1 0 29992 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_321
timestamp 1667941163
transform 1 0 30636 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_333
timestamp 1667941163
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_397
timestamp 1667941163
transform 1 0 37628 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1667941163
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_95
timestamp 1667941163
transform 1 0 9844 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_101
timestamp 1667941163
transform 1 0 10396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_108
timestamp 1667941163
transform 1 0 11040 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_115
timestamp 1667941163
transform 1 0 11684 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_128
timestamp 1667941163
transform 1 0 12880 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_134
timestamp 1667941163
transform 1 0 13432 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1667941163
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_167
timestamp 1667941163
transform 1 0 16468 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1667941163
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_202
timestamp 1667941163
transform 1 0 19688 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_206
timestamp 1667941163
transform 1 0 20056 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_210
timestamp 1667941163
transform 1 0 20424 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_217
timestamp 1667941163
transform 1 0 21068 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_221
timestamp 1667941163
transform 1 0 21436 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_258
timestamp 1667941163
transform 1 0 24840 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_266
timestamp 1667941163
transform 1 0 25576 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_276
timestamp 1667941163
transform 1 0 26496 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_289
timestamp 1667941163
transform 1 0 27692 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_296
timestamp 1667941163
transform 1 0 28336 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_303
timestamp 1667941163
transform 1 0 28980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1667941163
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_317
timestamp 1667941163
transform 1 0 30268 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_323
timestamp 1667941163
transform 1 0 30820 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_335
timestamp 1667941163
transform 1 0 31924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_347
timestamp 1667941163
transform 1 0 33028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_353
timestamp 1667941163
transform 1 0 33580 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_361
timestamp 1667941163
transform 1 0 34316 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_401
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1667941163
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1667941163
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1667941163
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1667941163
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_84
timestamp 1667941163
transform 1 0 8832 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_90
timestamp 1667941163
transform 1 0 9384 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_96
timestamp 1667941163
transform 1 0 9936 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_103
timestamp 1667941163
transform 1 0 10580 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1667941163
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_119
timestamp 1667941163
transform 1 0 12052 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_132
timestamp 1667941163
transform 1 0 13248 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_141
timestamp 1667941163
transform 1 0 14076 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1667941163
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_208
timestamp 1667941163
transform 1 0 20240 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_215
timestamp 1667941163
transform 1 0 20884 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1667941163
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_248
timestamp 1667941163
transform 1 0 23920 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_255
timestamp 1667941163
transform 1 0 24564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_268
timestamp 1667941163
transform 1 0 25760 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_275
timestamp 1667941163
transform 1 0 26404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_286
timestamp 1667941163
transform 1 0 27416 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_299
timestamp 1667941163
transform 1 0 28612 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_313
timestamp 1667941163
transform 1 0 29900 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_319
timestamp 1667941163
transform 1 0 30452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_325
timestamp 1667941163
transform 1 0 31004 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_331
timestamp 1667941163
transform 1 0 31556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_357
timestamp 1667941163
transform 1 0 33948 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_363
timestamp 1667941163
transform 1 0 34500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_375
timestamp 1667941163
transform 1 0 35604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_387
timestamp 1667941163
transform 1 0 36708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_7
timestamp 1667941163
transform 1 0 1748 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_19
timestamp 1667941163
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1667941163
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_77
timestamp 1667941163
transform 1 0 8188 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1667941163
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_90
timestamp 1667941163
transform 1 0 9384 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_104
timestamp 1667941163
transform 1 0 10672 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_111
timestamp 1667941163
transform 1 0 11316 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_124
timestamp 1667941163
transform 1 0 12512 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1667941163
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1667941163
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_167
timestamp 1667941163
transform 1 0 16468 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1667941163
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_202
timestamp 1667941163
transform 1 0 19688 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_208
timestamp 1667941163
transform 1 0 20240 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_218
timestamp 1667941163
transform 1 0 21160 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_222
timestamp 1667941163
transform 1 0 21528 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_244
timestamp 1667941163
transform 1 0 23552 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1667941163
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_257
timestamp 1667941163
transform 1 0 24748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_271
timestamp 1667941163
transform 1 0 26036 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_284
timestamp 1667941163
transform 1 0 27232 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_291
timestamp 1667941163
transform 1 0 27876 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_297
timestamp 1667941163
transform 1 0 28428 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1667941163
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_317
timestamp 1667941163
transform 1 0 30268 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_329
timestamp 1667941163
transform 1 0 31372 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_341
timestamp 1667941163
transform 1 0 32476 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_353
timestamp 1667941163
transform 1 0 33580 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_361
timestamp 1667941163
transform 1 0 34316 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_9
timestamp 1667941163
transform 1 0 1932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_21
timestamp 1667941163
transform 1 0 3036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_33
timestamp 1667941163
transform 1 0 4140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp 1667941163
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1667941163
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_75
timestamp 1667941163
transform 1 0 8004 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_78
timestamp 1667941163
transform 1 0 8280 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_84
timestamp 1667941163
transform 1 0 8832 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_92
timestamp 1667941163
transform 1 0 9568 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_96
timestamp 1667941163
transform 1 0 9936 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_103
timestamp 1667941163
transform 1 0 10580 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1667941163
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_117
timestamp 1667941163
transform 1 0 11868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_127
timestamp 1667941163
transform 1 0 12788 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_140
timestamp 1667941163
transform 1 0 13984 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1667941163
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1667941163
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1667941163
transform 1 0 19136 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_200
timestamp 1667941163
transform 1 0 19504 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1667941163
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_248
timestamp 1667941163
transform 1 0 23920 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_261
timestamp 1667941163
transform 1 0 25116 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_274
timestamp 1667941163
transform 1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_292
timestamp 1667941163
transform 1 0 27968 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_296
timestamp 1667941163
transform 1 0 28336 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_303
timestamp 1667941163
transform 1 0 28980 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_309
timestamp 1667941163
transform 1 0 29532 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_315
timestamp 1667941163
transform 1 0 30084 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_327
timestamp 1667941163
transform 1 0 31188 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1667941163
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_397
timestamp 1667941163
transform 1 0 37628 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1667941163
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1667941163
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_73
timestamp 1667941163
transform 1 0 7820 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_76
timestamp 1667941163
transform 1 0 8096 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1667941163
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_90
timestamp 1667941163
transform 1 0 9384 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_103
timestamp 1667941163
transform 1 0 10580 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_112
timestamp 1667941163
transform 1 0 11408 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_125
timestamp 1667941163
transform 1 0 12604 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1667941163
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_151
timestamp 1667941163
transform 1 0 14996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_164
timestamp 1667941163
transform 1 0 16192 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1667941163
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_207
timestamp 1667941163
transform 1 0 20148 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_220
timestamp 1667941163
transform 1 0 21344 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_233
timestamp 1667941163
transform 1 0 22540 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_246
timestamp 1667941163
transform 1 0 23736 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_264
timestamp 1667941163
transform 1 0 25392 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_277
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_290
timestamp 1667941163
transform 1 0 27784 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_297
timestamp 1667941163
transform 1 0 28428 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_303
timestamp 1667941163
transform 1 0 28980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1667941163
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_313
timestamp 1667941163
transform 1 0 29900 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_325
timestamp 1667941163
transform 1 0 31004 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_337
timestamp 1667941163
transform 1 0 32108 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_349
timestamp 1667941163
transform 1 0 33212 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_361
timestamp 1667941163
transform 1 0 34316 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_401
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_65
timestamp 1667941163
transform 1 0 7084 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_75
timestamp 1667941163
transform 1 0 8004 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_82
timestamp 1667941163
transform 1 0 8648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_89
timestamp 1667941163
transform 1 0 9292 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_96
timestamp 1667941163
transform 1 0 9936 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_103
timestamp 1667941163
transform 1 0 10580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1667941163
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_117
timestamp 1667941163
transform 1 0 11868 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_121
timestamp 1667941163
transform 1 0 12236 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_134
timestamp 1667941163
transform 1 0 13432 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_151
timestamp 1667941163
transform 1 0 14996 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1667941163
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_176
timestamp 1667941163
transform 1 0 17296 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_189
timestamp 1667941163
transform 1 0 18492 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_202
timestamp 1667941163
transform 1 0 19688 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_215
timestamp 1667941163
transform 1 0 20884 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1667941163
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_236
timestamp 1667941163
transform 1 0 22816 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_240
timestamp 1667941163
transform 1 0 23184 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_250
timestamp 1667941163
transform 1 0 24104 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_267
timestamp 1667941163
transform 1 0 25668 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_274
timestamp 1667941163
transform 1 0 26312 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_286
timestamp 1667941163
transform 1 0 27416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_300
timestamp 1667941163
transform 1 0 28704 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_306
timestamp 1667941163
transform 1 0 29256 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_312
timestamp 1667941163
transform 1 0 29808 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_324
timestamp 1667941163
transform 1 0 30912 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_397
timestamp 1667941163
transform 1 0 37628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_59
timestamp 1667941163
transform 1 0 6532 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_62
timestamp 1667941163
transform 1 0 6808 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_68
timestamp 1667941163
transform 1 0 7360 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_75
timestamp 1667941163
transform 1 0 8004 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1667941163
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_91
timestamp 1667941163
transform 1 0 9476 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_98
timestamp 1667941163
transform 1 0 10120 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_105
timestamp 1667941163
transform 1 0 10764 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_112
timestamp 1667941163
transform 1 0 11408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_125
timestamp 1667941163
transform 1 0 12604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1667941163
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_145
timestamp 1667941163
transform 1 0 14444 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_155
timestamp 1667941163
transform 1 0 15364 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_172
timestamp 1667941163
transform 1 0 16928 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_181
timestamp 1667941163
transform 1 0 17756 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1667941163
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1667941163
transform 1 0 19688 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_219
timestamp 1667941163
transform 1 0 21252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_231
timestamp 1667941163
transform 1 0 22356 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_237
timestamp 1667941163
transform 1 0 22908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1667941163
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_264
timestamp 1667941163
transform 1 0 25392 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_277
timestamp 1667941163
transform 1 0 26588 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_284
timestamp 1667941163
transform 1 0 27232 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_291
timestamp 1667941163
transform 1 0 27876 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_298
timestamp 1667941163
transform 1 0 28520 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_305
timestamp 1667941163
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_313
timestamp 1667941163
transform 1 0 29900 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_319
timestamp 1667941163
transform 1 0 30452 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_331
timestamp 1667941163
transform 1 0 31556 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_343
timestamp 1667941163
transform 1 0 32660 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_355
timestamp 1667941163
transform 1 0 33764 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1667941163
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_9
timestamp 1667941163
transform 1 0 1932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_21
timestamp 1667941163
transform 1 0 3036 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_33
timestamp 1667941163
transform 1 0 4140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1667941163
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1667941163
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_62
timestamp 1667941163
transform 1 0 6808 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_68
timestamp 1667941163
transform 1 0 7360 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_75
timestamp 1667941163
transform 1 0 8004 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_82
timestamp 1667941163
transform 1 0 8648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_89
timestamp 1667941163
transform 1 0 9292 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_96
timestamp 1667941163
transform 1 0 9936 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_103
timestamp 1667941163
transform 1 0 10580 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1667941163
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_124
timestamp 1667941163
transform 1 0 12512 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_130
timestamp 1667941163
transform 1 0 13064 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_140
timestamp 1667941163
transform 1 0 13984 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp 1667941163
transform 1 0 15180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1667941163
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1667941163
transform 1 0 17480 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_195
timestamp 1667941163
transform 1 0 19044 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_202
timestamp 1667941163
transform 1 0 19688 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_208
timestamp 1667941163
transform 1 0 20240 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1667941163
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_229
timestamp 1667941163
transform 1 0 22172 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_239
timestamp 1667941163
transform 1 0 23092 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_252
timestamp 1667941163
transform 1 0 24288 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_265
timestamp 1667941163
transform 1 0 25484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_272
timestamp 1667941163
transform 1 0 26128 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1667941163
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_286
timestamp 1667941163
transform 1 0 27416 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_300
timestamp 1667941163
transform 1 0 28704 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_306
timestamp 1667941163
transform 1 0 29256 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_312
timestamp 1667941163
transform 1 0 29808 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_318
timestamp 1667941163
transform 1 0 30360 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_324
timestamp 1667941163
transform 1 0 30912 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1667941163
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_61
timestamp 1667941163
transform 1 0 6716 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_64
timestamp 1667941163
transform 1 0 6992 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_70
timestamp 1667941163
transform 1 0 7544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_76
timestamp 1667941163
transform 1 0 8096 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1667941163
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_92
timestamp 1667941163
transform 1 0 9568 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_99
timestamp 1667941163
transform 1 0 10212 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_106
timestamp 1667941163
transform 1 0 10856 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_113
timestamp 1667941163
transform 1 0 11500 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_125
timestamp 1667941163
transform 1 0 12604 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1667941163
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_147
timestamp 1667941163
transform 1 0 14628 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_164
timestamp 1667941163
transform 1 0 16192 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_177
timestamp 1667941163
transform 1 0 17388 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1667941163
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_208
timestamp 1667941163
transform 1 0 20240 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_229
timestamp 1667941163
transform 1 0 22172 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1667941163
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_264
timestamp 1667941163
transform 1 0 25392 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_277
timestamp 1667941163
transform 1 0 26588 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_284
timestamp 1667941163
transform 1 0 27232 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_297
timestamp 1667941163
transform 1 0 28428 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1667941163
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_313
timestamp 1667941163
transform 1 0 29900 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_325
timestamp 1667941163
transform 1 0 31004 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_337
timestamp 1667941163
transform 1 0 32108 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_349
timestamp 1667941163
transform 1 0 33212 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_361
timestamp 1667941163
transform 1 0 34316 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1667941163
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1667941163
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1667941163
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1667941163
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1667941163
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_73
timestamp 1667941163
transform 1 0 7820 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_76
timestamp 1667941163
transform 1 0 8096 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_82
timestamp 1667941163
transform 1 0 8648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_89
timestamp 1667941163
transform 1 0 9292 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_96
timestamp 1667941163
transform 1 0 9936 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_103
timestamp 1667941163
transform 1 0 10580 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1667941163
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_117
timestamp 1667941163
transform 1 0 11868 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_130
timestamp 1667941163
transform 1 0 13064 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_147
timestamp 1667941163
transform 1 0 14628 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_155
timestamp 1667941163
transform 1 0 15364 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1667941163
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_180
timestamp 1667941163
transform 1 0 17664 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_188
timestamp 1667941163
transform 1 0 18400 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_192
timestamp 1667941163
transform 1 0 18768 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_205
timestamp 1667941163
transform 1 0 19964 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_214
timestamp 1667941163
transform 1 0 20792 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1667941163
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_235
timestamp 1667941163
transform 1 0 22724 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_239
timestamp 1667941163
transform 1 0 23092 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_249
timestamp 1667941163
transform 1 0 24012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_256
timestamp 1667941163
transform 1 0 24656 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_264
timestamp 1667941163
transform 1 0 25392 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_274
timestamp 1667941163
transform 1 0 26312 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_286
timestamp 1667941163
transform 1 0 27416 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_300
timestamp 1667941163
transform 1 0 28704 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_307
timestamp 1667941163
transform 1 0 29348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_313
timestamp 1667941163
transform 1 0 29900 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_319
timestamp 1667941163
transform 1 0 30452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_331
timestamp 1667941163
transform 1 0 31556 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_397
timestamp 1667941163
transform 1 0 37628 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_9
timestamp 1667941163
transform 1 0 1932 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1667941163
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1667941163
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1667941163
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_90
timestamp 1667941163
transform 1 0 9384 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_97
timestamp 1667941163
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_104
timestamp 1667941163
transform 1 0 10672 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_111
timestamp 1667941163
transform 1 0 11316 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_118
timestamp 1667941163
transform 1 0 11960 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_125
timestamp 1667941163
transform 1 0 12604 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1667941163
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_148
timestamp 1667941163
transform 1 0 14720 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_161
timestamp 1667941163
transform 1 0 15916 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_168
timestamp 1667941163
transform 1 0 16560 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_181
timestamp 1667941163
transform 1 0 17756 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1667941163
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_204
timestamp 1667941163
transform 1 0 19872 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_217
timestamp 1667941163
transform 1 0 21068 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_234
timestamp 1667941163
transform 1 0 22632 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_247
timestamp 1667941163
transform 1 0 23828 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1667941163
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_257
timestamp 1667941163
transform 1 0 24748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_267
timestamp 1667941163
transform 1 0 25668 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_280
timestamp 1667941163
transform 1 0 26864 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_287
timestamp 1667941163
transform 1 0 27508 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_294
timestamp 1667941163
transform 1 0 28152 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1667941163
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1667941163
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_313
timestamp 1667941163
transform 1 0 29900 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_325
timestamp 1667941163
transform 1 0 31004 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_337
timestamp 1667941163
transform 1 0 32108 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_349
timestamp 1667941163
transform 1 0 33212 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_361
timestamp 1667941163
transform 1 0 34316 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_401
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_84
timestamp 1667941163
transform 1 0 8832 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_90
timestamp 1667941163
transform 1 0 9384 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_96
timestamp 1667941163
transform 1 0 9936 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_103
timestamp 1667941163
transform 1 0 10580 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1667941163
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_119
timestamp 1667941163
transform 1 0 12052 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_123
timestamp 1667941163
transform 1 0 12420 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_136
timestamp 1667941163
transform 1 0 13616 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_149
timestamp 1667941163
transform 1 0 14812 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_162
timestamp 1667941163
transform 1 0 16008 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_184
timestamp 1667941163
transform 1 0 18032 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_197
timestamp 1667941163
transform 1 0 19228 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_204
timestamp 1667941163
transform 1 0 19872 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_211
timestamp 1667941163
transform 1 0 20516 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1667941163
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_240
timestamp 1667941163
transform 1 0 23184 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_246
timestamp 1667941163
transform 1 0 23736 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_259
timestamp 1667941163
transform 1 0 24932 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_272
timestamp 1667941163
transform 1 0 26128 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1667941163
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_286
timestamp 1667941163
transform 1 0 27416 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_300
timestamp 1667941163
transform 1 0 28704 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_306
timestamp 1667941163
transform 1 0 29256 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_312
timestamp 1667941163
transform 1 0 29808 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_324
timestamp 1667941163
transform 1 0 30912 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_65
timestamp 1667941163
transform 1 0 7084 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_73
timestamp 1667941163
transform 1 0 7820 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_78
timestamp 1667941163
transform 1 0 8280 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_95
timestamp 1667941163
transform 1 0 9844 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_102
timestamp 1667941163
transform 1 0 10488 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_108
timestamp 1667941163
transform 1 0 11040 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_112
timestamp 1667941163
transform 1 0 11408 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_119
timestamp 1667941163
transform 1 0 12052 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_126
timestamp 1667941163
transform 1 0 12696 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1667941163
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_152
timestamp 1667941163
transform 1 0 15088 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_158
timestamp 1667941163
transform 1 0 15640 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_168
timestamp 1667941163
transform 1 0 16560 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_181
timestamp 1667941163
transform 1 0 17756 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_187
timestamp 1667941163
transform 1 0 18308 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1667941163
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_203
timestamp 1667941163
transform 1 0 19780 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_210
timestamp 1667941163
transform 1 0 20424 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_223
timestamp 1667941163
transform 1 0 21620 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_234
timestamp 1667941163
transform 1 0 22632 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_247
timestamp 1667941163
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1667941163
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_264
timestamp 1667941163
transform 1 0 25392 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_277
timestamp 1667941163
transform 1 0 26588 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_284
timestamp 1667941163
transform 1 0 27232 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_291
timestamp 1667941163
transform 1 0 27876 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_298
timestamp 1667941163
transform 1 0 28520 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_304
timestamp 1667941163
transform 1 0 29072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_313
timestamp 1667941163
transform 1 0 29900 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_326
timestamp 1667941163
transform 1 0 31096 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_338
timestamp 1667941163
transform 1 0 32200 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_350
timestamp 1667941163
transform 1 0 33304 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1667941163
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1667941163
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1667941163
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1667941163
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1667941163
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_93
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_99
timestamp 1667941163
transform 1 0 10212 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_107
timestamp 1667941163
transform 1 0 10948 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1667941163
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1667941163
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_123
timestamp 1667941163
transform 1 0 12420 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_136
timestamp 1667941163
transform 1 0 13616 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_149
timestamp 1667941163
transform 1 0 14812 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1667941163
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_180
timestamp 1667941163
transform 1 0 17664 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_189
timestamp 1667941163
transform 1 0 18492 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_204
timestamp 1667941163
transform 1 0 19872 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_208
timestamp 1667941163
transform 1 0 20240 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_218
timestamp 1667941163
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_231
timestamp 1667941163
transform 1 0 22356 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_239
timestamp 1667941163
transform 1 0 23092 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_249
timestamp 1667941163
transform 1 0 24012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_257
timestamp 1667941163
transform 1 0 24748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_270
timestamp 1667941163
transform 1 0 25944 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_277
timestamp 1667941163
transform 1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_286
timestamp 1667941163
transform 1 0 27416 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_293
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_300
timestamp 1667941163
transform 1 0 28704 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_306
timestamp 1667941163
transform 1 0 29256 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_318
timestamp 1667941163
transform 1 0 30360 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_330
timestamp 1667941163
transform 1 0 31464 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1667941163
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_397
timestamp 1667941163
transform 1 0 37628 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1667941163
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1667941163
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_109
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_114
timestamp 1667941163
transform 1 0 11592 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_124
timestamp 1667941163
transform 1 0 12512 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_131
timestamp 1667941163
transform 1 0 13156 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1667941163
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_152
timestamp 1667941163
transform 1 0 15088 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1667941163
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_170
timestamp 1667941163
transform 1 0 16744 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_177
timestamp 1667941163
transform 1 0 17388 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1667941163
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_203
timestamp 1667941163
transform 1 0 19780 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_216
timestamp 1667941163
transform 1 0 20976 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_223
timestamp 1667941163
transform 1 0 21620 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_238
timestamp 1667941163
transform 1 0 23000 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1667941163
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1667941163
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_264
timestamp 1667941163
transform 1 0 25392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_277
timestamp 1667941163
transform 1 0 26588 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_284
timestamp 1667941163
transform 1 0 27232 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_291
timestamp 1667941163
transform 1 0 27876 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_297
timestamp 1667941163
transform 1 0 28428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_303
timestamp 1667941163
transform 1 0 28980 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1667941163
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1667941163
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1667941163
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1667941163
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1667941163
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1667941163
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1667941163
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_125
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_133
timestamp 1667941163
transform 1 0 13340 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_139
timestamp 1667941163
transform 1 0 13892 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_146
timestamp 1667941163
transform 1 0 14536 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_153
timestamp 1667941163
transform 1 0 15180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1667941163
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_180
timestamp 1667941163
transform 1 0 17664 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_186
timestamp 1667941163
transform 1 0 18216 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_193
timestamp 1667941163
transform 1 0 18860 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_206
timestamp 1667941163
transform 1 0 20056 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_214
timestamp 1667941163
transform 1 0 20792 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_218
timestamp 1667941163
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_231
timestamp 1667941163
transform 1 0 22356 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_237
timestamp 1667941163
transform 1 0 22908 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_250
timestamp 1667941163
transform 1 0 24104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_257
timestamp 1667941163
transform 1 0 24748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_261
timestamp 1667941163
transform 1 0 25116 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_271
timestamp 1667941163
transform 1 0 26036 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1667941163
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_285
timestamp 1667941163
transform 1 0 27324 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_297
timestamp 1667941163
transform 1 0 28428 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_309
timestamp 1667941163
transform 1 0 29532 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_321
timestamp 1667941163
transform 1 0 30636 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_333
timestamp 1667941163
transform 1 0 31740 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_397
timestamp 1667941163
transform 1 0 37628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_7
timestamp 1667941163
transform 1 0 1748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1667941163
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1667941163
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1667941163
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1667941163
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1667941163
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1667941163
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1667941163
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_146
timestamp 1667941163
transform 1 0 14536 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_152
timestamp 1667941163
transform 1 0 15088 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_159
timestamp 1667941163
transform 1 0 15732 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_170
timestamp 1667941163
transform 1 0 16744 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_177
timestamp 1667941163
transform 1 0 17388 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_183
timestamp 1667941163
transform 1 0 17940 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_190
timestamp 1667941163
transform 1 0 18584 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_203
timestamp 1667941163
transform 1 0 19780 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_216
timestamp 1667941163
transform 1 0 20976 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_223
timestamp 1667941163
transform 1 0 21620 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_229
timestamp 1667941163
transform 1 0 22172 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_233
timestamp 1667941163
transform 1 0 22540 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_246
timestamp 1667941163
transform 1 0 23736 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_264
timestamp 1667941163
transform 1 0 25392 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_271
timestamp 1667941163
transform 1 0 26036 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_277
timestamp 1667941163
transform 1 0 26588 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_283
timestamp 1667941163
transform 1 0 27140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_295
timestamp 1667941163
transform 1 0 28244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1667941163
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1667941163
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1667941163
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_9
timestamp 1667941163
transform 1 0 1932 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_21
timestamp 1667941163
transform 1 0 3036 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_33
timestamp 1667941163
transform 1 0 4140 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_37
timestamp 1667941163
transform 1 0 4508 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_41
timestamp 1667941163
transform 1 0 4876 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_47
timestamp 1667941163
transform 1 0 5428 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1667941163
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1667941163
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1667941163
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1667941163
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_149
timestamp 1667941163
transform 1 0 14812 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_159
timestamp 1667941163
transform 1 0 15732 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1667941163
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1667941163
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_184
timestamp 1667941163
transform 1 0 18032 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_187
timestamp 1667941163
transform 1 0 18308 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_200
timestamp 1667941163
transform 1 0 19504 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_213
timestamp 1667941163
transform 1 0 20700 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1667941163
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_236
timestamp 1667941163
transform 1 0 22816 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_242
timestamp 1667941163
transform 1 0 23368 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_249
timestamp 1667941163
transform 1 0 24012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_256
timestamp 1667941163
transform 1 0 24656 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_263
timestamp 1667941163
transform 1 0 25300 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_269
timestamp 1667941163
transform 1 0 25852 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_277
timestamp 1667941163
transform 1 0 26588 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1667941163
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1667941163
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1667941163
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1667941163
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1667941163
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1667941163
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1667941163
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1667941163
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1667941163
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1667941163
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1667941163
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_153
timestamp 1667941163
transform 1 0 15180 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_161
timestamp 1667941163
transform 1 0 15916 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_165
timestamp 1667941163
transform 1 0 16284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_169
timestamp 1667941163
transform 1 0 16652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_172
timestamp 1667941163
transform 1 0 16928 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_176
timestamp 1667941163
transform 1 0 17296 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_179
timestamp 1667941163
transform 1 0 17572 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_185
timestamp 1667941163
transform 1 0 18124 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_188
timestamp 1667941163
transform 1 0 18400 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1667941163
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_212
timestamp 1667941163
transform 1 0 20608 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_219
timestamp 1667941163
transform 1 0 21252 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_227
timestamp 1667941163
transform 1 0 21988 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_231
timestamp 1667941163
transform 1 0 22356 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_237
timestamp 1667941163
transform 1 0 22908 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_246
timestamp 1667941163
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_257
timestamp 1667941163
transform 1 0 24748 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_263
timestamp 1667941163
transform 1 0 25300 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_275
timestamp 1667941163
transform 1 0 26404 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_287
timestamp 1667941163
transform 1 0 27508 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_299
timestamp 1667941163
transform 1 0 28612 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1667941163
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1667941163
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_12
timestamp 1667941163
transform 1 0 2208 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_18
timestamp 1667941163
transform 1 0 2760 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_30
timestamp 1667941163
transform 1 0 3864 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_42
timestamp 1667941163
transform 1 0 4968 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1667941163
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_96
timestamp 1667941163
transform 1 0 9936 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1667941163
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_117
timestamp 1667941163
transform 1 0 11868 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_120
timestamp 1667941163
transform 1 0 12144 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_128
timestamp 1667941163
transform 1 0 12880 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_140
timestamp 1667941163
transform 1 0 13984 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_152
timestamp 1667941163
transform 1 0 15088 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1667941163
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1667941163
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_193
timestamp 1667941163
transform 1 0 18860 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_197
timestamp 1667941163
transform 1 0 19228 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_204
timestamp 1667941163
transform 1 0 19872 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_211
timestamp 1667941163
transform 1 0 20516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1667941163
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1667941163
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_229
timestamp 1667941163
transform 1 0 22172 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_237
timestamp 1667941163
transform 1 0 22908 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_240
timestamp 1667941163
transform 1 0 23184 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_246
timestamp 1667941163
transform 1 0 23736 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_258
timestamp 1667941163
transform 1 0 24840 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_270
timestamp 1667941163
transform 1 0 25944 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1667941163
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1667941163
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1667941163
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1667941163
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1667941163
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_9
timestamp 1667941163
transform 1 0 1932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_16
timestamp 1667941163
transform 1 0 2576 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_22
timestamp 1667941163
transform 1 0 3128 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1667941163
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1667941163
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1667941163
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1667941163
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1667941163
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1667941163
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1667941163
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1667941163
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_177
timestamp 1667941163
transform 1 0 17388 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_187
timestamp 1667941163
transform 1 0 18308 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1667941163
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_202
timestamp 1667941163
transform 1 0 19688 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_209
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_215
timestamp 1667941163
transform 1 0 20884 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_227
timestamp 1667941163
transform 1 0 21988 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_235
timestamp 1667941163
transform 1 0 22724 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_241
timestamp 1667941163
transform 1 0 23276 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_247
timestamp 1667941163
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1667941163
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1667941163
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1667941163
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1667941163
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1667941163
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1667941163
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1667941163
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1667941163
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1667941163
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1667941163
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1667941163
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1667941163
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1667941163
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1667941163
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1667941163
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_181
timestamp 1667941163
transform 1 0 17756 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_189
timestamp 1667941163
transform 1 0 18492 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_201
timestamp 1667941163
transform 1 0 19596 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_207
timestamp 1667941163
transform 1 0 20148 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_219
timestamp 1667941163
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1667941163
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1667941163
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1667941163
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1667941163
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1667941163
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1667941163
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1667941163
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_10
timestamp 1667941163
transform 1 0 2024 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_22
timestamp 1667941163
transform 1 0 3128 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1667941163
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1667941163
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1667941163
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1667941163
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1667941163
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1667941163
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1667941163
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1667941163
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1667941163
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1667941163
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1667941163
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_202
timestamp 1667941163
transform 1 0 19688 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_214
timestamp 1667941163
transform 1 0 20792 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_226
timestamp 1667941163
transform 1 0 21896 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_238
timestamp 1667941163
transform 1 0 23000 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1667941163
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1667941163
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1667941163
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1667941163
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1667941163
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_9
timestamp 1667941163
transform 1 0 1932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_21
timestamp 1667941163
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_33
timestamp 1667941163
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_45
timestamp 1667941163
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1667941163
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_62
timestamp 1667941163
transform 1 0 6808 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_68
timestamp 1667941163
transform 1 0 7360 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_80
timestamp 1667941163
transform 1 0 8464 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_92
timestamp 1667941163
transform 1 0 9568 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_104
timestamp 1667941163
transform 1 0 10672 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1667941163
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1667941163
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1667941163
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1667941163
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_193
timestamp 1667941163
transform 1 0 18860 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_201
timestamp 1667941163
transform 1 0 19596 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_206
timestamp 1667941163
transform 1 0 20056 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_212
timestamp 1667941163
transform 1 0 20608 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1667941163
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1667941163
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_261
timestamp 1667941163
transform 1 0 25116 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_270
timestamp 1667941163
transform 1 0 25944 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1667941163
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1667941163
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_397
timestamp 1667941163
transform 1 0 37628 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1667941163
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1667941163
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1667941163
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1667941163
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1667941163
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1667941163
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1667941163
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1667941163
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1667941163
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1667941163
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1667941163
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1667941163
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1667941163
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1667941163
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1667941163
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1667941163
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1667941163
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_401
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1667941163
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1667941163
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1667941163
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1667941163
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1667941163
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1667941163
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1667941163
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1667941163
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_137
timestamp 1667941163
transform 1 0 13708 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_145
timestamp 1667941163
transform 1 0 14444 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_150
timestamp 1667941163
transform 1 0 14904 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_156
timestamp 1667941163
transform 1 0 15456 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1667941163
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1667941163
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1667941163
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1667941163
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1667941163
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1667941163
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1667941163
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1667941163
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1667941163
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1667941163
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1667941163
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_397
timestamp 1667941163
transform 1 0 37628 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1667941163
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1667941163
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1667941163
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1667941163
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1667941163
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1667941163
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1667941163
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1667941163
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1667941163
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1667941163
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1667941163
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1667941163
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1667941163
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1667941163
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1667941163
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1667941163
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_9
timestamp 1667941163
transform 1 0 1932 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_21
timestamp 1667941163
transform 1 0 3036 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_33
timestamp 1667941163
transform 1 0 4140 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_45
timestamp 1667941163
transform 1 0 5244 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_53
timestamp 1667941163
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1667941163
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1667941163
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1667941163
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1667941163
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1667941163
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1667941163
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1667941163
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1667941163
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1667941163
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1667941163
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1667941163
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1667941163
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1667941163
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1667941163
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1667941163
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1667941163
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1667941163
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1667941163
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1667941163
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1667941163
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1667941163
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1667941163
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1667941163
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1667941163
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1667941163
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1667941163
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1667941163
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1667941163
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1667941163
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1667941163
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1667941163
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1667941163
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1667941163
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_317
timestamp 1667941163
transform 1 0 30268 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_323
timestamp 1667941163
transform 1 0 30820 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_329
timestamp 1667941163
transform 1 0 31372 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_341
timestamp 1667941163
transform 1 0 32476 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_353
timestamp 1667941163
transform 1 0 33580 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_361
timestamp 1667941163
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_401
timestamp 1667941163
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_7
timestamp 1667941163
transform 1 0 1748 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_19
timestamp 1667941163
transform 1 0 2852 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_31
timestamp 1667941163
transform 1 0 3956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_43
timestamp 1667941163
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1667941163
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1667941163
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1667941163
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1667941163
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1667941163
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1667941163
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1667941163
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1667941163
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1667941163
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1667941163
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1667941163
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1667941163
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1667941163
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1667941163
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1667941163
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1667941163
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1667941163
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1667941163
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_397
timestamp 1667941163
transform 1 0 37628 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1667941163
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_121
timestamp 1667941163
transform 1 0 12236 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_131
timestamp 1667941163
transform 1 0 13156 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1667941163
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_153
timestamp 1667941163
transform 1 0 15180 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_161
timestamp 1667941163
transform 1 0 15916 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_166
timestamp 1667941163
transform 1 0 16376 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_172
timestamp 1667941163
transform 1 0 16928 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_184
timestamp 1667941163
transform 1 0 18032 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1667941163
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1667941163
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1667941163
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1667941163
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1667941163
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_292
timestamp 1667941163
transform 1 0 27968 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_298
timestamp 1667941163
transform 1 0 28520 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 1667941163
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1667941163
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1667941163
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1667941163
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_401
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1667941163
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1667941163
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1667941163
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1667941163
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1667941163
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1667941163
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_196
timestamp 1667941163
transform 1 0 19136 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_202
timestamp 1667941163
transform 1 0 19688 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_214
timestamp 1667941163
transform 1 0 20792 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1667941163
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1667941163
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1667941163
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1667941163
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1667941163
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1667941163
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1667941163
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1667941163
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1667941163
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_153
timestamp 1667941163
transform 1 0 15180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_157
timestamp 1667941163
transform 1 0 15548 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_160
timestamp 1667941163
transform 1 0 15824 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_168
timestamp 1667941163
transform 1 0 16560 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_180
timestamp 1667941163
transform 1 0 17664 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1667941163
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1667941163
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1667941163
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1667941163
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1667941163
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1667941163
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1667941163
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1667941163
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1667941163
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_401
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_405
timestamp 1667941163
transform 1 0 38364 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_9
timestamp 1667941163
transform 1 0 1932 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_21
timestamp 1667941163
transform 1 0 3036 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_33
timestamp 1667941163
transform 1 0 4140 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_45
timestamp 1667941163
transform 1 0 5244 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1667941163
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1667941163
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1667941163
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1667941163
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1667941163
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1667941163
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1667941163
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1667941163
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1667941163
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1667941163
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1667941163
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1667941163
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_232
timestamp 1667941163
transform 1 0 22448 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_238
timestamp 1667941163
transform 1 0 23000 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_250
timestamp 1667941163
transform 1 0 24104 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_262
timestamp 1667941163
transform 1 0 25208 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_274
timestamp 1667941163
transform 1 0 26312 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_322
timestamp 1667941163
transform 1 0 30728 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_334
timestamp 1667941163
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1667941163
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1667941163
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1667941163
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1667941163
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1667941163
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1667941163
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1667941163
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1667941163
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1667941163
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1667941163
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1667941163
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1667941163
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1667941163
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1667941163
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1667941163
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1667941163
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_137
timestamp 1667941163
transform 1 0 13708 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_143
timestamp 1667941163
transform 1 0 14260 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_147
timestamp 1667941163
transform 1 0 14628 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_153
timestamp 1667941163
transform 1 0 15180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_165
timestamp 1667941163
transform 1 0 16284 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1667941163
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1667941163
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1667941163
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1667941163
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1667941163
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1667941163
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1667941163
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1667941163
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1667941163
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_397
timestamp 1667941163
transform 1 0 37628 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_7
timestamp 1667941163
transform 1 0 1748 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_19
timestamp 1667941163
transform 1 0 2852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1667941163
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_121
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_129
timestamp 1667941163
transform 1 0 12972 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_135
timestamp 1667941163
transform 1 0 13524 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1667941163
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1667941163
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1667941163
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_221
timestamp 1667941163
transform 1 0 21436 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_226
timestamp 1667941163
transform 1 0 21896 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_232
timestamp 1667941163
transform 1 0 22448 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_244
timestamp 1667941163
transform 1 0 23552 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1667941163
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1667941163
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1667941163
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1667941163
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1667941163
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1667941163
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1667941163
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1667941163
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1667941163
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1667941163
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_212
timestamp 1667941163
transform 1 0 20608 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_401
timestamp 1667941163
transform 1 0 37996 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_404
timestamp 1667941163
transform 1 0 38272 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1667941163
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1667941163
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1667941163
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1667941163
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1667941163
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1667941163
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1667941163
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1667941163
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1667941163
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1667941163
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1667941163
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_397
timestamp 1667941163
transform 1 0 37628 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_402
timestamp 1667941163
transform 1 0 38088 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_406
timestamp 1667941163
transform 1 0 38456 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_7
timestamp 1667941163
transform 1 0 1748 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_19
timestamp 1667941163
transform 1 0 2852 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_31
timestamp 1667941163
transform 1 0 3956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_43
timestamp 1667941163
transform 1 0 5060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1667941163
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1667941163
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1667941163
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_137
timestamp 1667941163
transform 1 0 13708 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_145
timestamp 1667941163
transform 1 0 14444 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_150
timestamp 1667941163
transform 1 0 14904 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_158
timestamp 1667941163
transform 1 0 15640 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1667941163
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1667941163
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1667941163
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1667941163
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1667941163
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1667941163
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1667941163
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1667941163
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1667941163
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_9
timestamp 1667941163
transform 1 0 1932 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1667941163
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1667941163
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1667941163
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1667941163
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1667941163
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1667941163
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1667941163
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1667941163
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1667941163
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_283
timestamp 1667941163
transform 1 0 27140 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_287
timestamp 1667941163
transform 1 0 27508 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_293
timestamp 1667941163
transform 1 0 28060 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_305
timestamp 1667941163
transform 1 0 29164 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_325
timestamp 1667941163
transform 1 0 31004 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_331
timestamp 1667941163
transform 1 0 31556 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_343
timestamp 1667941163
transform 1 0 32660 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_355
timestamp 1667941163
transform 1 0 33764 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1667941163
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1667941163
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1667941163
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1667941163
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1667941163
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1667941163
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_7
timestamp 1667941163
transform 1 0 1748 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_19
timestamp 1667941163
transform 1 0 2852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1667941163
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1667941163
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1667941163
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1667941163
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1667941163
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_405
timestamp 1667941163
transform 1 0 38364 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_9
timestamp 1667941163
transform 1 0 1932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_21
timestamp 1667941163
transform 1 0 3036 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_33
timestamp 1667941163
transform 1 0 4140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1667941163
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1667941163
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1667941163
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1667941163
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1667941163
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1667941163
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1667941163
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_397
timestamp 1667941163
transform 1 0 37628 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_61
timestamp 1667941163
transform 1 0 6716 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_66
timestamp 1667941163
transform 1 0 7176 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_72
timestamp 1667941163
transform 1 0 7728 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_9
timestamp 1667941163
transform 1 0 1932 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1667941163
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1667941163
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1667941163
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1667941163
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1667941163
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_205
timestamp 1667941163
transform 1 0 19964 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_215
timestamp 1667941163
transform 1 0 20884 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_227
timestamp 1667941163
transform 1 0 21988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_239
timestamp 1667941163
transform 1 0 23092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_314
timestamp 1667941163
transform 1 0 29992 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_320
timestamp 1667941163
transform 1 0 30544 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_332
timestamp 1667941163
transform 1 0 31648 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_344
timestamp 1667941163
transform 1 0 32752 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_356
timestamp 1667941163
transform 1 0 33856 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_401
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_405
timestamp 1667941163
transform 1 0 38364 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_9
timestamp 1667941163
transform 1 0 1932 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_13
timestamp 1667941163
transform 1 0 2300 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_19
timestamp 1667941163
transform 1 0 2852 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_31
timestamp 1667941163
transform 1 0 3956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_43
timestamp 1667941163
transform 1 0 5060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1667941163
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_9
timestamp 1667941163
transform 1 0 1932 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1667941163
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1667941163
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_385
timestamp 1667941163
transform 1 0 36524 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_397
timestamp 1667941163
transform 1 0 37628 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_17
timestamp 1667941163
transform 1 0 2668 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_23
timestamp 1667941163
transform 1 0 3220 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_35
timestamp 1667941163
transform 1 0 4324 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_47
timestamp 1667941163
transform 1 0 5428 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1667941163
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_93
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_104
timestamp 1667941163
transform 1 0 10672 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1667941163
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1667941163
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1667941163
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1667941163
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1667941163
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1667941163
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1667941163
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_230
timestamp 1667941163
transform 1 0 22264 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_236
timestamp 1667941163
transform 1 0 22816 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_248
timestamp 1667941163
transform 1 0 23920 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_260
timestamp 1667941163
transform 1 0 25024 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_272
timestamp 1667941163
transform 1 0 26128 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_289
timestamp 1667941163
transform 1 0 27692 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1667941163
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1667941163
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1667941163
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1667941163
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1667941163
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1667941163
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_385
timestamp 1667941163
transform 1 0 36524 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1667941163
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_399
timestamp 1667941163
transform 1 0 37812 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_9
timestamp 1667941163
transform 1 0 1932 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_21
timestamp 1667941163
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1667941163
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_37
timestamp 1667941163
transform 1 0 4508 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_42
timestamp 1667941163
transform 1 0 4968 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_48
timestamp 1667941163
transform 1 0 5520 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_63
timestamp 1667941163
transform 1 0 6900 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_69
timestamp 1667941163
transform 1 0 7452 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1667941163
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1667941163
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_93
timestamp 1667941163
transform 1 0 9660 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_98
timestamp 1667941163
transform 1 0 10120 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_110
timestamp 1667941163
transform 1 0 11224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_119
timestamp 1667941163
transform 1 0 12052 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_125
timestamp 1667941163
transform 1 0 12604 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1667941163
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1667941163
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_146
timestamp 1667941163
transform 1 0 14536 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_160
timestamp 1667941163
transform 1 0 15824 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_166
timestamp 1667941163
transform 1 0 16376 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_175
timestamp 1667941163
transform 1 0 17204 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_181
timestamp 1667941163
transform 1 0 17756 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1667941163
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1667941163
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_205
timestamp 1667941163
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_210
timestamp 1667941163
transform 1 0 20424 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_218
timestamp 1667941163
transform 1 0 21160 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1667941163
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_237
timestamp 1667941163
transform 1 0 22908 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1667941163
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1667941163
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_261
timestamp 1667941163
transform 1 0 25116 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_266
timestamp 1667941163
transform 1 0 25576 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_278
timestamp 1667941163
transform 1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_287
timestamp 1667941163
transform 1 0 27508 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_295
timestamp 1667941163
transform 1 0 28244 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1667941163
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1667941163
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_317
timestamp 1667941163
transform 1 0 30268 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_322
timestamp 1667941163
transform 1 0 30728 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_334
timestamp 1667941163
transform 1 0 31832 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_343
timestamp 1667941163
transform 1 0 32660 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_351
timestamp 1667941163
transform 1 0 33396 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1667941163
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1667941163
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_370
timestamp 1667941163
transform 1 0 35144 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_384
timestamp 1667941163
transform 1 0 36432 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_390
timestamp 1667941163
transform 1 0 36984 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1667941163
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _216_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 10580 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1667941163
transform -1 0 26680 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1667941163
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1667941163
transform 1 0 25024 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1667941163
transform -1 0 17388 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _221_
timestamp 1667941163
transform 1 0 22264 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1667941163
transform -1 0 19688 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _223_
timestamp 1667941163
transform 1 0 14904 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _224_
timestamp 1667941163
transform -1 0 12604 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1667941163
transform -1 0 28060 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1667941163
transform 1 0 16100 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1667941163
transform -1 0 24656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1667941163
transform 1 0 26956 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1667941163
transform -1 0 27508 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp 1667941163
transform 1 0 22356 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp 1667941163
transform -1 0 27232 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _232_
timestamp 1667941163
transform -1 0 20700 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _233_
timestamp 1667941163
transform -1 0 20516 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _234_
timestamp 1667941163
transform -1 0 20424 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1667941163
transform -1 0 16100 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1667941163
transform 1 0 10948 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 1667941163
transform 1 0 14444 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 1667941163
transform 1 0 28428 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 1667941163
transform 1 0 18584 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1667941163
transform 1 0 9292 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1667941163
transform 1 0 27784 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 1667941163
transform 1 0 20792 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 1667941163
transform -1 0 18768 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1667941163
transform 1 0 9936 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 1667941163
transform -1 0 19688 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 1667941163
transform -1 0 21344 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1667941163
transform 1 0 24380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1667941163
transform -1 0 17112 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 1667941163
transform 1 0 26036 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1667941163
transform 1 0 9844 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 1667941163
transform 1 0 27600 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 1667941163
transform -1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1667941163
transform 1 0 17112 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1667941163
transform 1 0 18308 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1667941163
transform 1 0 19412 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1667941163
transform -1 0 28704 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1667941163
transform -1 0 14536 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 1667941163
transform -1 0 16744 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1667941163
transform -1 0 9936 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1667941163
transform -1 0 28060 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1667941163
transform -1 0 13800 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1667941163
transform -1 0 27876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1667941163
transform -1 0 18400 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1667941163
transform -1 0 11224 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1667941163
transform -1 0 26312 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1667941163
transform 1 0 10948 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1667941163
transform -1 0 28060 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1667941163
transform -1 0 12052 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1667941163
transform 1 0 9200 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1667941163
transform -1 0 10672 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1667941163
transform -1 0 27416 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1667941163
transform -1 0 10580 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1667941163
transform 1 0 9016 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1667941163
transform 1 0 11776 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1667941163
transform 1 0 10304 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1667941163
transform -1 0 11408 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1667941163
transform 1 0 23736 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _278_
timestamp 1667941163
transform 1 0 24288 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1667941163
transform -1 0 16744 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1667941163
transform -1 0 13432 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _281_
timestamp 1667941163
transform 1 0 19504 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1667941163
transform 1 0 8372 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1667941163
transform -1 0 11040 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp 1667941163
transform -1 0 10580 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1667941163
transform -1 0 27416 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1667941163
transform 1 0 11040 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _287_
timestamp 1667941163
transform 1 0 13524 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _288_
timestamp 1667941163
transform -1 0 24104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _289_
timestamp 1667941163
transform 1 0 26312 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _290_
timestamp 1667941163
transform -1 0 26036 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _291_
timestamp 1667941163
transform -1 0 28520 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1667941163
transform 1 0 24840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _293_
timestamp 1667941163
transform -1 0 23736 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1667941163
transform -1 0 24748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1667941163
transform 1 0 12144 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 1667941163
transform 1 0 24564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 1667941163
transform -1 0 21344 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1667941163
transform -1 0 21160 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1667941163
transform -1 0 28152 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 1667941163
transform 1 0 20148 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1667941163
transform -1 0 27416 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 1667941163
transform -1 0 28060 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _303_
timestamp 1667941163
transform 1 0 27140 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1667941163
transform 1 0 17480 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1667941163
transform -1 0 22356 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _306_
timestamp 1667941163
transform 1 0 19596 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1667941163
transform -1 0 18492 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1667941163
transform 1 0 20608 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1667941163
transform 1 0 27600 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 1667941163
transform -1 0 28704 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 1667941163
transform -1 0 21620 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 1667941163
transform -1 0 11408 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1667941163
transform -1 0 21528 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1667941163
transform 1 0 20516 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1667941163
transform -1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1667941163
transform -1 0 11224 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 1667941163
transform -1 0 26128 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _318_
timestamp 1667941163
transform -1 0 21620 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 1667941163
transform 1 0 21252 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1667941163
transform -1 0 10764 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1667941163
transform 1 0 28520 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 1667941163
transform -1 0 15732 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1667941163
transform 1 0 27784 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1667941163
transform 1 0 24748 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 1667941163
transform 1 0 19596 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1667941163
transform 1 0 17480 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1667941163
transform -1 0 28520 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1667941163
transform 1 0 28060 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 1667941163
transform 1 0 19412 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp 1667941163
transform 1 0 17020 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp 1667941163
transform -1 0 28428 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1667941163
transform 1 0 27600 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1667941163
transform 1 0 10396 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1667941163
transform 1 0 10948 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1667941163
transform -1 0 11316 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp 1667941163
transform -1 0 13432 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp 1667941163
transform 1 0 16284 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp 1667941163
transform -1 0 12788 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1667941163
transform -1 0 8648 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1667941163
transform -1 0 10580 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp 1667941163
transform 1 0 9752 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1667941163
transform 1 0 21252 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp 1667941163
transform 1 0 9108 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp 1667941163
transform -1 0 10580 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1667941163
transform -1 0 13156 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1667941163
transform 1 0 11224 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1667941163
transform 1 0 12420 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1667941163
transform 1 0 11132 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1667941163
transform -1 0 13800 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1667941163
transform 1 0 11408 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp 1667941163
transform -1 0 2944 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _352_
timestamp 1667941163
transform -1 0 28336 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp 1667941163
transform -1 0 19872 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1667941163
transform -1 0 19688 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1667941163
transform -1 0 14904 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1667941163
transform 1 0 9016 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp 1667941163
transform 1 0 30728 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1667941163
transform -1 0 26404 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1667941163
transform -1 0 27416 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _360_
timestamp 1667941163
transform 1 0 9752 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _361_
timestamp 1667941163
transform -1 0 27232 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _362_
timestamp 1667941163
transform -1 0 24840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1667941163
transform 1 0 7728 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _364_
timestamp 1667941163
transform -1 0 7176 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1667941163
transform 1 0 8372 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _367_
timestamp 1667941163
transform -1 0 23276 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1667941163
transform -1 0 28704 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1667941163
transform -1 0 27416 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1667941163
transform -1 0 30820 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1667941163
transform -1 0 14628 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1667941163
transform 1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _373_
timestamp 1667941163
transform -1 0 26312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _374_
timestamp 1667941163
transform -1 0 20332 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp 1667941163
transform -1 0 29348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _376_
timestamp 1667941163
transform -1 0 30728 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp 1667941163
transform 1 0 12144 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _378_
timestamp 1667941163
transform 1 0 30360 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _379_
timestamp 1667941163
transform -1 0 21896 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _380_
timestamp 1667941163
transform 1 0 16100 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _381_
timestamp 1667941163
transform -1 0 27232 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _382_
timestamp 1667941163
transform -1 0 20516 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _383_
timestamp 1667941163
transform -1 0 27968 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _384_
timestamp 1667941163
transform 1 0 10212 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _385_
timestamp 1667941163
transform -1 0 8004 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _386_
timestamp 1667941163
transform -1 0 20608 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _387_
timestamp 1667941163
transform 1 0 9660 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp 1667941163
transform 1 0 13248 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _389_
timestamp 1667941163
transform -1 0 17480 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _390_
timestamp 1667941163
transform -1 0 25668 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _391_
timestamp 1667941163
transform 1 0 11684 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _392_
timestamp 1667941163
transform -1 0 2300 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _393_
timestamp 1667941163
transform 1 0 30820 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _394_
timestamp 1667941163
transform -1 0 11592 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _395_
timestamp 1667941163
transform 1 0 9292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _396_
timestamp 1667941163
transform -1 0 8280 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _397_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 33028 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _398_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 30268 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _399_
timestamp 1667941163
transform -1 0 31372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _400_
timestamp 1667941163
transform -1 0 30636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _401_
timestamp 1667941163
transform -1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _402_
timestamp 1667941163
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _403_
timestamp 1667941163
transform -1 0 26312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _404_
timestamp 1667941163
transform 1 0 34224 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _405_
timestamp 1667941163
transform -1 0 30728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _406_
timestamp 1667941163
transform -1 0 29992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _407_
timestamp 1667941163
transform -1 0 27508 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _408_
timestamp 1667941163
transform -1 0 26956 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _409_
timestamp 1667941163
transform -1 0 28980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _410_
timestamp 1667941163
transform 1 0 29072 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _411_
timestamp 1667941163
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _412_
timestamp 1667941163
transform -1 0 28060 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _413_
timestamp 1667941163
transform -1 0 27692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _414_
timestamp 1667941163
transform -1 0 26864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _415_
timestamp 1667941163
transform -1 0 28244 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _416_
timestamp 1667941163
transform -1 0 28060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _417_
timestamp 1667941163
transform -1 0 28060 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _418_
timestamp 1667941163
transform -1 0 28980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _419_
timestamp 1667941163
transform 1 0 29164 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _420_
timestamp 1667941163
transform -1 0 30268 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _421_
timestamp 1667941163
transform -1 0 28152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _422_
timestamp 1667941163
transform -1 0 28704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _423_
timestamp 1667941163
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _424_
timestamp 1667941163
transform -1 0 27416 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _425_
timestamp 1667941163
transform -1 0 29624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _426_
timestamp 1667941163
transform -1 0 28980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _427_
timestamp 1667941163
transform -1 0 29992 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _428_
timestamp 1667941163
transform -1 0 27600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _429_
timestamp 1667941163
transform -1 0 28980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 1667941163
transform -1 0 26864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _431_
timestamp 1667941163
transform -1 0 29072 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 1667941163
transform 1 0 29808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _434_
timestamp 1667941163
transform -1 0 27416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _435_
timestamp 1667941163
transform -1 0 28060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _436_
timestamp 1667941163
transform -1 0 27416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _437_
timestamp 1667941163
transform -1 0 28336 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _438_
timestamp 1667941163
transform -1 0 27692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _439_
timestamp 1667941163
transform -1 0 27232 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _440_
timestamp 1667941163
transform -1 0 25944 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _441_
timestamp 1667941163
transform -1 0 28704 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _442_
timestamp 1667941163
transform -1 0 32568 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _443_
timestamp 1667941163
transform -1 0 30636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _444_
timestamp 1667941163
transform -1 0 29256 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _445_
timestamp 1667941163
transform -1 0 31280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _446_
timestamp 1667941163
transform -1 0 31924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _447_
timestamp 1667941163
transform -1 0 28980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _448_
timestamp 1667941163
transform -1 0 29256 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _449_
timestamp 1667941163
transform -1 0 30636 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _450_
timestamp 1667941163
transform -1 0 29348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _451_
timestamp 1667941163
transform -1 0 29992 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _452_
timestamp 1667941163
transform -1 0 30636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _453_
timestamp 1667941163
transform 1 0 32292 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _454_
timestamp 1667941163
transform -1 0 32568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _455_
timestamp 1667941163
transform -1 0 29992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _456_
timestamp 1667941163
transform -1 0 29992 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _457_
timestamp 1667941163
transform -1 0 31280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _458_
timestamp 1667941163
transform -1 0 30268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _459_
timestamp 1667941163
transform -1 0 32568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _460_
timestamp 1667941163
transform -1 0 29348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _461_
timestamp 1667941163
transform -1 0 29992 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _462_
timestamp 1667941163
transform -1 0 30636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _463_
timestamp 1667941163
transform 1 0 32936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _464_
timestamp 1667941163
transform -1 0 24564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _465_
timestamp 1667941163
transform -1 0 26496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _466_
timestamp 1667941163
transform -1 0 25760 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _467_
timestamp 1667941163
transform -1 0 25208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _468_
timestamp 1667941163
transform -1 0 27416 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _469_
timestamp 1667941163
transform -1 0 25024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _470_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14536 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _471_
timestamp 1667941163
transform 1 0 11960 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _472_
timestamp 1667941163
transform -1 0 16468 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _473_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 18492 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _474_
timestamp 1667941163
transform 1 0 17204 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _475_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _476_
timestamp 1667941163
transform -1 0 26404 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _477_
timestamp 1667941163
transform 1 0 24564 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _478_
timestamp 1667941163
transform 1 0 21988 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _479_
timestamp 1667941163
transform 1 0 14352 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _480_
timestamp 1667941163
transform 1 0 14536 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _481_
timestamp 1667941163
transform 1 0 18584 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _482_
timestamp 1667941163
transform 1 0 17112 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _483_
timestamp 1667941163
transform 1 0 14904 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _484_
timestamp 1667941163
transform 1 0 12328 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _485_
timestamp 1667941163
transform -1 0 20240 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _486_
timestamp 1667941163
transform 1 0 21712 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _487_
timestamp 1667941163
transform -1 0 23920 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _488_
timestamp 1667941163
transform 1 0 11960 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _489_
timestamp 1667941163
transform 1 0 17112 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _490_
timestamp 1667941163
transform 1 0 14536 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _491_
timestamp 1667941163
transform 1 0 17940 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _492_
timestamp 1667941163
transform 1 0 21620 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _493_
timestamp 1667941163
transform 1 0 21160 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _494_
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _495_
timestamp 1667941163
transform 1 0 24196 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _496_
timestamp 1667941163
transform -1 0 26312 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _497_
timestamp 1667941163
transform 1 0 21988 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _498_
timestamp 1667941163
transform 1 0 21988 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _499_
timestamp 1667941163
transform 1 0 21988 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _500_
timestamp 1667941163
transform 1 0 12328 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _501_
timestamp 1667941163
transform -1 0 13800 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _502_
timestamp 1667941163
transform 1 0 11960 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _503_
timestamp 1667941163
transform 1 0 19412 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _504_
timestamp 1667941163
transform 1 0 14444 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _505_
timestamp 1667941163
transform -1 0 24104 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _506_
timestamp 1667941163
transform 1 0 12328 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _507_
timestamp 1667941163
transform -1 0 13800 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _508_
timestamp 1667941163
transform 1 0 17388 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _509_
timestamp 1667941163
transform 1 0 14536 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _510_
timestamp 1667941163
transform 1 0 16836 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _511_
timestamp 1667941163
transform 1 0 15548 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _512_
timestamp 1667941163
transform 1 0 14536 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _513_
timestamp 1667941163
transform 1 0 14628 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _514_
timestamp 1667941163
transform 1 0 19596 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _515_
timestamp 1667941163
transform 1 0 17020 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _516_
timestamp 1667941163
transform 1 0 14444 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _517_
timestamp 1667941163
transform 1 0 14444 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _518_
timestamp 1667941163
transform 1 0 17112 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _519_
timestamp 1667941163
transform 1 0 17204 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _520_
timestamp 1667941163
transform 1 0 14536 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _521_
timestamp 1667941163
transform -1 0 23644 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _522_
timestamp 1667941163
transform 1 0 18768 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _523_
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _524_
timestamp 1667941163
transform -1 0 23828 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _525_
timestamp 1667941163
transform -1 0 23184 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _526_
timestamp 1667941163
transform 1 0 21528 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _527_
timestamp 1667941163
transform 1 0 21988 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _528_
timestamp 1667941163
transform 1 0 17020 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _529_
timestamp 1667941163
transform 1 0 19412 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _530_
timestamp 1667941163
transform 1 0 16836 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _531_
timestamp 1667941163
transform 1 0 12236 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _532_
timestamp 1667941163
transform -1 0 13892 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _533_
timestamp 1667941163
transform 1 0 14260 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _534_
timestamp 1667941163
transform 1 0 20976 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _535_
timestamp 1667941163
transform 1 0 19596 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  _547_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 19780 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _548_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9108 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _549_
timestamp 1667941163
transform 1 0 6532 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _550_
timestamp 1667941163
transform -1 0 28060 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _551_
timestamp 1667941163
transform -1 0 22264 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _552_
timestamp 1667941163
transform 1 0 18860 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _553_
timestamp 1667941163
transform -1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _554_
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _555_
timestamp 1667941163
transform -1 0 17572 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _556_
timestamp 1667941163
transform 1 0 10396 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _557_
timestamp 1667941163
transform -1 0 22356 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _558_
timestamp 1667941163
transform -1 0 22356 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _559_
timestamp 1667941163
transform -1 0 22448 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _560_
timestamp 1667941163
transform -1 0 27048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _561_
timestamp 1667941163
transform 1 0 15272 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _562_
timestamp 1667941163
transform 1 0 28244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _563_
timestamp 1667941163
transform -1 0 29992 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _564_
timestamp 1667941163
transform -1 0 36984 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _565_
timestamp 1667941163
transform -1 0 14628 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _566_
timestamp 1667941163
transform 1 0 10948 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _567_
timestamp 1667941163
transform -1 0 28704 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _568_
timestamp 1667941163
transform 1 0 31096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _569_
timestamp 1667941163
transform 1 0 5060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _570_
timestamp 1667941163
transform 1 0 1932 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _571_
timestamp 1667941163
transform 1 0 4600 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _572_
timestamp 1667941163
transform -1 0 38088 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _573_
timestamp 1667941163
transform 1 0 2300 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _574_
timestamp 1667941163
transform -1 0 20332 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _575_
timestamp 1667941163
transform -1 0 28796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _576_
timestamp 1667941163
transform 1 0 16192 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _577_
timestamp 1667941163
transform -1 0 33856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _578_
timestamp 1667941163
transform 1 0 1748 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _579_
timestamp 1667941163
transform 1 0 27876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _580_
timestamp 1667941163
transform 1 0 12512 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _581_
timestamp 1667941163
transform -1 0 20056 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _582_
timestamp 1667941163
transform 1 0 24380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _583_
timestamp 1667941163
transform -1 0 27508 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _584_
timestamp 1667941163
transform -1 0 25944 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _585_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14260 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _586_
timestamp 1667941163
transform -1 0 17756 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _587_
timestamp 1667941163
transform 1 0 12788 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _588_
timestamp 1667941163
transform 1 0 12788 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _589_
timestamp 1667941163
transform 1 0 14352 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _589__91 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 14076 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _590_
timestamp 1667941163
transform -1 0 25116 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _591_
timestamp 1667941163
transform -1 0 10580 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _592_
timestamp 1667941163
transform -1 0 12512 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _593_
timestamp 1667941163
transform -1 0 18952 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _594_
timestamp 1667941163
transform 1 0 12880 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _595_
timestamp 1667941163
transform 1 0 11776 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _596_
timestamp 1667941163
transform -1 0 12788 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _597_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22908 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _598_
timestamp 1667941163
transform 1 0 12972 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _599_
timestamp 1667941163
transform 1 0 27140 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _600_
timestamp 1667941163
transform 1 0 20516 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _601_
timestamp 1667941163
transform 1 0 15364 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _601__92
timestamp 1667941163
transform -1 0 10856 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _602_
timestamp 1667941163
transform 1 0 28704 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _603_
timestamp 1667941163
transform -1 0 25392 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _604_
timestamp 1667941163
transform 1 0 18860 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _605_
timestamp 1667941163
transform 1 0 24840 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _606_
timestamp 1667941163
transform 1 0 12972 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _607_
timestamp 1667941163
transform 1 0 21988 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _608_
timestamp 1667941163
transform 1 0 20056 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _609_
timestamp 1667941163
transform 1 0 16836 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _610_
timestamp 1667941163
transform 1 0 20056 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _611_
timestamp 1667941163
transform -1 0 23000 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _612_
timestamp 1667941163
transform 1 0 20148 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _612__93
timestamp 1667941163
transform -1 0 19780 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _613_
timestamp 1667941163
transform 1 0 23000 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _614_
timestamp 1667941163
transform 1 0 15180 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _615_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 20148 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _616_
timestamp 1667941163
transform -1 0 22724 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _617_
timestamp 1667941163
transform 1 0 20332 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _618_
timestamp 1667941163
transform 1 0 15364 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _619_
timestamp 1667941163
transform -1 0 25668 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _620_
timestamp 1667941163
transform -1 0 22356 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _621_
timestamp 1667941163
transform -1 0 23184 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _622_
timestamp 1667941163
transform 1 0 17756 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _623_
timestamp 1667941163
transform 1 0 16836 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _624__94
timestamp 1667941163
transform 1 0 20976 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _624_
timestamp 1667941163
transform -1 0 20608 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _625_
timestamp 1667941163
transform 1 0 20240 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _626_
timestamp 1667941163
transform -1 0 26312 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _627_
timestamp 1667941163
transform -1 0 26588 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _628_
timestamp 1667941163
transform -1 0 25944 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _629_
timestamp 1667941163
transform -1 0 22172 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _630_
timestamp 1667941163
transform -1 0 21160 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _631_
timestamp 1667941163
transform -1 0 26864 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _632_
timestamp 1667941163
transform -1 0 24288 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _633_
timestamp 1667941163
transform 1 0 24840 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _634_
timestamp 1667941163
transform 1 0 25668 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _635_
timestamp 1667941163
transform 1 0 16836 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _636_
timestamp 1667941163
transform 1 0 23276 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _636__95
timestamp 1667941163
transform 1 0 23368 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _637_
timestamp 1667941163
transform -1 0 24932 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _638_
timestamp 1667941163
transform 1 0 18676 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _639_
timestamp 1667941163
transform -1 0 28428 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _640_
timestamp 1667941163
transform 1 0 25208 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _641_
timestamp 1667941163
transform 1 0 26864 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _642_
timestamp 1667941163
transform 1 0 22908 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _643_
timestamp 1667941163
transform -1 0 20056 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _644_
timestamp 1667941163
transform -1 0 26588 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _645_
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _646_
timestamp 1667941163
transform -1 0 13248 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _647_
timestamp 1667941163
transform 1 0 12052 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _648__96
timestamp 1667941163
transform -1 0 9292 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _648_
timestamp 1667941163
transform 1 0 11684 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _649_
timestamp 1667941163
transform 1 0 14260 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _650_
timestamp 1667941163
transform 1 0 11776 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _651_
timestamp 1667941163
transform -1 0 16376 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _652_
timestamp 1667941163
transform 1 0 25484 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _653_
timestamp 1667941163
transform -1 0 15364 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _654_
timestamp 1667941163
transform 1 0 20148 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _655_
timestamp 1667941163
transform -1 0 23092 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _656_
timestamp 1667941163
transform -1 0 25392 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _657_
timestamp 1667941163
transform 1 0 13432 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _658_
timestamp 1667941163
transform 1 0 13800 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _659_
timestamp 1667941163
transform -1 0 26588 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _660__97
timestamp 1667941163
transform -1 0 9936 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _660_
timestamp 1667941163
transform 1 0 12972 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _661_
timestamp 1667941163
transform 1 0 11868 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _662_
timestamp 1667941163
transform 1 0 13064 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _663_
timestamp 1667941163
transform 1 0 23276 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _664_
timestamp 1667941163
transform 1 0 13984 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _665_
timestamp 1667941163
transform -1 0 16928 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _666_
timestamp 1667941163
transform 1 0 13156 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _667_
timestamp 1667941163
transform -1 0 14996 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _668_
timestamp 1667941163
transform -1 0 25668 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _669_
timestamp 1667941163
transform 1 0 26956 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _670_
timestamp 1667941163
transform 1 0 25760 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _671_
timestamp 1667941163
transform 1 0 13156 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _672__98
timestamp 1667941163
transform -1 0 11960 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _672_
timestamp 1667941163
transform 1 0 15456 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _673_
timestamp 1667941163
transform -1 0 18492 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _674_
timestamp 1667941163
transform -1 0 25760 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _675_
timestamp 1667941163
transform 1 0 18124 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _676_
timestamp 1667941163
transform 1 0 18400 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _677_
timestamp 1667941163
transform 1 0 25760 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _678_
timestamp 1667941163
transform 1 0 13984 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _679_
timestamp 1667941163
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _680_
timestamp 1667941163
transform 1 0 19412 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _681_
timestamp 1667941163
transform -1 0 15180 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _682_
timestamp 1667941163
transform -1 0 15916 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _683_
timestamp 1667941163
transform -1 0 25484 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _684_
timestamp 1667941163
transform 1 0 15548 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _684__99
timestamp 1667941163
transform -1 0 12236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _685_
timestamp 1667941163
transform 1 0 23184 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _686_
timestamp 1667941163
transform 1 0 12972 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _687_
timestamp 1667941163
transform 1 0 21712 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _688_
timestamp 1667941163
transform -1 0 21160 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _689_
timestamp 1667941163
transform -1 0 13064 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _690_
timestamp 1667941163
transform 1 0 15548 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _691_
timestamp 1667941163
transform -1 0 27232 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _692_
timestamp 1667941163
transform -1 0 23736 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _693_
timestamp 1667941163
transform 1 0 17848 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _694_
timestamp 1667941163
transform -1 0 18952 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _695_
timestamp 1667941163
transform 1 0 15548 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _696_
timestamp 1667941163
transform -1 0 19964 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _696__100
timestamp 1667941163
transform -1 0 19688 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _697_
timestamp 1667941163
transform 1 0 20792 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _698_
timestamp 1667941163
transform -1 0 24104 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _699_
timestamp 1667941163
transform -1 0 26128 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _700_
timestamp 1667941163
transform 1 0 23000 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _701_
timestamp 1667941163
transform -1 0 22632 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _702_
timestamp 1667941163
transform -1 0 19872 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _703_
timestamp 1667941163
transform 1 0 16560 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _704_
timestamp 1667941163
transform -1 0 25392 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _705_
timestamp 1667941163
transform -1 0 17756 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _706_
timestamp 1667941163
transform -1 0 17756 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _707_
timestamp 1667941163
transform 1 0 16836 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _708_
timestamp 1667941163
transform -1 0 19596 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _708__101
timestamp 1667941163
transform 1 0 19412 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _709_
timestamp 1667941163
transform -1 0 24012 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _710_
timestamp 1667941163
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _711_
timestamp 1667941163
transform -1 0 25392 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _712_
timestamp 1667941163
transform 1 0 19872 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _713_
timestamp 1667941163
transform -1 0 16560 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _714_
timestamp 1667941163
transform -1 0 22816 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _715_
timestamp 1667941163
transform -1 0 25392 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _716_
timestamp 1667941163
transform -1 0 25392 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform -1 0 1840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1667941163
transform 1 0 1564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1667941163
transform -1 0 35972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14904 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1667941163
transform -1 0 18492 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1667941163
transform 1 0 16836 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1667941163
transform -1 0 38364 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1667941163
transform 1 0 35512 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1667941163
transform -1 0 11224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1667941163
transform -1 0 38364 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1667941163
transform -1 0 38364 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1667941163
transform -1 0 38364 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1667941163
transform -1 0 38364 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1667941163
transform -1 0 38364 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1667941163
transform 1 0 1564 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1667941163
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1667941163
transform -1 0 38364 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1667941163
transform 1 0 1564 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1667941163
transform -1 0 38364 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1667941163
transform 1 0 1564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1667941163
transform 1 0 1564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1667941163
transform 1 0 1564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1667941163
transform -1 0 38364 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1667941163
transform 1 0 7820 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1667941163
transform -1 0 3496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1667941163
transform -1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1667941163
transform 1 0 32936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1667941163
transform -1 0 38364 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1667941163
transform -1 0 38364 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1667941163
transform -1 0 28244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1667941163
transform 1 0 2300 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1667941163
transform -1 0 38364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1667941163
transform 1 0 1564 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1667941163
transform -1 0 38364 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1667941163
transform 1 0 1564 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1667941163
transform -1 0 32568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1667941163
transform -1 0 38364 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 37812 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1667941163
transform -1 0 1932 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1667941163
transform 1 0 37996 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1667941163
transform 1 0 37444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1667941163
transform 1 0 25208 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1667941163
transform -1 0 1932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1667941163
transform 1 0 37996 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1667941163
transform -1 0 1932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1667941163
transform -1 0 1932 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1667941163
transform -1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1667941163
transform -1 0 30728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1667941163
transform -1 0 1932 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1667941163
transform 1 0 28428 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1667941163
transform 1 0 37996 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1667941163
transform -1 0 27508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1667941163
transform -1 0 1932 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1667941163
transform 1 0 36616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1667941163
transform 1 0 37996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1667941163
transform -1 0 12052 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1667941163
transform -1 0 6900 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1667941163
transform 1 0 19412 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1667941163
transform -1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1667941163
transform -1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1667941163
transform -1 0 13340 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1667941163
transform 1 0 23276 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1667941163
transform 1 0 33580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1667941163
transform -1 0 1932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1667941163
transform -1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1667941163
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1667941163
transform 1 0 30360 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1667941163
transform -1 0 20516 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1667941163
transform 1 0 37260 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1667941163
transform 1 0 37996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1667941163
transform -1 0 4968 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1667941163
transform 1 0 37996 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1667941163
transform -1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1667941163
transform 1 0 10856 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1667941163
transform -1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1667941163
transform -1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform -1 0 3036 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform -1 0 10120 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform -1 0 27508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform -1 0 1932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform -1 0 1932 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform 1 0 37996 0 -1 19584
box -38 -48 406 592
<< labels >>
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 ccff_head
port 0 nsew signal input
flabel metal2 s 37370 39200 37426 39800 0 FreeSans 224 90 0 0 ccff_tail
port 1 nsew signal tristate
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 chany_bottom_in[0]
port 2 nsew signal input
flabel metal2 s 35438 200 35494 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 3 nsew signal input
flabel metal2 s 14830 39200 14886 39800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 4 nsew signal input
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 5 nsew signal input
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 6 nsew signal input
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 7 nsew signal input
flabel metal3 s 39200 8168 39800 8288 0 FreeSans 480 0 0 0 chany_bottom_in[15]
port 8 nsew signal input
flabel metal2 s 35438 39200 35494 39800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 9 nsew signal input
flabel metal2 s 21914 39200 21970 39800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 10 nsew signal input
flabel metal2 s 13542 200 13598 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 11 nsew signal input
flabel metal3 s 39200 11568 39800 11688 0 FreeSans 480 0 0 0 chany_bottom_in[1]
port 12 nsew signal input
flabel metal3 s 39200 17008 39800 17128 0 FreeSans 480 0 0 0 chany_bottom_in[2]
port 13 nsew signal input
flabel metal3 s 39200 35368 39800 35488 0 FreeSans 480 0 0 0 chany_bottom_in[3]
port 14 nsew signal input
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chany_bottom_in[4]
port 15 nsew signal input
flabel metal3 s 39200 4768 39800 4888 0 FreeSans 480 0 0 0 chany_bottom_in[5]
port 16 nsew signal input
flabel metal3 s 200 28568 800 28688 0 FreeSans 480 0 0 0 chany_bottom_in[6]
port 17 nsew signal input
flabel metal2 s 8390 200 8446 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 18 nsew signal input
flabel metal3 s 39200 26528 39800 26648 0 FreeSans 480 0 0 0 chany_bottom_in[8]
port 19 nsew signal input
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 chany_bottom_in[9]
port 20 nsew signal input
flabel metal3 s 200 14288 800 14408 0 FreeSans 480 0 0 0 chany_bottom_out[0]
port 21 nsew signal tristate
flabel metal3 s 39200 27888 39800 28008 0 FreeSans 480 0 0 0 chany_bottom_out[10]
port 22 nsew signal tristate
flabel metal2 s 37370 200 37426 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 23 nsew signal tristate
flabel metal2 s 25134 39200 25190 39800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 24 nsew signal tristate
flabel metal2 s 1306 39200 1362 39800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 25 nsew signal tristate
flabel metal3 s 39200 29928 39800 30048 0 FreeSans 480 0 0 0 chany_bottom_out[14]
port 26 nsew signal tristate
flabel metal3 s 200 19728 800 19848 0 FreeSans 480 0 0 0 chany_bottom_out[15]
port 27 nsew signal tristate
flabel metal3 s 200 23128 800 23248 0 FreeSans 480 0 0 0 chany_bottom_out[16]
port 28 nsew signal tristate
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 chany_bottom_out[17]
port 29 nsew signal tristate
flabel metal2 s 30286 200 30342 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 30 nsew signal tristate
flabel metal3 s 200 34008 800 34128 0 FreeSans 480 0 0 0 chany_bottom_out[1]
port 31 nsew signal tristate
flabel metal2 s 27066 39200 27122 39800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 32 nsew signal tristate
flabel metal2 s 28354 39200 28410 39800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 33 nsew signal tristate
flabel metal2 s 34150 200 34206 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 34 nsew signal tristate
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 35 nsew signal tristate
flabel metal3 s 39200 33328 39800 33448 0 FreeSans 480 0 0 0 chany_bottom_out[6]
port 36 nsew signal tristate
flabel metal2 s 23846 200 23902 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 37 nsew signal tristate
flabel metal3 s 200 21088 800 21208 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 38 nsew signal tristate
flabel metal3 s 39200 688 39800 808 0 FreeSans 480 0 0 0 chany_bottom_out[9]
port 39 nsew signal tristate
flabel metal3 s 39200 15648 39800 15768 0 FreeSans 480 0 0 0 chany_top_in[0]
port 40 nsew signal input
flabel metal3 s 200 39448 800 39568 0 FreeSans 480 0 0 0 chany_top_in[10]
port 41 nsew signal input
flabel metal3 s 200 10208 800 10328 0 FreeSans 480 0 0 0 chany_top_in[11]
port 42 nsew signal input
flabel metal3 s 200 31968 800 32088 0 FreeSans 480 0 0 0 chany_top_in[12]
port 43 nsew signal input
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 chany_top_in[13]
port 44 nsew signal input
flabel metal3 s 39200 37408 39800 37528 0 FreeSans 480 0 0 0 chany_top_in[14]
port 45 nsew signal input
flabel metal2 s 7746 39200 7802 39800 0 FreeSans 224 90 0 0 chany_top_in[15]
port 46 nsew signal input
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chany_top_in[16]
port 47 nsew signal input
flabel metal2 s 9678 200 9734 800 0 FreeSans 224 90 0 0 chany_top_in[17]
port 48 nsew signal input
flabel metal2 s 32218 200 32274 800 0 FreeSans 224 90 0 0 chany_top_in[18]
port 49 nsew signal input
flabel metal3 s 39200 13608 39800 13728 0 FreeSans 480 0 0 0 chany_top_in[1]
port 50 nsew signal input
flabel metal3 s 39200 6128 39800 6248 0 FreeSans 480 0 0 0 chany_top_in[2]
port 51 nsew signal input
flabel metal2 s 25134 200 25190 800 0 FreeSans 224 90 0 0 chany_top_in[3]
port 52 nsew signal input
flabel metal3 s 200 37408 800 37528 0 FreeSans 480 0 0 0 chany_top_in[4]
port 53 nsew signal input
flabel metal2 s 39302 200 39358 800 0 FreeSans 224 90 0 0 chany_top_in[5]
port 54 nsew signal input
flabel metal3 s 200 8848 800 8968 0 FreeSans 480 0 0 0 chany_top_in[6]
port 55 nsew signal input
flabel metal3 s 39200 10208 39800 10328 0 FreeSans 480 0 0 0 chany_top_in[7]
port 56 nsew signal input
flabel metal3 s 200 25168 800 25288 0 FreeSans 480 0 0 0 chany_top_in[8]
port 57 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 chany_top_in[9]
port 58 nsew signal input
flabel metal3 s 39200 24488 39800 24608 0 FreeSans 480 0 0 0 chany_top_out[0]
port 59 nsew signal tristate
flabel metal2 s 11610 39200 11666 39800 0 FreeSans 224 90 0 0 chany_top_out[10]
port 60 nsew signal tristate
flabel metal2 s 6458 39200 6514 39800 0 FreeSans 224 90 0 0 chany_top_out[11]
port 61 nsew signal tristate
flabel metal2 s 18694 200 18750 800 0 FreeSans 224 90 0 0 chany_top_out[12]
port 62 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_top_out[13]
port 63 nsew signal tristate
flabel metal2 s 21914 200 21970 800 0 FreeSans 224 90 0 0 chany_top_out[14]
port 64 nsew signal tristate
flabel metal2 s 12898 39200 12954 39800 0 FreeSans 224 90 0 0 chany_top_out[15]
port 65 nsew signal tristate
flabel metal2 s 23202 39200 23258 39800 0 FreeSans 224 90 0 0 chany_top_out[16]
port 66 nsew signal tristate
flabel metal2 s 33506 39200 33562 39800 0 FreeSans 224 90 0 0 chany_top_out[17]
port 67 nsew signal tristate
flabel metal3 s 200 26528 800 26648 0 FreeSans 480 0 0 0 chany_top_out[18]
port 68 nsew signal tristate
flabel metal2 s 4526 200 4582 800 0 FreeSans 224 90 0 0 chany_top_out[1]
port 69 nsew signal tristate
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 chany_top_out[2]
port 70 nsew signal tristate
flabel metal2 s 38658 39200 38714 39800 0 FreeSans 224 90 0 0 chany_top_out[3]
port 71 nsew signal tristate
flabel metal2 s 30286 39200 30342 39800 0 FreeSans 224 90 0 0 chany_top_out[4]
port 72 nsew signal tristate
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 chany_top_out[5]
port 73 nsew signal tristate
flabel metal3 s 39200 38768 39800 38888 0 FreeSans 480 0 0 0 chany_top_out[6]
port 74 nsew signal tristate
flabel metal3 s 39200 2728 39800 2848 0 FreeSans 480 0 0 0 chany_top_out[7]
port 75 nsew signal tristate
flabel metal2 s 4526 39200 4582 39800 0 FreeSans 224 90 0 0 chany_top_out[8]
port 76 nsew signal tristate
flabel metal3 s 39200 21088 39800 21208 0 FreeSans 480 0 0 0 chany_top_out[9]
port 77 nsew signal tristate
flabel metal2 s 6458 200 6514 800 0 FreeSans 224 90 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_1_
port 78 nsew signal tristate
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_5_
port 79 nsew signal tristate
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 left_grid_right_width_0_height_0_subtile_0__pin_I_9_
port 80 nsew signal tristate
flabel metal3 s 39200 22448 39800 22568 0 FreeSans 480 0 0 0 pReset
port 81 nsew signal input
flabel metal2 s 19982 200 20038 800 0 FreeSans 224 90 0 0 prog_clk
port 82 nsew signal input
flabel metal3 s 200 4768 800 4888 0 FreeSans 480 0 0 0 right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_
port 83 nsew signal tristate
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_
port 84 nsew signal tristate
flabel metal2 s 2594 39200 2650 39800 0 FreeSans 224 90 0 0 right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_
port 85 nsew signal tristate
flabel metal2 s 9678 39200 9734 39800 0 FreeSans 224 90 0 0 right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_
port 86 nsew signal tristate
flabel metal2 s 27066 200 27122 800 0 FreeSans 224 90 0 0 right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_
port 87 nsew signal tristate
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_
port 88 nsew signal tristate
flabel metal3 s 200 36048 800 36168 0 FreeSans 480 0 0 0 right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_
port 89 nsew signal tristate
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_
port 90 nsew signal tristate
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 91 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 91 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 92 nsew ground bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal2 17342 2210 17342 2210 0 _000_
rlabel metal2 13386 2686 13386 2686 0 _001_
rlabel metal1 15877 4522 15877 4522 0 _002_
rlabel metal1 17855 11050 17855 11050 0 _003_
rlabel metal1 26128 8058 26128 8058 0 _004_
rlabel metal1 21167 2346 21167 2346 0 _005_
rlabel metal2 25622 2108 25622 2108 0 _006_
rlabel metal1 27285 3434 27285 3434 0 _007_
rlabel metal2 27370 6392 27370 6392 0 _008_
rlabel metal1 16245 8942 16245 8942 0 _009_
rlabel metal1 16291 9962 16291 9962 0 _010_
rlabel metal2 28750 2176 28750 2176 0 _011_
rlabel metal2 21206 4692 21206 4692 0 _012_
rlabel metal1 16889 5610 16889 5610 0 _013_
rlabel metal2 13754 6086 13754 6086 0 _014_
rlabel metal1 20838 9554 20838 9554 0 _015_
rlabel metal1 25261 7786 25261 7786 0 _016_
rlabel metal1 25537 6358 25537 6358 0 _017_
rlabel metal1 13531 4590 13531 4590 0 _018_
rlabel metal1 18538 2523 18538 2523 0 _019_
rlabel metal1 20470 6392 20470 6392 0 _020_
rlabel metal1 27922 7514 27922 7514 0 _021_
rlabel metal1 28106 7922 28106 7922 0 _022_
rlabel metal2 27278 6494 27278 6494 0 _023_
rlabel metal1 23973 2414 23973 2414 0 _024_
rlabel metal2 28842 4590 28842 4590 0 _025_
rlabel metal2 25530 3332 25530 3332 0 _026_
rlabel via2 27462 7701 27462 7701 0 _027_
rlabel metal1 28290 9078 28290 9078 0 _028_
rlabel metal1 26174 6902 26174 6902 0 _029_
rlabel metal2 13754 2771 13754 2771 0 _030_
rlabel via2 12374 2397 12374 2397 0 _031_
rlabel metal1 14589 6698 14589 6698 0 _032_
rlabel metal2 27922 7497 27922 7497 0 _033_
rlabel metal2 21298 7072 21298 7072 0 _034_
rlabel metal2 23322 3400 23322 3400 0 _035_
rlabel metal2 13754 5151 13754 5151 0 _036_
rlabel metal2 12374 5729 12374 5729 0 _037_
rlabel metal1 20286 5304 20286 5304 0 _038_
rlabel metal1 16659 7786 16659 7786 0 _039_
rlabel metal1 18591 8874 18591 8874 0 _040_
rlabel metal1 18177 6698 18177 6698 0 _041_
rlabel via2 16514 5253 16514 5253 0 _042_
rlabel metal2 31786 2652 31786 2652 0 _043_
rlabel metal2 22402 5202 22402 5202 0 _044_
rlabel metal2 18354 10047 18354 10047 0 _045_
rlabel metal2 20102 8313 20102 8313 0 _046_
rlabel metal2 18538 7973 18538 7973 0 _047_
rlabel metal2 21298 5593 21298 5593 0 _048_
rlabel metal2 20378 3774 20378 3774 0 _049_
rlabel metal2 19826 2992 19826 2992 0 _050_
rlabel metal1 23053 8874 23053 8874 0 _051_
rlabel via2 28750 8381 28750 8381 0 _052_
rlabel via2 19182 6307 19182 6307 0 _053_
rlabel metal1 23743 4182 23743 4182 0 _054_
rlabel metal2 30406 3978 30406 3978 0 _055_
rlabel metal1 29164 4114 29164 4114 0 _056_
rlabel metal2 29854 8024 29854 8024 0 _057_
rlabel metal1 18959 7786 18959 7786 0 _058_
rlabel metal2 28658 3213 28658 3213 0 _059_
rlabel metal1 18262 3543 18262 3543 0 _060_
rlabel metal2 26358 7735 26358 7735 0 _061_
rlabel metal1 13301 4182 13301 4182 0 _062_
rlabel via1 21942 5083 21942 5083 0 _063_
rlabel metal1 22823 3502 22823 3502 0 _064_
rlabel metal2 21022 10166 21022 10166 0 _065_
rlabel metal2 30222 9486 30222 9486 0 _066_
rlabel metal2 29946 9758 29946 9758 0 _067_
rlabel metal1 28796 10574 28796 10574 0 _068_
rlabel metal1 29762 5202 29762 5202 0 _069_
rlabel metal1 28704 9962 28704 9962 0 _070_
rlabel metal2 31878 4046 31878 4046 0 _071_
rlabel metal1 32522 3468 32522 3468 0 _072_
rlabel metal1 13524 15674 13524 15674 0 _073_
rlabel metal1 15686 9112 15686 9112 0 _074_
rlabel metal2 13018 16286 13018 16286 0 _075_
rlabel metal1 10396 13974 10396 13974 0 _076_
rlabel metal1 14582 10744 14582 10744 0 _077_
rlabel via2 22218 9605 22218 9605 0 _078_
rlabel metal1 10396 9622 10396 9622 0 _079_
rlabel metal2 12282 9010 12282 9010 0 _080_
rlabel metal1 18722 14280 18722 14280 0 _081_
rlabel metal2 13386 10744 13386 10744 0 _082_
rlabel metal2 9890 10540 9890 10540 0 _083_
rlabel metal1 13202 7514 13202 7514 0 _084_
rlabel metal1 27370 13770 27370 13770 0 _085_
rlabel metal1 13202 13192 13202 13192 0 _086_
rlabel metal1 27830 10710 27830 10710 0 _087_
rlabel metal2 20746 11288 20746 11288 0 _088_
rlabel metal1 13294 13770 13294 13770 0 _089_
rlabel metal2 28198 9282 28198 9282 0 _090_
rlabel metal1 25162 11016 25162 11016 0 _091_
rlabel metal2 19090 11934 19090 11934 0 _092_
rlabel metal1 24978 8058 24978 8058 0 _093_
rlabel via2 13202 14331 13202 14331 0 _094_
rlabel metal2 20838 11934 20838 11934 0 _095_
rlabel metal1 19964 14246 19964 14246 0 _096_
rlabel metal2 16054 13753 16054 13753 0 _097_
rlabel metal2 19734 12274 19734 12274 0 _098_
rlabel metal2 21390 15810 21390 15810 0 _099_
rlabel metal1 20562 16490 20562 16490 0 _100_
rlabel metal1 27094 15062 27094 15062 0 _101_
rlabel metal2 15410 16286 15410 16286 0 _102_
rlabel metal2 19918 11254 19918 11254 0 _103_
rlabel metal1 21367 13974 21367 13974 0 _104_
rlabel metal1 19734 12920 19734 12920 0 _105_
rlabel metal1 19826 11288 19826 11288 0 _106_
rlabel metal1 25438 14280 25438 14280 0 _107_
rlabel metal2 21390 11968 21390 11968 0 _108_
rlabel metal2 20746 9214 20746 9214 0 _109_
rlabel metal1 17848 16422 17848 16422 0 _110_
rlabel metal2 18354 16728 18354 16728 0 _111_
rlabel metal1 20286 18666 20286 18666 0 _112_
rlabel metal1 20654 14314 20654 14314 0 _113_
rlabel metal1 27324 13974 27324 13974 0 _114_
rlabel metal2 26358 15640 26358 15640 0 _115_
rlabel metal1 26818 16150 26818 16150 0 _116_
rlabel metal1 21528 13226 21528 13226 0 _117_
rlabel metal1 21505 16150 21505 16150 0 _118_
rlabel metal2 26634 15368 26634 15368 0 _119_
rlabel metal1 24104 12886 24104 12886 0 _120_
rlabel metal2 24702 7106 24702 7106 0 _121_
rlabel metal1 25070 6834 25070 6834 0 _122_
rlabel metal2 17066 14382 17066 14382 0 _123_
rlabel metal1 24058 17238 24058 17238 0 _124_
rlabel metal1 26358 14586 26358 14586 0 _125_
rlabel metal2 21022 17850 21022 17850 0 _126_
rlabel metal2 28198 14280 28198 14280 0 _127_
rlabel metal2 25438 17374 25438 17374 0 _128_
rlabel metal1 25254 6630 25254 6630 0 _129_
rlabel metal1 23322 17578 23322 17578 0 _130_
rlabel metal1 20516 17238 20516 17238 0 _131_
rlabel metal1 26404 16218 26404 16218 0 _132_
rlabel metal2 12558 11186 12558 11186 0 _133_
rlabel metal2 13294 8806 13294 8806 0 _134_
rlabel metal1 12282 8840 12282 8840 0 _135_
rlabel metal1 12006 12886 12006 12886 0 _136_
rlabel metal1 14536 15402 14536 15402 0 _137_
rlabel metal1 11684 10166 11684 10166 0 _138_
rlabel metal2 16606 16898 16606 16898 0 _139_
rlabel metal3 25116 10268 25116 10268 0 _140_
rlabel metal2 13478 11696 13478 11696 0 _141_
rlabel metal1 20378 17544 20378 17544 0 _142_
rlabel metal1 22908 12886 22908 12886 0 _143_
rlabel metal1 25116 17578 25116 17578 0 _144_
rlabel metal1 10396 11866 10396 11866 0 _145_
rlabel metal2 13938 10574 13938 10574 0 _146_
rlabel metal1 26864 9622 26864 9622 0 _147_
rlabel metal1 11178 9962 11178 9962 0 _148_
rlabel metal2 12098 14076 12098 14076 0 _149_
rlabel metal1 12604 15538 12604 15538 0 _150_
rlabel via2 23506 12155 23506 12155 0 _151_
rlabel metal1 14214 16184 14214 16184 0 _152_
rlabel metal2 16698 11186 16698 11186 0 _153_
rlabel metal2 10166 11679 10166 11679 0 _154_
rlabel metal1 14168 11186 14168 11186 0 _155_
rlabel metal1 25806 11798 25806 11798 0 _156_
rlabel metal1 27784 9622 27784 9622 0 _157_
rlabel metal1 28060 12954 28060 12954 0 _158_
rlabel metal1 12926 12818 12926 12818 0 _159_
rlabel metal1 16192 13974 16192 13974 0 _160_
rlabel metal2 18262 9656 18262 9656 0 _161_
rlabel metal1 25898 9622 25898 9622 0 _162_
rlabel metal1 19642 9894 19642 9894 0 _163_
rlabel metal2 18630 16286 18630 16286 0 _164_
rlabel metal1 27508 12138 27508 12138 0 _165_
rlabel metal2 14214 16014 14214 16014 0 _166_
rlabel metal1 14168 9010 14168 9010 0 _167_
rlabel metal2 17250 16014 17250 16014 0 _168_
rlabel metal1 15180 12886 15180 12886 0 _169_
rlabel metal2 14214 13685 14214 13685 0 _170_
rlabel metal1 25173 12886 25173 12886 0 _171_
rlabel via2 21206 8483 21206 8483 0 _172_
rlabel metal2 23414 14025 23414 14025 0 _173_
rlabel metal1 13202 12104 13202 12104 0 _174_
rlabel metal1 21620 13838 21620 13838 0 _175_
rlabel metal2 20930 9418 20930 9418 0 _176_
rlabel metal1 10212 13498 10212 13498 0 _177_
rlabel metal1 16514 12886 16514 12886 0 _178_
rlabel metal1 26220 8262 26220 8262 0 _179_
rlabel metal2 23506 11288 23506 11288 0 _180_
rlabel metal1 15778 12682 15778 12682 0 _181_
rlabel metal1 19642 13158 19642 13158 0 _182_
rlabel metal2 15778 16286 15778 16286 0 _183_
rlabel metal1 20010 13974 20010 13974 0 _184_
rlabel metal2 21022 16184 21022 16184 0 _185_
rlabel metal1 23874 11832 23874 11832 0 _186_
rlabel metal1 25944 15062 25944 15062 0 _187_
rlabel metal1 23092 14314 23092 14314 0 _188_
rlabel metal2 27094 13583 27094 13583 0 _189_
rlabel metal2 20378 15640 20378 15640 0 _190_
rlabel metal2 16790 13838 16790 13838 0 _191_
rlabel metal2 25162 13838 25162 13838 0 _192_
rlabel metal2 17526 14416 17526 14416 0 _193_
rlabel metal2 17526 16456 17526 16456 0 _194_
rlabel metal1 16744 16150 16744 16150 0 _195_
rlabel metal1 19458 20026 19458 20026 0 _196_
rlabel metal1 23920 16150 23920 16150 0 _197_
rlabel metal1 16652 18326 16652 18326 0 _198_
rlabel metal2 25162 16728 25162 16728 0 _199_
rlabel metal2 20102 19006 20102 19006 0 _200_
rlabel metal1 10626 12614 10626 12614 0 _201_
rlabel metal1 22494 17850 22494 17850 0 _202_
rlabel metal1 26542 12274 26542 12274 0 _203_
rlabel metal1 25162 16456 25162 16456 0 _204_
rlabel via2 1610 3485 1610 3485 0 ccff_head
rlabel metal1 37490 36890 37490 36890 0 ccff_tail
rlabel via2 1610 17765 1610 17765 0 chany_bottom_in[0]
rlabel metal1 35650 2346 35650 2346 0 chany_bottom_in[10]
rlabel metal1 14904 37298 14904 37298 0 chany_bottom_in[11]
rlabel metal2 16698 37383 16698 37383 0 chany_bottom_in[12]
rlabel metal1 17894 37434 17894 37434 0 chany_bottom_in[13]
rlabel metal2 16882 4199 16882 4199 0 chany_bottom_in[14]
rlabel metal2 38226 8347 38226 8347 0 chany_bottom_in[15]
rlabel metal1 35512 37298 35512 37298 0 chany_bottom_in[16]
rlabel metal1 21988 37298 21988 37298 0 chany_bottom_in[17]
rlabel metal1 11132 2414 11132 2414 0 chany_bottom_in[18]
rlabel metal2 38226 11679 38226 11679 0 chany_bottom_in[1]
rlabel metal2 38226 17119 38226 17119 0 chany_bottom_in[2]
rlabel metal2 38318 35343 38318 35343 0 chany_bottom_in[3]
rlabel via2 38318 32011 38318 32011 0 chany_bottom_in[4]
rlabel via2 38318 4811 38318 4811 0 chany_bottom_in[5]
rlabel via2 1610 28645 1610 28645 0 chany_bottom_in[6]
rlabel metal2 8418 1554 8418 1554 0 chany_bottom_in[7]
rlabel via2 38318 26571 38318 26571 0 chany_bottom_in[8]
rlabel via2 1702 30651 1702 30651 0 chany_bottom_in[9]
rlabel metal3 1188 14348 1188 14348 0 chany_bottom_out[0]
rlabel via2 38226 27931 38226 27931 0 chany_bottom_out[10]
rlabel metal2 37398 1520 37398 1520 0 chany_bottom_out[11]
rlabel metal1 25300 37094 25300 37094 0 chany_bottom_out[12]
rlabel metal1 1518 37094 1518 37094 0 chany_bottom_out[13]
rlabel via2 38226 30005 38226 30005 0 chany_bottom_out[14]
rlabel metal3 1188 19788 1188 19788 0 chany_bottom_out[15]
rlabel metal3 1188 23188 1188 23188 0 chany_bottom_out[16]
rlabel metal3 1188 1428 1188 1428 0 chany_bottom_out[17]
rlabel metal2 30314 1520 30314 1520 0 chany_bottom_out[18]
rlabel metal3 1188 34068 1188 34068 0 chany_bottom_out[1]
rlabel metal1 27232 37094 27232 37094 0 chany_bottom_out[2]
rlabel metal1 28520 37094 28520 37094 0 chany_bottom_out[3]
rlabel metal2 34178 1520 34178 1520 0 chany_bottom_out[4]
rlabel metal1 20148 37094 20148 37094 0 chany_bottom_out[5]
rlabel via2 38226 33371 38226 33371 0 chany_bottom_out[6]
rlabel metal2 23874 1520 23874 1520 0 chany_bottom_out[7]
rlabel metal3 1188 21148 1188 21148 0 chany_bottom_out[8]
rlabel metal1 37030 2278 37030 2278 0 chany_bottom_out[9]
rlabel metal2 38226 15895 38226 15895 0 chany_top_in[0]
rlabel metal1 2346 36754 2346 36754 0 chany_top_in[10]
rlabel via2 1610 10251 1610 10251 0 chany_top_in[11]
rlabel via2 1610 32011 1610 32011 0 chany_top_in[12]
rlabel metal3 1142 6868 1142 6868 0 chany_top_in[13]
rlabel metal2 38318 37383 38318 37383 0 chany_top_in[14]
rlabel metal1 7866 37230 7866 37230 0 chany_top_in[15]
rlabel metal1 3312 2414 3312 2414 0 chany_top_in[16]
rlabel metal2 9706 1367 9706 1367 0 chany_top_in[17]
rlabel metal1 33764 2414 33764 2414 0 chany_top_in[18]
rlabel metal2 38226 13787 38226 13787 0 chany_top_in[1]
rlabel metal2 38226 6239 38226 6239 0 chany_top_in[2]
rlabel metal2 34086 2924 34086 2924 0 chany_top_in[3]
rlabel metal1 2668 36822 2668 36822 0 chany_top_in[4]
rlabel metal1 38778 3434 38778 3434 0 chany_top_in[5]
rlabel via2 1610 8925 1610 8925 0 chany_top_in[6]
rlabel metal2 38226 10455 38226 10455 0 chany_top_in[7]
rlabel via2 1610 25245 1610 25245 0 chany_top_in[8]
rlabel metal2 32338 2074 32338 2074 0 chany_top_in[9]
rlabel via2 38226 24565 38226 24565 0 chany_top_out[0]
rlabel metal1 11730 37094 11730 37094 0 chany_top_out[10]
rlabel metal1 6578 37094 6578 37094 0 chany_top_out[11]
rlabel metal1 19182 3366 19182 3366 0 chany_top_out[12]
rlabel metal2 46 1656 46 1656 0 chany_top_out[13]
rlabel metal2 21942 2064 21942 2064 0 chany_top_out[14]
rlabel metal1 13018 37094 13018 37094 0 chany_top_out[15]
rlabel metal1 23368 37094 23368 37094 0 chany_top_out[16]
rlabel metal1 33672 37094 33672 37094 0 chany_top_out[17]
rlabel metal3 1188 26588 1188 26588 0 chany_top_out[18]
rlabel metal2 4554 1520 4554 1520 0 chany_top_out[1]
rlabel metal2 1334 1520 1334 1520 0 chany_top_out[2]
rlabel metal1 38456 36346 38456 36346 0 chany_top_out[3]
rlabel metal1 30498 37094 30498 37094 0 chany_top_out[4]
rlabel metal2 16790 823 16790 823 0 chany_top_out[5]
rlabel metal1 37352 36346 37352 36346 0 chany_top_out[6]
rlabel via2 38226 2805 38226 2805 0 chany_top_out[7]
rlabel metal1 4692 37094 4692 37094 0 chany_top_out[8]
rlabel metal2 38226 21233 38226 21233 0 chany_top_out[9]
rlabel metal2 6486 1520 6486 1520 0 left_grid_right_width_0_height_0_subtile_0__pin_I_1_
rlabel metal1 11362 2822 11362 2822 0 left_grid_right_width_0_height_0_subtile_0__pin_I_5_
rlabel metal3 1188 15708 1188 15708 0 left_grid_right_width_0_height_0_subtile_0__pin_I_9_
rlabel metal2 21482 2176 21482 2176 0 mem_left_ipin_0.DFFR_0_.Q
rlabel via2 12558 13685 12558 13685 0 mem_left_ipin_0.DFFR_1_.Q
rlabel metal1 12604 15470 12604 15470 0 mem_left_ipin_0.DFFR_2_.Q
rlabel via2 14674 4437 14674 4437 0 mem_left_ipin_0.DFFR_3_.Q
rlabel metal1 14066 2618 14066 2618 0 mem_left_ipin_0.DFFR_4_.Q
rlabel metal1 13846 2278 13846 2278 0 mem_left_ipin_0.DFFR_5_.Q
rlabel metal2 20608 8772 20608 8772 0 mem_left_ipin_1.DFFR_0_.Q
rlabel metal1 14628 8874 14628 8874 0 mem_left_ipin_1.DFFR_1_.Q
rlabel metal2 19366 8942 19366 8942 0 mem_left_ipin_1.DFFR_2_.Q
rlabel metal2 23782 6426 23782 6426 0 mem_left_ipin_1.DFFR_3_.Q
rlabel metal1 26266 2346 26266 2346 0 mem_left_ipin_1.DFFR_4_.Q
rlabel metal1 24058 2550 24058 2550 0 mem_left_ipin_1.DFFR_5_.Q
rlabel metal1 21896 7786 21896 7786 0 mem_left_ipin_2.DFFR_0_.Q
rlabel metal1 20332 9486 20332 9486 0 mem_left_ipin_2.DFFR_1_.Q
rlabel metal1 15364 17646 15364 17646 0 mem_left_ipin_2.DFFR_2_.Q
rlabel metal2 15226 5916 15226 5916 0 mem_left_ipin_2.DFFR_3_.Q
rlabel metal2 16698 5933 16698 5933 0 mem_left_ipin_2.DFFR_4_.Q
rlabel metal1 21390 6834 21390 6834 0 mem_left_ipin_2.DFFR_5_.Q
rlabel metal1 21712 9962 21712 9962 0 mem_left_ipin_3.DFFR_0_.Q
rlabel metal2 21574 16388 21574 16388 0 mem_left_ipin_3.DFFR_1_.Q
rlabel metal2 19274 13005 19274 13005 0 mem_left_ipin_3.DFFR_2_.Q
rlabel metal1 19366 6664 19366 6664 0 mem_left_ipin_3.DFFR_3_.Q
rlabel metal1 19412 2278 19412 2278 0 mem_left_ipin_3.DFFR_4_.Q
rlabel metal1 17526 7344 17526 7344 0 mem_left_ipin_3.DFFR_5_.Q
rlabel metal1 21298 18326 21298 18326 0 mem_left_ipin_4.DFFR_0_.Q
rlabel metal2 21390 14790 21390 14790 0 mem_left_ipin_4.DFFR_1_.Q
rlabel metal1 23828 7514 23828 7514 0 mem_left_ipin_4.DFFR_2_.Q
rlabel metal2 24518 5474 24518 5474 0 mem_left_ipin_4.DFFR_3_.Q
rlabel metal1 23368 2482 23368 2482 0 mem_left_ipin_4.DFFR_4_.Q
rlabel metal1 23966 2958 23966 2958 0 mem_left_ipin_4.DFFR_5_.Q
rlabel metal1 19826 17646 19826 17646 0 mem_left_ipin_5.DFFR_0_.Q
rlabel metal1 16698 16524 16698 16524 0 mem_left_ipin_5.DFFR_1_.Q
rlabel metal1 21160 7718 21160 7718 0 mem_left_ipin_5.DFFR_2_.Q
rlabel metal1 13524 2346 13524 2346 0 mem_left_ipin_5.DFFR_3_.Q
rlabel metal1 11362 10506 11362 10506 0 mem_left_ipin_5.DFFR_4_.Q
rlabel metal1 15824 6698 15824 6698 0 mem_left_ipin_5.DFFR_5_.Q
rlabel metal1 17296 8874 17296 8874 0 mem_left_ipin_6.DFFR_0_.Q
rlabel metal1 10304 14994 10304 14994 0 mem_left_ipin_6.DFFR_1_.Q
rlabel metal1 15272 8058 15272 8058 0 mem_left_ipin_6.DFFR_2_.Q
rlabel metal1 13616 5610 13616 5610 0 mem_left_ipin_6.DFFR_3_.Q
rlabel metal1 11776 5542 11776 5542 0 mem_left_ipin_6.DFFR_4_.Q
rlabel metal1 13156 9690 13156 9690 0 mem_left_ipin_6.DFFR_5_.Q
rlabel metal1 17158 16626 17158 16626 0 mem_left_ipin_7.DFFR_0_.Q
rlabel metal1 16514 9486 16514 9486 0 mem_left_ipin_7.DFFR_1_.Q
rlabel metal1 18538 17646 18538 17646 0 mem_left_ipin_7.DFFR_2_.Q
rlabel metal2 21390 7616 21390 7616 0 mem_left_ipin_7.DFFR_3_.Q
rlabel metal1 16882 3366 16882 3366 0 mem_left_ipin_7.DFFR_4_.Q
rlabel metal1 20194 13498 20194 13498 0 mem_left_ipin_7.DFFR_5_.Q
rlabel metal2 19642 6885 19642 6885 0 mem_right_ipin_0.DFFR_0_.Q
rlabel metal2 18722 14212 18722 14212 0 mem_right_ipin_0.DFFR_1_.Q
rlabel metal1 14398 3094 14398 3094 0 mem_right_ipin_0.DFFR_2_.Q
rlabel metal1 14582 3162 14582 3162 0 mem_right_ipin_0.DFFR_3_.Q
rlabel metal2 17434 4403 17434 4403 0 mem_right_ipin_0.DFFR_4_.Q
rlabel metal1 18538 5746 18538 5746 0 mem_right_ipin_0.DFFR_5_.Q
rlabel metal1 14168 14382 14168 14382 0 mem_right_ipin_1.DFFR_0_.Q
rlabel metal1 18630 17204 18630 17204 0 mem_right_ipin_1.DFFR_1_.Q
rlabel metal1 21965 5610 21965 5610 0 mem_right_ipin_1.DFFR_2_.Q
rlabel metal3 25070 12852 25070 12852 0 mem_right_ipin_1.DFFR_3_.Q
rlabel metal1 18630 4760 18630 4760 0 mem_right_ipin_1.DFFR_4_.Q
rlabel metal1 20746 8466 20746 8466 0 mem_right_ipin_1.DFFR_5_.Q
rlabel metal1 21528 10778 21528 10778 0 mem_right_ipin_2.DFFR_0_.Q
rlabel metal2 14950 17119 14950 17119 0 mem_right_ipin_2.DFFR_1_.Q
rlabel metal1 15916 18258 15916 18258 0 mem_right_ipin_2.DFFR_2_.Q
rlabel metal1 12696 10438 12696 10438 0 mem_right_ipin_2.DFFR_3_.Q
rlabel metal1 14122 8602 14122 8602 0 mem_right_ipin_2.DFFR_4_.Q
rlabel metal1 19734 13362 19734 13362 0 mux_left_ipin_0.INVTX1_0_.out
rlabel metal1 17894 9622 17894 9622 0 mux_left_ipin_0.INVTX1_1_.out
rlabel metal1 14582 22406 14582 22406 0 mux_left_ipin_0.INVTX1_2_.out
rlabel metal1 12926 9962 12926 9962 0 mux_left_ipin_0.INVTX1_3_.out
rlabel metal2 12466 15130 12466 15130 0 mux_left_ipin_0.INVTX1_4_.out
rlabel metal1 13294 25126 13294 25126 0 mux_left_ipin_0.INVTX1_5_.out
rlabel via2 13294 10557 13294 10557 0 mux_left_ipin_0.INVTX1_6_.out
rlabel metal1 28244 3366 28244 3366 0 mux_left_ipin_0.INVTX1_7_.out
rlabel metal1 16606 9554 16606 9554 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 13570 15504 13570 15504 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 15042 10472 15042 10472 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 9798 9758 9798 9758 0 mux_left_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 22954 11186 22954 11186 0 mux_left_ipin_1.INVTX1_2_.out
rlabel metal1 20976 11186 20976 11186 0 mux_left_ipin_1.INVTX1_3_.out
rlabel metal1 19688 11050 19688 11050 0 mux_left_ipin_1.INVTX1_4_.out
rlabel metal2 27094 10268 27094 10268 0 mux_left_ipin_1.INVTX1_5_.out
rlabel metal1 11500 14314 11500 14314 0 mux_left_ipin_1.INVTX1_6_.out
rlabel metal1 7912 12954 7912 12954 0 mux_left_ipin_1.INVTX1_7_.out
rlabel metal1 20470 11628 20470 11628 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 27922 10030 27922 10030 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 20654 13549 20654 13549 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 27370 24106 27370 24106 0 mux_left_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 23828 12750 23828 12750 0 mux_left_ipin_2.INVTX1_2_.out
rlabel metal2 26450 15266 26450 15266 0 mux_left_ipin_2.INVTX1_3_.out
rlabel metal2 23138 17612 23138 17612 0 mux_left_ipin_2.INVTX1_4_.out
rlabel metal1 13892 19482 13892 19482 0 mux_left_ipin_2.INVTX1_5_.out
rlabel metal1 15594 12750 15594 12750 0 mux_left_ipin_2.INVTX1_6_.out
rlabel metal1 27784 24038 27784 24038 0 mux_left_ipin_2.INVTX1_7_.out
rlabel metal2 20470 13464 20470 13464 0 mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 23414 15419 23414 15419 0 mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 21574 16694 21574 16694 0 mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 12466 24106 12466 24106 0 mux_left_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 28520 26758 28520 26758 0 mux_left_ipin_3.INVTX1_2_.out
rlabel metal1 26818 14314 26818 14314 0 mux_left_ipin_3.INVTX1_3_.out
rlabel metal2 20010 18972 20010 18972 0 mux_left_ipin_3.INVTX1_4_.out
rlabel metal2 25668 13838 25668 13838 0 mux_left_ipin_3.INVTX1_5_.out
rlabel metal1 20378 16014 20378 16014 0 mux_left_ipin_3.INVTX1_6_.out
rlabel viali 15686 16008 15686 16008 0 mux_left_ipin_3.INVTX1_7_.out
rlabel metal2 23506 13022 23506 13022 0 mux_left_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 23046 14892 23046 14892 0 mux_left_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 20470 17374 20470 17374 0 mux_left_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 14858 28050 14858 28050 0 mux_left_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 26542 25126 26542 25126 0 mux_left_ipin_4.INVTX1_2_.out
rlabel metal2 19918 17204 19918 17204 0 mux_left_ipin_4.INVTX1_3_.out
rlabel metal2 24794 15538 24794 15538 0 mux_left_ipin_4.INVTX1_4_.out
rlabel metal1 16606 25194 16606 25194 0 mux_left_ipin_4.INVTX1_5_.out
rlabel metal1 22218 28390 22218 28390 0 mux_left_ipin_4.INVTX1_6_.out
rlabel metal2 16928 16014 16928 16014 0 mux_left_ipin_4.INVTX1_7_.out
rlabel metal1 27738 13226 27738 13226 0 mux_left_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 19366 16048 19366 16048 0 mux_left_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel via2 19182 13821 19182 13821 0 mux_left_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 30590 6562 30590 6562 0 mux_left_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 25622 9316 25622 9316 0 mux_left_ipin_5.INVTX1_2_.out
rlabel metal1 22954 12716 22954 12716 0 mux_left_ipin_5.INVTX1_3_.out
rlabel metal1 13846 28390 13846 28390 0 mux_left_ipin_5.INVTX1_4_.out
rlabel metal1 10396 10506 10396 10506 0 mux_left_ipin_5.INVTX1_5_.out
rlabel metal1 20378 29002 20378 29002 0 mux_left_ipin_5.INVTX1_6_.out
rlabel metal1 12006 3162 12006 3162 0 mux_left_ipin_5.INVTX1_7_.out
rlabel metal2 15962 17442 15962 17442 0 mux_left_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel via2 22310 12733 22310 12733 0 mux_left_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 12466 13311 12466 13311 0 mux_left_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 12742 9418 12742 9418 0 mux_left_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 16054 16218 16054 16218 0 mux_left_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 13616 13838 13616 13838 0 mux_left_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 15778 11662 15778 11662 0 mux_left_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 3128 35462 3128 35462 0 mux_left_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 19044 15062 19044 15062 0 mux_left_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 17894 11373 17894 11373 0 mux_left_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 16284 13906 16284 13906 0 mux_left_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 26680 13294 26680 13294 0 mux_left_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 22724 11050 22724 11050 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 24656 13974 24656 13974 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 21758 13719 21758 13719 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 14766 13532 14766 13532 0 mux_right_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 24978 14144 24978 14144 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 18124 12750 18124 12750 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 18814 16082 18814 16082 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 18676 12750 18676 12750 0 mux_right_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 16974 15470 16974 15470 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 17526 14450 17526 14450 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 19182 19210 19182 19210 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 15732 15606 15732 15606 0 mux_right_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 1794 3400 1794 3400 0 net1
rlabel metal1 21436 37230 21436 37230 0 net10
rlabel metal1 19550 12954 19550 12954 0 net100
rlabel metal2 19458 20638 19458 20638 0 net101
rlabel metal1 10856 2550 10856 2550 0 net11
rlabel metal2 18170 8704 18170 8704 0 net12
rlabel metal1 36984 17034 36984 17034 0 net13
rlabel metal1 37352 36686 37352 36686 0 net14
rlabel metal1 29072 25466 29072 25466 0 net15
rlabel metal2 38042 4896 38042 4896 0 net16
rlabel metal1 15088 22610 15088 22610 0 net17
rlabel metal2 9338 1972 9338 1972 0 net18
rlabel metal1 23184 26758 23184 26758 0 net19
rlabel metal2 1794 18598 1794 18598 0 net2
rlabel metal2 1886 23868 1886 23868 0 net20
rlabel via2 38042 15963 38042 15963 0 net21
rlabel metal1 16238 25262 16238 25262 0 net22
rlabel metal1 14030 5304 14030 5304 0 net23
rlabel metal1 20056 35054 20056 35054 0 net24
rlabel metal1 2576 19822 2576 19822 0 net25
rlabel metal1 37950 37230 37950 37230 0 net26
rlabel metal1 11684 16082 11684 16082 0 net27
rlabel metal1 2714 2618 2714 2618 0 net28
rlabel metal1 7682 3094 7682 3094 0 net29
rlabel metal1 33304 2550 33304 2550 0 net3
rlabel metal2 31326 2516 31326 2516 0 net30
rlabel metal1 19872 16490 19872 16490 0 net31
rlabel metal1 26036 21522 26036 21522 0 net32
rlabel metal1 28658 30566 28658 30566 0 net33
rlabel metal2 2530 28016 2530 28016 0 net34
rlabel metal1 37996 3638 37996 3638 0 net35
rlabel metal1 12535 19346 12535 19346 0 net36
rlabel metal2 37030 10064 37030 10064 0 net37
rlabel metal1 2024 20910 2024 20910 0 net38
rlabel metal1 32844 2278 32844 2278 0 net39
rlabel metal1 14306 37230 14306 37230 0 net4
rlabel metal1 37996 22474 37996 22474 0 net40
rlabel metal1 37996 36754 37996 36754 0 net41
rlabel metal1 1886 14450 1886 14450 0 net42
rlabel metal1 37766 28050 37766 28050 0 net43
rlabel metal2 37490 2244 37490 2244 0 net44
rlabel metal1 23000 37162 23000 37162 0 net45
rlabel metal1 2116 37230 2116 37230 0 net46
rlabel metal2 38042 30022 38042 30022 0 net47
rlabel metal1 1886 19788 1886 19788 0 net48
rlabel metal1 1932 19482 1932 19482 0 net49
rlabel metal1 16974 37298 16974 37298 0 net5
rlabel metal1 1886 2992 1886 2992 0 net50
rlabel metal1 30912 2414 30912 2414 0 net51
rlabel metal1 2300 34510 2300 34510 0 net52
rlabel metal1 26542 37230 26542 37230 0 net53
rlabel metal1 27968 37230 27968 37230 0 net54
rlabel metal1 34868 3706 34868 3706 0 net55
rlabel metal2 20056 26220 20056 26220 0 net56
rlabel metal1 37766 33490 37766 33490 0 net57
rlabel metal1 27692 2414 27692 2414 0 net58
rlabel metal2 1794 21318 1794 21318 0 net59
rlabel metal2 12558 15895 12558 15895 0 net6
rlabel metal2 36662 2652 36662 2652 0 net60
rlabel metal1 37812 24786 37812 24786 0 net61
rlabel metal1 12052 37230 12052 37230 0 net62
rlabel metal1 8878 36550 8878 36550 0 net63
rlabel metal1 18998 3502 18998 3502 0 net64
rlabel metal1 2760 2414 2760 2414 0 net65
rlabel via2 32982 3587 32982 3587 0 net66
rlabel metal1 16100 26010 16100 26010 0 net67
rlabel metal1 22770 36890 22770 36890 0 net68
rlabel metal1 30820 36890 30820 36890 0 net69
rlabel via2 12650 3723 12650 3723 0 net7
rlabel metal1 4232 26962 4232 26962 0 net70
rlabel metal1 4922 2448 4922 2448 0 net71
rlabel metal1 1886 2448 1886 2448 0 net72
rlabel metal2 38042 36346 38042 36346 0 net73
rlabel metal1 30452 37230 30452 37230 0 net74
rlabel metal2 20470 3162 20470 3162 0 net75
rlabel metal1 37030 36142 37030 36142 0 net76
rlabel metal2 38042 3502 38042 3502 0 net77
rlabel metal2 5474 36992 5474 36992 0 net78
rlabel metal2 37490 19992 37490 19992 0 net79
rlabel metal1 18676 25874 18676 25874 0 net8
rlabel metal1 7544 2414 7544 2414 0 net80
rlabel metal1 10166 3026 10166 3026 0 net81
rlabel metal2 8142 15878 8142 15878 0 net82
rlabel metal2 2806 6766 2806 6766 0 net83
rlabel metal1 31602 37230 31602 37230 0 net84
rlabel metal1 4876 37162 4876 37162 0 net85
rlabel metal1 11638 37162 11638 37162 0 net86
rlabel metal2 27462 3502 27462 3502 0 net87
rlabel metal1 3726 12818 3726 12818 0 net88
rlabel metal1 2024 35802 2024 35802 0 net89
rlabel metal2 22770 36448 22770 36448 0 net9
rlabel metal1 37352 19346 37352 19346 0 net90
rlabel metal2 14030 10132 14030 10132 0 net91
rlabel metal1 10994 13294 10994 13294 0 net92
rlabel metal1 20010 15538 20010 15538 0 net93
rlabel metal1 20746 18666 20746 18666 0 net94
rlabel metal2 23414 16762 23414 16762 0 net95
rlabel metal1 11730 12886 11730 12886 0 net96
rlabel metal2 12282 11492 12282 11492 0 net97
rlabel via2 12466 14059 12466 14059 0 net98
rlabel metal1 15686 11832 15686 11832 0 net99
rlabel metal2 38226 22559 38226 22559 0 pReset
rlabel metal1 19458 2380 19458 2380 0 prog_clk
rlabel metal3 1188 4828 1188 4828 0 right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 32384 37094 32384 37094 0 right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal2 2806 37145 2806 37145 0 right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 9798 37094 9798 37094 0 right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 27186 2822 27186 2822 0 right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_
rlabel metal3 1188 12308 1188 12308 0 right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_
rlabel metal3 1188 36108 1188 36108 0 right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_
rlabel via2 38226 19125 38226 19125 0 right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
