magic
tech sky130A
magscale 1 2
timestamp 1672417756
<< viali >>
rect 1777 37417 1811 37451
rect 18889 37281 18923 37315
rect 22017 37281 22051 37315
rect 27445 37281 27479 37315
rect 1593 37213 1627 37247
rect 2881 37213 2915 37247
rect 3985 37213 4019 37247
rect 4905 37213 4939 37247
rect 6009 37213 6043 37247
rect 6745 37213 6779 37247
rect 7849 37213 7883 37247
rect 9781 37213 9815 37247
rect 11713 37213 11747 37247
rect 12633 37213 12667 37247
rect 13737 37213 13771 37247
rect 14289 37213 14323 37247
rect 15577 37213 15611 37247
rect 17509 37213 17543 37247
rect 18705 37213 18739 37247
rect 20085 37213 20119 37247
rect 22293 37213 22327 37247
rect 24593 37213 24627 37247
rect 25513 37213 25547 37247
rect 27261 37213 27295 37247
rect 27905 37213 27939 37247
rect 28825 37213 28859 37247
rect 29929 37213 29963 37247
rect 31217 37213 31251 37247
rect 32321 37213 32355 37247
rect 33057 37213 33091 37247
rect 34897 37213 34931 37247
rect 35449 37213 35483 37247
rect 35817 37213 35851 37247
rect 36277 37213 36311 37247
rect 37565 37213 37599 37247
rect 2697 37077 2731 37111
rect 4169 37077 4203 37111
rect 4721 37077 4755 37111
rect 5825 37077 5859 37111
rect 6561 37077 6595 37111
rect 8033 37077 8067 37111
rect 9965 37077 9999 37111
rect 11897 37077 11931 37111
rect 12449 37077 12483 37111
rect 13553 37077 13587 37111
rect 14473 37077 14507 37111
rect 15761 37077 15795 37111
rect 17693 37077 17727 37111
rect 20269 37077 20303 37111
rect 24777 37077 24811 37111
rect 25329 37077 25363 37111
rect 28089 37077 28123 37111
rect 28641 37077 28675 37111
rect 29745 37077 29779 37111
rect 31033 37077 31067 37111
rect 32505 37077 32539 37111
rect 33241 37077 33275 37111
rect 35081 37077 35115 37111
rect 36369 37077 36403 37111
rect 37657 37077 37691 37111
rect 1777 36873 1811 36907
rect 9321 36873 9355 36907
rect 14841 36873 14875 36907
rect 17049 36873 17083 36907
rect 27169 36873 27203 36907
rect 38117 36805 38151 36839
rect 1593 36737 1627 36771
rect 2513 36737 2547 36771
rect 3157 36737 3191 36771
rect 9137 36737 9171 36771
rect 14105 36737 14139 36771
rect 14197 36737 14231 36771
rect 15025 36737 15059 36771
rect 16865 36737 16899 36771
rect 17877 36737 17911 36771
rect 22201 36737 22235 36771
rect 23305 36737 23339 36771
rect 27353 36737 27387 36771
rect 35725 36737 35759 36771
rect 36921 36737 36955 36771
rect 23581 36669 23615 36703
rect 17693 36601 17727 36635
rect 36737 36601 36771 36635
rect 38301 36601 38335 36635
rect 2329 36533 2363 36567
rect 2973 36533 3007 36567
rect 22017 36533 22051 36567
rect 35541 36533 35575 36567
rect 19717 36329 19751 36363
rect 37473 36329 37507 36363
rect 1777 36125 1811 36159
rect 19901 36125 19935 36159
rect 37289 36125 37323 36159
rect 38025 36125 38059 36159
rect 1593 35989 1627 36023
rect 38209 35989 38243 36023
rect 38117 35649 38151 35683
rect 1593 35581 1627 35615
rect 1869 35581 1903 35615
rect 38209 35445 38243 35479
rect 3157 35241 3191 35275
rect 19533 35241 19567 35275
rect 1777 35037 1811 35071
rect 3341 35037 3375 35071
rect 19441 35037 19475 35071
rect 38301 35037 38335 35071
rect 1593 34901 1627 34935
rect 38117 34901 38151 34935
rect 4353 34697 4387 34731
rect 4537 34561 4571 34595
rect 38025 34561 38059 34595
rect 38209 34357 38243 34391
rect 22017 34153 22051 34187
rect 22201 33949 22235 33983
rect 1593 33473 1627 33507
rect 8585 33473 8619 33507
rect 1777 33337 1811 33371
rect 8677 33269 8711 33303
rect 33241 33065 33275 33099
rect 9597 32861 9631 32895
rect 11069 32861 11103 32895
rect 28273 32861 28307 32895
rect 33425 32861 33459 32895
rect 38117 32793 38151 32827
rect 9689 32725 9723 32759
rect 11161 32725 11195 32759
rect 28365 32725 28399 32759
rect 38209 32725 38243 32759
rect 9045 32521 9079 32555
rect 10609 32521 10643 32555
rect 1593 32385 1627 32419
rect 9229 32385 9263 32419
rect 10793 32385 10827 32419
rect 20729 32385 20763 32419
rect 23489 32385 23523 32419
rect 38117 32385 38151 32419
rect 1777 32181 1811 32215
rect 2237 32181 2271 32215
rect 20821 32181 20855 32215
rect 23581 32181 23615 32215
rect 38209 32181 38243 32215
rect 24685 31977 24719 32011
rect 1869 31841 1903 31875
rect 21465 31841 21499 31875
rect 28089 31841 28123 31875
rect 1593 31773 1627 31807
rect 21373 31773 21407 31807
rect 24593 31773 24627 31807
rect 27997 31773 28031 31807
rect 29285 31297 29319 31331
rect 29377 31093 29411 31127
rect 8401 30889 8435 30923
rect 25973 30889 26007 30923
rect 5917 30821 5951 30855
rect 37749 30753 37783 30787
rect 3985 30685 4019 30719
rect 5825 30685 5859 30719
rect 6469 30685 6503 30719
rect 7113 30685 7147 30719
rect 8309 30685 8343 30719
rect 9689 30685 9723 30719
rect 12909 30685 12943 30719
rect 26157 30685 26191 30719
rect 27997 30685 28031 30719
rect 37473 30685 37507 30719
rect 7205 30617 7239 30651
rect 4077 30549 4111 30583
rect 6561 30549 6595 30583
rect 9781 30549 9815 30583
rect 13001 30549 13035 30583
rect 28089 30549 28123 30583
rect 1593 30209 1627 30243
rect 4353 30209 4387 30243
rect 1777 30005 1811 30039
rect 4445 30005 4479 30039
rect 4905 29801 4939 29835
rect 27445 29801 27479 29835
rect 1777 29597 1811 29631
rect 5089 29597 5123 29631
rect 9137 29597 9171 29631
rect 11805 29597 11839 29631
rect 17877 29597 17911 29631
rect 27353 29597 27387 29631
rect 38025 29597 38059 29631
rect 9229 29529 9263 29563
rect 1593 29461 1627 29495
rect 11621 29461 11655 29495
rect 17693 29461 17727 29495
rect 38209 29461 38243 29495
rect 8217 29257 8251 29291
rect 16865 29257 16899 29291
rect 1777 29121 1811 29155
rect 8125 29121 8159 29155
rect 11897 29121 11931 29155
rect 17049 29121 17083 29155
rect 17693 29121 17727 29155
rect 1593 28985 1627 29019
rect 11713 28985 11747 29019
rect 17509 28917 17543 28951
rect 17233 28645 17267 28679
rect 17049 28577 17083 28611
rect 1869 28509 1903 28543
rect 2513 28509 2547 28543
rect 16221 28509 16255 28543
rect 16865 28509 16899 28543
rect 1961 28441 1995 28475
rect 2605 28373 2639 28407
rect 16313 28373 16347 28407
rect 5825 28169 5859 28203
rect 16957 28169 16991 28203
rect 21373 28169 21407 28203
rect 1961 28033 1995 28067
rect 2605 28033 2639 28067
rect 3433 28033 3467 28067
rect 4077 28033 4111 28067
rect 5733 28033 5767 28067
rect 8309 28033 8343 28067
rect 8953 28033 8987 28067
rect 12633 28033 12667 28067
rect 17693 28033 17727 28067
rect 19257 28033 19291 28067
rect 21281 28033 21315 28067
rect 10425 27965 10459 27999
rect 10609 27965 10643 27999
rect 12725 27965 12759 27999
rect 37473 27965 37507 27999
rect 37749 27965 37783 27999
rect 2697 27897 2731 27931
rect 8125 27897 8159 27931
rect 2053 27829 2087 27863
rect 3249 27829 3283 27863
rect 3893 27829 3927 27863
rect 8769 27829 8803 27863
rect 11069 27829 11103 27863
rect 17785 27829 17819 27863
rect 19073 27829 19107 27863
rect 18705 27625 18739 27659
rect 11069 27557 11103 27591
rect 17325 27557 17359 27591
rect 37381 27557 37415 27591
rect 10425 27489 10459 27523
rect 10609 27489 10643 27523
rect 17141 27489 17175 27523
rect 1869 27421 1903 27455
rect 2513 27421 2547 27455
rect 3157 27421 3191 27455
rect 3985 27421 4019 27455
rect 7757 27421 7791 27455
rect 9965 27421 9999 27455
rect 13001 27421 13035 27455
rect 16957 27421 16991 27455
rect 18061 27421 18095 27455
rect 18889 27421 18923 27455
rect 19441 27421 19475 27455
rect 22109 27421 22143 27455
rect 37565 27421 37599 27455
rect 38025 27421 38059 27455
rect 1961 27285 1995 27319
rect 2605 27285 2639 27319
rect 3249 27285 3283 27319
rect 7849 27285 7883 27319
rect 9781 27285 9815 27319
rect 12817 27285 12851 27319
rect 18153 27285 18187 27319
rect 19533 27285 19567 27319
rect 22201 27285 22235 27319
rect 38209 27285 38243 27319
rect 5181 27081 5215 27115
rect 37565 27081 37599 27115
rect 12725 27013 12759 27047
rect 17049 27013 17083 27047
rect 17601 27013 17635 27047
rect 1869 26945 1903 26979
rect 2513 26945 2547 26979
rect 3801 26945 3835 26979
rect 4445 26945 4479 26979
rect 5365 26945 5399 26979
rect 7113 26945 7147 26979
rect 11897 26945 11931 26979
rect 18797 26945 18831 26979
rect 37473 26945 37507 26979
rect 3157 26877 3191 26911
rect 12633 26877 12667 26911
rect 12909 26877 12943 26911
rect 16957 26877 16991 26911
rect 18981 26877 19015 26911
rect 2605 26809 2639 26843
rect 1961 26741 1995 26775
rect 3893 26741 3927 26775
rect 4537 26741 4571 26775
rect 7205 26741 7239 26775
rect 11989 26741 12023 26775
rect 19349 26741 19383 26775
rect 8309 26537 8343 26571
rect 13185 26537 13219 26571
rect 5825 26469 5859 26503
rect 7021 26469 7055 26503
rect 14473 26469 14507 26503
rect 15945 26469 15979 26503
rect 38117 26469 38151 26503
rect 3249 26401 3283 26435
rect 7849 26401 7883 26435
rect 12081 26401 12115 26435
rect 12449 26401 12483 26435
rect 20637 26401 20671 26435
rect 20913 26401 20947 26435
rect 1869 26333 1903 26367
rect 2513 26333 2547 26367
rect 3157 26333 3191 26367
rect 4077 26333 4111 26367
rect 5181 26333 5215 26367
rect 5273 26333 5307 26367
rect 6009 26333 6043 26367
rect 6929 26333 6963 26367
rect 7665 26333 7699 26367
rect 13369 26333 13403 26367
rect 14381 26333 14415 26367
rect 16129 26333 16163 26367
rect 16773 26333 16807 26367
rect 38301 26333 38335 26367
rect 1961 26265 1995 26299
rect 2605 26265 2639 26299
rect 4169 26265 4203 26299
rect 12173 26265 12207 26299
rect 20729 26265 20763 26299
rect 16589 26197 16623 26231
rect 17785 26197 17819 26231
rect 7849 25993 7883 26027
rect 13369 25993 13403 26027
rect 17785 25925 17819 25959
rect 17877 25925 17911 25959
rect 2145 25857 2179 25891
rect 3249 25857 3283 25891
rect 4169 25857 4203 25891
rect 4813 25857 4847 25891
rect 5641 25857 5675 25891
rect 6561 25857 6595 25891
rect 7757 25857 7791 25891
rect 10977 25857 11011 25891
rect 13553 25857 13587 25891
rect 14013 25857 14047 25891
rect 14657 25857 14691 25891
rect 15485 25857 15519 25891
rect 6653 25789 6687 25823
rect 9689 25789 9723 25823
rect 9873 25789 9907 25823
rect 16865 25789 16899 25823
rect 18061 25789 18095 25823
rect 4905 25721 4939 25755
rect 10793 25721 10827 25755
rect 2237 25653 2271 25687
rect 3341 25653 3375 25687
rect 4261 25653 4295 25687
rect 5733 25653 5767 25687
rect 10057 25653 10091 25687
rect 14105 25653 14139 25687
rect 14749 25653 14783 25687
rect 15301 25653 15335 25687
rect 10701 25449 10735 25483
rect 20085 25449 20119 25483
rect 29929 25449 29963 25483
rect 5365 25381 5399 25415
rect 6193 25313 6227 25347
rect 13645 25313 13679 25347
rect 16313 25313 16347 25347
rect 16957 25313 16991 25347
rect 1593 25245 1627 25279
rect 2329 25245 2363 25279
rect 4537 25245 4571 25279
rect 5549 25245 5583 25279
rect 6009 25245 6043 25279
rect 7113 25245 7147 25279
rect 9137 25245 9171 25279
rect 10885 25245 10919 25279
rect 15117 25245 15151 25279
rect 15577 25245 15611 25279
rect 18705 25245 18739 25279
rect 19993 25245 20027 25279
rect 21465 25245 21499 25279
rect 30113 25245 30147 25279
rect 6653 25177 6687 25211
rect 9229 25177 9263 25211
rect 12265 25177 12299 25211
rect 13001 25177 13035 25211
rect 13093 25177 13127 25211
rect 16405 25177 16439 25211
rect 1777 25109 1811 25143
rect 2421 25109 2455 25143
rect 2973 25109 3007 25143
rect 4629 25109 4663 25143
rect 7205 25109 7239 25143
rect 8125 25109 8159 25143
rect 14289 25109 14323 25143
rect 14933 25109 14967 25143
rect 15669 25109 15703 25143
rect 18797 25109 18831 25143
rect 21557 25109 21591 25143
rect 4721 24837 4755 24871
rect 13461 24837 13495 24871
rect 15209 24837 15243 24871
rect 17969 24837 18003 24871
rect 1961 24769 1995 24803
rect 3341 24769 3375 24803
rect 3985 24769 4019 24803
rect 4629 24769 4663 24803
rect 5273 24769 5307 24803
rect 8033 24769 8067 24803
rect 8217 24769 8251 24803
rect 9321 24769 9355 24803
rect 10057 24769 10091 24803
rect 15761 24769 15795 24803
rect 17049 24769 17083 24803
rect 38025 24769 38059 24803
rect 2513 24701 2547 24735
rect 5365 24701 5399 24735
rect 7021 24701 7055 24735
rect 13369 24701 13403 24735
rect 14381 24701 14415 24735
rect 15117 24701 15151 24735
rect 17877 24701 17911 24735
rect 18705 24701 18739 24735
rect 8401 24633 8435 24667
rect 1777 24565 1811 24599
rect 3433 24565 3467 24599
rect 4077 24565 4111 24599
rect 9137 24565 9171 24599
rect 9873 24565 9907 24599
rect 16865 24565 16899 24599
rect 38209 24565 38243 24599
rect 5917 24361 5951 24395
rect 9137 24361 9171 24395
rect 19441 24361 19475 24395
rect 20361 24361 20395 24395
rect 4077 24293 4111 24327
rect 18613 24293 18647 24327
rect 7021 24225 7055 24259
rect 13461 24225 13495 24259
rect 14381 24225 14415 24259
rect 14841 24225 14875 24259
rect 16681 24225 16715 24259
rect 1593 24157 1627 24191
rect 2513 24157 2547 24191
rect 3157 24157 3191 24191
rect 3985 24157 4019 24191
rect 4629 24157 4663 24191
rect 5273 24157 5307 24191
rect 6101 24157 6135 24191
rect 7665 24157 7699 24191
rect 8217 24157 8251 24191
rect 9321 24157 9355 24191
rect 10057 24157 10091 24191
rect 11069 24157 11103 24191
rect 15853 24157 15887 24191
rect 17509 24157 17543 24191
rect 18521 24157 18555 24191
rect 19625 24157 19659 24191
rect 20269 24157 20303 24191
rect 31033 24157 31067 24191
rect 38025 24157 38059 24191
rect 4721 24089 4755 24123
rect 7113 24089 7147 24123
rect 8401 24089 8435 24123
rect 12817 24089 12851 24123
rect 12909 24089 12943 24123
rect 14473 24089 14507 24123
rect 16405 24089 16439 24123
rect 16497 24089 16531 24123
rect 1777 24021 1811 24055
rect 2605 24021 2639 24055
rect 3249 24021 3283 24055
rect 5365 24021 5399 24055
rect 10149 24021 10183 24055
rect 11161 24021 11195 24055
rect 15669 24021 15703 24055
rect 17601 24021 17635 24055
rect 31125 24021 31159 24055
rect 38209 24021 38243 24055
rect 3985 23817 4019 23851
rect 6653 23817 6687 23851
rect 7481 23817 7515 23851
rect 8861 23817 8895 23851
rect 9965 23817 9999 23851
rect 13369 23817 13403 23851
rect 22109 23817 22143 23851
rect 32689 23817 32723 23851
rect 15393 23749 15427 23783
rect 15485 23749 15519 23783
rect 17233 23749 17267 23783
rect 18981 23749 19015 23783
rect 1685 23681 1719 23715
rect 2605 23681 2639 23715
rect 3249 23681 3283 23715
rect 3893 23681 3927 23715
rect 4721 23681 4755 23715
rect 5181 23681 5215 23715
rect 5825 23681 5859 23715
rect 6561 23681 6595 23715
rect 7389 23681 7423 23715
rect 8401 23681 8435 23715
rect 9321 23681 9355 23715
rect 9505 23681 9539 23715
rect 10517 23681 10551 23715
rect 11713 23681 11747 23715
rect 13277 23681 13311 23715
rect 14105 23681 14139 23715
rect 14565 23681 14599 23715
rect 22017 23681 22051 23715
rect 23305 23681 23339 23715
rect 24501 23681 24535 23715
rect 32873 23681 32907 23715
rect 1869 23613 1903 23647
rect 8217 23613 8251 23647
rect 15669 23613 15703 23647
rect 17141 23613 17175 23647
rect 18061 23613 18095 23647
rect 18889 23613 18923 23647
rect 19349 23613 19383 23647
rect 23489 23613 23523 23647
rect 24593 23613 24627 23647
rect 3341 23545 3375 23579
rect 13921 23545 13955 23579
rect 2697 23477 2731 23511
rect 4537 23477 4571 23511
rect 5273 23477 5307 23511
rect 5917 23477 5951 23511
rect 10609 23477 10643 23511
rect 11805 23477 11839 23511
rect 14657 23477 14691 23511
rect 23949 23477 23983 23511
rect 6101 23273 6135 23307
rect 17785 23273 17819 23307
rect 18429 23273 18463 23307
rect 16773 23205 16807 23239
rect 27353 23205 27387 23239
rect 5641 23137 5675 23171
rect 9505 23137 9539 23171
rect 10517 23137 10551 23171
rect 12541 23137 12575 23171
rect 14381 23137 14415 23171
rect 14749 23137 14783 23171
rect 3249 23069 3283 23103
rect 4169 23069 4203 23103
rect 4813 23069 4847 23103
rect 5457 23069 5491 23103
rect 7757 23069 7791 23103
rect 8401 23069 8435 23103
rect 11069 23069 11103 23103
rect 11805 23069 11839 23103
rect 15485 23069 15519 23103
rect 18337 23069 18371 23103
rect 24777 23069 24811 23103
rect 25421 23069 25455 23103
rect 27261 23069 27295 23103
rect 1777 23001 1811 23035
rect 1869 23001 1903 23035
rect 2421 23001 2455 23035
rect 4905 23001 4939 23035
rect 9597 23001 9631 23035
rect 12633 23001 12667 23035
rect 13553 23001 13587 23035
rect 14473 23001 14507 23035
rect 16589 23001 16623 23035
rect 17693 23001 17727 23035
rect 3341 22933 3375 22967
rect 4261 22933 4295 22967
rect 7113 22933 7147 22967
rect 7849 22933 7883 22967
rect 8493 22933 8527 22967
rect 11161 22933 11195 22967
rect 11897 22933 11931 22967
rect 15577 22933 15611 22967
rect 24593 22933 24627 22967
rect 25237 22933 25271 22967
rect 6837 22729 6871 22763
rect 1777 22661 1811 22695
rect 2881 22661 2915 22695
rect 2973 22661 3007 22695
rect 3525 22661 3559 22695
rect 7481 22661 7515 22695
rect 7573 22661 7607 22695
rect 9045 22661 9079 22695
rect 10149 22661 10183 22695
rect 10241 22661 10275 22695
rect 12357 22661 12391 22695
rect 12909 22661 12943 22695
rect 17969 22661 18003 22695
rect 18705 22661 18739 22695
rect 21189 22661 21223 22695
rect 22201 22661 22235 22695
rect 4537 22593 4571 22627
rect 5181 22593 5215 22627
rect 5825 22593 5859 22627
rect 6745 22593 6779 22627
rect 13737 22593 13771 22627
rect 17877 22593 17911 22627
rect 23673 22593 23707 22627
rect 24593 22593 24627 22627
rect 38025 22593 38059 22627
rect 1685 22525 1719 22559
rect 8493 22525 8527 22559
rect 10425 22525 10459 22559
rect 12265 22525 12299 22559
rect 18613 22525 18647 22559
rect 18889 22525 18923 22559
rect 22109 22525 22143 22559
rect 22385 22525 22419 22559
rect 2237 22457 2271 22491
rect 21373 22457 21407 22491
rect 38209 22457 38243 22491
rect 4629 22389 4663 22423
rect 5273 22389 5307 22423
rect 5917 22389 5951 22423
rect 9137 22389 9171 22423
rect 13829 22389 13863 22423
rect 23765 22389 23799 22423
rect 24685 22389 24719 22423
rect 1869 22049 1903 22083
rect 2421 22049 2455 22083
rect 4997 22049 5031 22083
rect 6745 22049 6779 22083
rect 7389 22049 7423 22083
rect 9689 22049 9723 22083
rect 14657 22049 14691 22083
rect 1777 21981 1811 22015
rect 4261 21981 4295 22015
rect 8401 21981 8435 22015
rect 14565 21981 14599 22015
rect 15209 21981 15243 22015
rect 22109 21981 22143 22015
rect 23213 21981 23247 22015
rect 38025 21981 38059 22015
rect 2513 21913 2547 21947
rect 3065 21913 3099 21947
rect 5089 21913 5123 21947
rect 5641 21913 5675 21947
rect 6837 21913 6871 21947
rect 9413 21913 9447 21947
rect 9505 21913 9539 21947
rect 10701 21913 10735 21947
rect 10793 21913 10827 21947
rect 11713 21913 11747 21947
rect 12357 21913 12391 21947
rect 12449 21913 12483 21947
rect 13369 21913 13403 21947
rect 4353 21845 4387 21879
rect 8493 21845 8527 21879
rect 15301 21845 15335 21879
rect 21925 21845 21959 21879
rect 23305 21845 23339 21879
rect 37841 21845 37875 21879
rect 5917 21641 5951 21675
rect 11897 21641 11931 21675
rect 28825 21641 28859 21675
rect 1869 21573 1903 21607
rect 3341 21573 3375 21607
rect 3433 21573 3467 21607
rect 4629 21573 4663 21607
rect 6745 21573 6779 21607
rect 8762 21573 8796 21607
rect 9965 21573 9999 21607
rect 11069 21573 11103 21607
rect 14657 21573 14691 21607
rect 15209 21573 15243 21607
rect 17509 21573 17543 21607
rect 17601 21573 17635 21607
rect 22201 21573 22235 21607
rect 23121 21573 23155 21607
rect 5825 21505 5859 21539
rect 10977 21505 11011 21539
rect 11805 21505 11839 21539
rect 12449 21505 12483 21539
rect 13277 21505 13311 21539
rect 13737 21505 13771 21539
rect 15853 21505 15887 21539
rect 25329 21505 25363 21539
rect 27997 21505 28031 21539
rect 28733 21505 28767 21539
rect 32505 21505 32539 21539
rect 38025 21505 38059 21539
rect 1777 21437 1811 21471
rect 2421 21437 2455 21471
rect 3617 21437 3651 21471
rect 4537 21437 4571 21471
rect 6653 21437 6687 21471
rect 7665 21437 7699 21471
rect 8677 21437 8711 21471
rect 9873 21437 9907 21471
rect 14565 21437 14599 21471
rect 17969 21437 18003 21471
rect 22109 21437 22143 21471
rect 24041 21437 24075 21471
rect 24225 21437 24259 21471
rect 25421 21437 25455 21471
rect 5089 21369 5123 21403
rect 9229 21369 9263 21403
rect 10425 21369 10459 21403
rect 32321 21369 32355 21403
rect 12541 21301 12575 21335
rect 13093 21301 13127 21335
rect 13829 21301 13863 21335
rect 15669 21301 15703 21335
rect 24501 21301 24535 21335
rect 27813 21301 27847 21335
rect 38209 21301 38243 21335
rect 1777 21097 1811 21131
rect 9413 21097 9447 21131
rect 17325 21097 17359 21131
rect 31401 21097 31435 21131
rect 37381 21097 37415 21131
rect 7757 21029 7791 21063
rect 2421 20961 2455 20995
rect 5273 20961 5307 20995
rect 5549 20961 5583 20995
rect 7205 20961 7239 20995
rect 10150 20961 10184 20995
rect 11161 20961 11195 20995
rect 12633 20961 12667 20995
rect 14473 20961 14507 20995
rect 19441 20961 19475 20995
rect 20729 20961 20763 20995
rect 1593 20893 1627 20927
rect 6469 20893 6503 20927
rect 8401 20893 8435 20927
rect 9605 20889 9639 20923
rect 13737 20893 13771 20927
rect 14289 20893 14323 20927
rect 14933 20893 14967 20927
rect 15393 20893 15427 20927
rect 16589 20893 16623 20927
rect 17233 20893 17267 20927
rect 19625 20893 19659 20927
rect 20913 20893 20947 20927
rect 22201 20893 22235 20927
rect 22385 20893 22419 20927
rect 26065 20893 26099 20927
rect 31309 20893 31343 20927
rect 37565 20893 37599 20927
rect 38025 20893 38059 20927
rect 2513 20825 2547 20859
rect 3065 20825 3099 20859
rect 4077 20825 4111 20859
rect 4169 20825 4203 20859
rect 4721 20825 4755 20859
rect 5365 20825 5399 20859
rect 7297 20825 7331 20859
rect 8493 20825 8527 20859
rect 10241 20825 10275 20859
rect 11713 20825 11747 20859
rect 11805 20825 11839 20859
rect 6561 20757 6595 20791
rect 13553 20757 13587 20791
rect 15485 20757 15519 20791
rect 16681 20757 16715 20791
rect 20085 20757 20119 20791
rect 21373 20757 21407 20791
rect 22845 20757 22879 20791
rect 26157 20757 26191 20791
rect 38209 20757 38243 20791
rect 14105 20553 14139 20587
rect 21097 20553 21131 20587
rect 22017 20553 22051 20587
rect 37749 20553 37783 20587
rect 1685 20485 1719 20519
rect 1777 20485 1811 20519
rect 3341 20485 3375 20519
rect 3893 20485 3927 20519
rect 5457 20485 5491 20519
rect 6009 20485 6043 20519
rect 7021 20485 7055 20519
rect 7573 20485 7607 20519
rect 8217 20485 8251 20519
rect 9413 20485 9447 20519
rect 10333 20485 10367 20519
rect 11897 20485 11931 20519
rect 11989 20485 12023 20519
rect 15209 20485 15243 20519
rect 16129 20485 16163 20519
rect 17417 20485 17451 20519
rect 19533 20485 19567 20519
rect 19625 20485 19659 20519
rect 4629 20417 4663 20451
rect 8769 20417 8803 20451
rect 10977 20417 11011 20451
rect 13645 20417 13679 20451
rect 18797 20417 18831 20451
rect 18889 20417 18923 20451
rect 21005 20417 21039 20451
rect 22201 20417 22235 20451
rect 27813 20417 27847 20451
rect 35357 20417 35391 20451
rect 37933 20417 37967 20451
rect 2697 20349 2731 20383
rect 3249 20349 3283 20383
rect 5365 20349 5399 20383
rect 6929 20349 6963 20383
rect 8125 20349 8159 20383
rect 9321 20349 9355 20383
rect 12173 20349 12207 20383
rect 13461 20349 13495 20383
rect 15117 20349 15151 20383
rect 17325 20349 17359 20383
rect 18153 20349 18187 20383
rect 19809 20349 19843 20383
rect 11069 20281 11103 20315
rect 4721 20213 4755 20247
rect 27629 20213 27663 20247
rect 35173 20213 35207 20247
rect 9229 20009 9263 20043
rect 37749 20009 37783 20043
rect 1777 19873 1811 19907
rect 2789 19873 2823 19907
rect 4077 19873 4111 19907
rect 6745 19873 6779 19907
rect 7941 19873 7975 19907
rect 9873 19873 9907 19907
rect 10885 19873 10919 19907
rect 13277 19873 13311 19907
rect 19533 19873 19567 19907
rect 21281 19873 21315 19907
rect 22477 19873 22511 19907
rect 22661 19873 22695 19907
rect 24961 19873 24995 19907
rect 26801 19873 26835 19907
rect 3249 19805 3283 19839
rect 6009 19805 6043 19839
rect 9137 19805 9171 19839
rect 15485 19805 15519 19839
rect 16313 19805 16347 19839
rect 16773 19805 16807 19839
rect 18153 19805 18187 19839
rect 20177 19805 20211 19839
rect 25973 19805 26007 19839
rect 26617 19805 26651 19839
rect 36921 19805 36955 19839
rect 37013 19805 37047 19839
rect 37933 19805 37967 19839
rect 1869 19737 1903 19771
rect 4169 19737 4203 19771
rect 5089 19737 5123 19771
rect 6846 19737 6880 19771
rect 7389 19737 7423 19771
rect 8033 19737 8067 19771
rect 8585 19737 8619 19771
rect 9965 19737 9999 19771
rect 11805 19737 11839 19771
rect 11897 19737 11931 19771
rect 12449 19737 12483 19771
rect 13001 19737 13035 19771
rect 13093 19737 13127 19771
rect 14381 19737 14415 19771
rect 14473 19737 14507 19771
rect 15025 19737 15059 19771
rect 19625 19737 19659 19771
rect 21005 19737 21039 19771
rect 21097 19737 21131 19771
rect 24685 19737 24719 19771
rect 24777 19737 24811 19771
rect 3341 19669 3375 19703
rect 6101 19669 6135 19703
rect 15577 19669 15611 19703
rect 16129 19669 16163 19703
rect 16865 19669 16899 19703
rect 18245 19669 18279 19703
rect 23121 19669 23155 19703
rect 27261 19669 27295 19703
rect 4721 19465 4755 19499
rect 26065 19465 26099 19499
rect 36829 19465 36863 19499
rect 37841 19465 37875 19499
rect 1685 19397 1719 19431
rect 2881 19397 2915 19431
rect 3801 19397 3835 19431
rect 5457 19397 5491 19431
rect 6009 19397 6043 19431
rect 6653 19397 6687 19431
rect 7389 19397 7423 19431
rect 9045 19397 9079 19431
rect 11805 19397 11839 19431
rect 11897 19397 11931 19431
rect 14013 19397 14047 19431
rect 15577 19397 15611 19431
rect 17049 19397 17083 19431
rect 18337 19397 18371 19431
rect 18429 19397 18463 19431
rect 19901 19397 19935 19431
rect 4629 19329 4663 19363
rect 6561 19329 6595 19363
rect 10977 19329 11011 19363
rect 11069 19329 11103 19363
rect 13185 19329 13219 19363
rect 19809 19329 19843 19363
rect 24133 19329 24167 19363
rect 25605 19329 25639 19363
rect 26249 19329 26283 19363
rect 36737 19329 36771 19363
rect 38025 19329 38059 19363
rect 2789 19261 2823 19295
rect 5365 19261 5399 19295
rect 7297 19261 7331 19295
rect 7573 19261 7607 19295
rect 8769 19261 8803 19295
rect 12173 19261 12207 19295
rect 13277 19261 13311 19295
rect 13921 19261 13955 19295
rect 14381 19261 14415 19295
rect 15485 19261 15519 19295
rect 15761 19261 15795 19295
rect 16957 19261 16991 19295
rect 17325 19261 17359 19295
rect 19257 19261 19291 19295
rect 24777 19261 24811 19295
rect 1869 19193 1903 19227
rect 10517 19125 10551 19159
rect 24225 19125 24259 19159
rect 25421 19125 25455 19159
rect 4353 18921 4387 18955
rect 10885 18921 10919 18955
rect 21557 18921 21591 18955
rect 37473 18921 37507 18955
rect 2237 18785 2271 18819
rect 4997 18785 5031 18819
rect 5641 18785 5675 18819
rect 9413 18785 9447 18819
rect 11529 18785 11563 18819
rect 12725 18785 12759 18819
rect 13553 18785 13587 18819
rect 24685 18785 24719 18819
rect 4261 18717 4295 18751
rect 6101 18717 6135 18751
rect 8401 18717 8435 18751
rect 9137 18717 9171 18751
rect 12173 18717 12207 18751
rect 14381 18717 14415 18751
rect 16037 18717 16071 18751
rect 16957 18717 16991 18751
rect 18245 18717 18279 18751
rect 21465 18717 21499 18751
rect 26801 18717 26835 18751
rect 37657 18717 37691 18751
rect 38301 18717 38335 18751
rect 2329 18649 2363 18683
rect 2881 18649 2915 18683
rect 5089 18649 5123 18683
rect 6837 18649 6871 18683
rect 6929 18649 6963 18683
rect 7849 18649 7883 18683
rect 11621 18649 11655 18683
rect 12817 18649 12851 18683
rect 15393 18649 15427 18683
rect 15485 18649 15519 18683
rect 23397 18649 23431 18683
rect 23489 18649 23523 18683
rect 24041 18649 24075 18683
rect 24777 18649 24811 18683
rect 25329 18649 25363 18683
rect 6193 18581 6227 18615
rect 8493 18581 8527 18615
rect 14473 18581 14507 18615
rect 17049 18581 17083 18615
rect 18337 18581 18371 18615
rect 26893 18581 26927 18615
rect 38117 18581 38151 18615
rect 2053 18377 2087 18411
rect 16957 18377 16991 18411
rect 20545 18377 20579 18411
rect 38117 18377 38151 18411
rect 2789 18309 2823 18343
rect 3341 18309 3375 18343
rect 4077 18309 4111 18343
rect 6745 18309 6779 18343
rect 10618 18309 10652 18343
rect 11897 18309 11931 18343
rect 11989 18309 12023 18343
rect 13553 18309 13587 18343
rect 22201 18309 22235 18343
rect 23121 18309 23155 18343
rect 23857 18309 23891 18343
rect 24961 18309 24995 18343
rect 27813 18309 27847 18343
rect 1869 18241 1903 18275
rect 5089 18241 5123 18275
rect 15025 18241 15059 18275
rect 15209 18241 15243 18275
rect 15669 18241 15703 18275
rect 16865 18241 16899 18275
rect 17509 18241 17543 18275
rect 20453 18241 20487 18275
rect 24869 18241 24903 18275
rect 27353 18241 27387 18275
rect 31493 18241 31527 18275
rect 38301 18241 38335 18275
rect 2697 18173 2731 18207
rect 3985 18173 4019 18207
rect 4629 18173 4663 18207
rect 5917 18173 5951 18207
rect 6653 18173 6687 18207
rect 7849 18173 7883 18207
rect 8125 18173 8159 18207
rect 10517 18173 10551 18207
rect 12909 18173 12943 18207
rect 13461 18173 13495 18207
rect 14381 18173 14415 18207
rect 22109 18173 22143 18207
rect 23765 18173 23799 18207
rect 24409 18173 24443 18207
rect 27169 18173 27203 18207
rect 7205 18105 7239 18139
rect 11069 18105 11103 18139
rect 17601 18105 17635 18139
rect 9597 18037 9631 18071
rect 15761 18037 15795 18071
rect 31585 18037 31619 18071
rect 3341 17833 3375 17867
rect 5733 17833 5767 17867
rect 18061 17833 18095 17867
rect 8585 17765 8619 17799
rect 15577 17765 15611 17799
rect 16773 17765 16807 17799
rect 22109 17765 22143 17799
rect 6285 17697 6319 17731
rect 13553 17697 13587 17731
rect 19901 17697 19935 17731
rect 30757 17697 30791 17731
rect 1593 17629 1627 17663
rect 3985 17629 4019 17663
rect 6193 17629 6227 17663
rect 6837 17629 6871 17663
rect 9505 17629 9539 17663
rect 11805 17629 11839 17663
rect 14289 17629 14323 17663
rect 17325 17629 17359 17663
rect 17969 17629 18003 17663
rect 22017 17629 22051 17663
rect 22937 17629 22971 17663
rect 28089 17629 28123 17663
rect 1869 17561 1903 17595
rect 4261 17561 4295 17595
rect 7113 17561 7147 17595
rect 9781 17561 9815 17595
rect 12081 17561 12115 17595
rect 15025 17561 15059 17595
rect 15117 17561 15151 17595
rect 16221 17561 16255 17595
rect 16313 17561 16347 17595
rect 19993 17561 20027 17595
rect 20545 17561 20579 17595
rect 23121 17561 23155 17595
rect 30573 17561 30607 17595
rect 11253 17493 11287 17527
rect 14381 17493 14415 17527
rect 17417 17493 17451 17527
rect 27905 17493 27939 17527
rect 3709 17289 3743 17323
rect 6009 17289 6043 17323
rect 18429 17289 18463 17323
rect 25053 17289 25087 17323
rect 28273 17289 28307 17323
rect 4537 17221 4571 17255
rect 14565 17221 14599 17255
rect 19165 17221 19199 17255
rect 22201 17221 22235 17255
rect 6561 17153 6595 17187
rect 11989 17153 12023 17187
rect 17049 17153 17083 17187
rect 17693 17153 17727 17187
rect 18337 17153 18371 17187
rect 20177 17153 20211 17187
rect 24961 17153 24995 17187
rect 27353 17153 27387 17187
rect 28457 17153 28491 17187
rect 1961 17085 1995 17119
rect 2237 17085 2271 17119
rect 4261 17085 4295 17119
rect 6837 17085 6871 17119
rect 8861 17085 8895 17119
rect 9137 17085 9171 17119
rect 10885 17085 10919 17119
rect 12265 17085 12299 17119
rect 13737 17085 13771 17119
rect 14289 17085 14323 17119
rect 17141 17085 17175 17119
rect 17785 17085 17819 17119
rect 19073 17085 19107 17119
rect 22109 17085 22143 17119
rect 22385 17085 22419 17119
rect 27169 17085 27203 17119
rect 19625 17017 19659 17051
rect 8309 16949 8343 16983
rect 16037 16949 16071 16983
rect 20269 16949 20303 16983
rect 27629 16949 27663 16983
rect 4892 16745 4926 16779
rect 18705 16745 18739 16779
rect 1869 16609 1903 16643
rect 4629 16609 4663 16643
rect 7113 16609 7147 16643
rect 9873 16609 9907 16643
rect 10977 16609 11011 16643
rect 19533 16609 19567 16643
rect 24593 16609 24627 16643
rect 24777 16609 24811 16643
rect 1593 16541 1627 16575
rect 3985 16541 4019 16575
rect 6837 16541 6871 16575
rect 10701 16541 10735 16575
rect 13553 16541 13587 16575
rect 14289 16541 14323 16575
rect 16865 16541 16899 16575
rect 16957 16541 16991 16575
rect 17509 16541 17543 16575
rect 18889 16541 18923 16575
rect 22477 16541 22511 16575
rect 25237 16541 25271 16575
rect 38025 16541 38059 16575
rect 9137 16473 9171 16507
rect 13645 16473 13679 16507
rect 14565 16473 14599 16507
rect 17601 16473 17635 16507
rect 19618 16473 19652 16507
rect 20545 16473 20579 16507
rect 3341 16405 3375 16439
rect 4077 16405 4111 16439
rect 6377 16405 6411 16439
rect 8585 16405 8619 16439
rect 12449 16405 12483 16439
rect 16037 16405 16071 16439
rect 22569 16405 22603 16439
rect 38209 16405 38243 16439
rect 6009 16201 6043 16235
rect 6653 16201 6687 16235
rect 10425 16201 10459 16235
rect 16221 16201 16255 16235
rect 20821 16201 20855 16235
rect 27261 16201 27295 16235
rect 4537 16133 4571 16167
rect 13829 16133 13863 16167
rect 17141 16133 17175 16167
rect 17877 16133 17911 16167
rect 17969 16133 18003 16167
rect 19441 16133 19475 16167
rect 22201 16133 22235 16167
rect 23121 16133 23155 16167
rect 4261 16065 4295 16099
rect 6561 16065 6595 16099
rect 7205 16065 7239 16099
rect 9689 16065 9723 16099
rect 10333 16065 10367 16099
rect 10977 16065 11011 16099
rect 12173 16065 12207 16099
rect 16129 16065 16163 16099
rect 16865 16065 16899 16099
rect 19349 16065 19383 16099
rect 19993 16065 20027 16099
rect 20729 16065 20763 16099
rect 27169 16065 27203 16099
rect 27905 16065 27939 16099
rect 28733 16065 28767 16099
rect 38301 16065 38335 16099
rect 2053 15997 2087 16031
rect 7481 15997 7515 16031
rect 9229 15997 9263 16031
rect 12909 15997 12943 16031
rect 13553 15997 13587 16031
rect 18521 15997 18555 16031
rect 22109 15997 22143 16031
rect 27997 15997 28031 16031
rect 20085 15929 20119 15963
rect 28549 15929 28583 15963
rect 2316 15861 2350 15895
rect 3801 15861 3835 15895
rect 9781 15861 9815 15895
rect 11069 15861 11103 15895
rect 15301 15861 15335 15895
rect 38117 15861 38151 15895
rect 9137 15657 9171 15691
rect 13001 15657 13035 15691
rect 21097 15657 21131 15691
rect 29837 15589 29871 15623
rect 1869 15521 1903 15555
rect 3341 15521 3375 15555
rect 4169 15521 4203 15555
rect 4445 15521 4479 15555
rect 5917 15521 5951 15555
rect 7021 15521 7055 15555
rect 10885 15521 10919 15555
rect 12357 15521 12391 15555
rect 15209 15521 15243 15555
rect 16129 15521 16163 15555
rect 20177 15521 20211 15555
rect 21741 15521 21775 15555
rect 22753 15521 22787 15555
rect 1593 15453 1627 15487
rect 6745 15453 6779 15487
rect 9321 15453 9355 15487
rect 9781 15453 9815 15487
rect 10609 15453 10643 15487
rect 12909 15453 12943 15487
rect 13553 15453 13587 15487
rect 14473 15453 14507 15487
rect 16773 15453 16807 15487
rect 19441 15453 19475 15487
rect 20085 15453 20119 15487
rect 21005 15453 21039 15487
rect 27813 15453 27847 15487
rect 29745 15453 29779 15487
rect 13645 15385 13679 15419
rect 15301 15385 15335 15419
rect 17049 15385 17083 15419
rect 18245 15385 18279 15419
rect 18337 15385 18371 15419
rect 18889 15385 18923 15419
rect 21833 15385 21867 15419
rect 8493 15317 8527 15351
rect 9873 15317 9907 15351
rect 14565 15317 14599 15351
rect 19533 15317 19567 15351
rect 27629 15317 27663 15351
rect 3341 15113 3375 15147
rect 5549 15113 5583 15147
rect 8585 15113 8619 15147
rect 15577 15113 15611 15147
rect 19349 15113 19383 15147
rect 4077 15045 4111 15079
rect 16221 15045 16255 15079
rect 17049 15045 17083 15079
rect 12173 14977 12207 15011
rect 14841 14977 14875 15011
rect 15485 14977 15519 15011
rect 16129 14977 16163 15011
rect 18429 14977 18463 15011
rect 19533 14977 19567 15011
rect 20177 14977 20211 15011
rect 20637 14977 20671 15011
rect 22201 14977 22235 15011
rect 27997 14977 28031 15011
rect 1593 14909 1627 14943
rect 1869 14909 1903 14943
rect 3801 14909 3835 14943
rect 6837 14909 6871 14943
rect 7113 14909 7147 14943
rect 9045 14909 9079 14943
rect 12449 14909 12483 14943
rect 16957 14909 16991 14943
rect 17877 14909 17911 14943
rect 18613 14909 18647 14943
rect 25697 14909 25731 14943
rect 10793 14841 10827 14875
rect 13921 14841 13955 14875
rect 20729 14841 20763 14875
rect 9302 14773 9336 14807
rect 14933 14773 14967 14807
rect 19993 14773 20027 14807
rect 22017 14773 22051 14807
rect 27813 14773 27847 14807
rect 3341 14569 3375 14603
rect 5549 14569 5583 14603
rect 6193 14569 6227 14603
rect 9400 14569 9434 14603
rect 14552 14569 14586 14603
rect 16037 14569 16071 14603
rect 21925 14569 21959 14603
rect 25513 14569 25547 14603
rect 26341 14569 26375 14603
rect 11437 14501 11471 14535
rect 19441 14501 19475 14535
rect 1593 14433 1627 14467
rect 4721 14433 4755 14467
rect 6745 14433 6779 14467
rect 7021 14433 7055 14467
rect 9137 14433 9171 14467
rect 10885 14433 10919 14467
rect 16773 14433 16807 14467
rect 25973 14433 26007 14467
rect 26157 14433 26191 14467
rect 3985 14365 4019 14399
rect 6101 14365 6135 14399
rect 11345 14365 11379 14399
rect 11989 14365 12023 14399
rect 13553 14365 13587 14399
rect 14289 14365 14323 14399
rect 16589 14365 16623 14399
rect 19625 14365 19659 14399
rect 21281 14365 21315 14399
rect 22109 14365 22143 14399
rect 24869 14365 24903 14399
rect 25053 14365 25087 14399
rect 27077 14365 27111 14399
rect 38025 14365 38059 14399
rect 1869 14297 1903 14331
rect 5457 14297 5491 14331
rect 17785 14297 17819 14331
rect 17877 14297 17911 14331
rect 18429 14297 18463 14331
rect 27169 14297 27203 14331
rect 8493 14229 8527 14263
rect 12081 14229 12115 14263
rect 13645 14229 13679 14263
rect 17233 14229 17267 14263
rect 20637 14229 20671 14263
rect 21373 14229 21407 14263
rect 38209 14229 38243 14263
rect 1777 14025 1811 14059
rect 4629 14025 4663 14059
rect 5825 14025 5859 14059
rect 6745 14025 6779 14059
rect 7389 14025 7423 14059
rect 8033 14025 8067 14059
rect 10333 14025 10367 14059
rect 10977 14025 11011 14059
rect 2237 13957 2271 13991
rect 8861 13957 8895 13991
rect 14749 13957 14783 13991
rect 17049 13957 17083 13991
rect 17693 13957 17727 13991
rect 17785 13957 17819 13991
rect 19809 13957 19843 13991
rect 20453 13957 20487 13991
rect 20545 13957 20579 13991
rect 21465 13957 21499 13991
rect 1593 13889 1627 13923
rect 2881 13889 2915 13923
rect 5089 13889 5123 13923
rect 5733 13889 5767 13923
rect 6653 13889 6687 13923
rect 7297 13889 7331 13923
rect 7941 13889 7975 13923
rect 10885 13889 10919 13923
rect 11989 13889 12023 13923
rect 16129 13889 16163 13923
rect 16957 13889 16991 13923
rect 18797 13889 18831 13923
rect 19073 13889 19107 13923
rect 19717 13889 19751 13923
rect 22017 13889 22051 13923
rect 5181 13821 5215 13855
rect 8585 13821 8619 13855
rect 13737 13821 13771 13855
rect 14657 13821 14691 13855
rect 15669 13821 15703 13855
rect 17969 13821 18003 13855
rect 16221 13753 16255 13787
rect 3144 13685 3178 13719
rect 12252 13685 12286 13719
rect 22109 13685 22143 13719
rect 3341 13481 3375 13515
rect 8125 13481 8159 13515
rect 9768 13481 9802 13515
rect 20729 13481 20763 13515
rect 22201 13481 22235 13515
rect 5825 13413 5859 13447
rect 11253 13413 11287 13447
rect 26433 13413 26467 13447
rect 1869 13345 1903 13379
rect 9505 13345 9539 13379
rect 11713 13345 11747 13379
rect 16589 13345 16623 13379
rect 26065 13345 26099 13379
rect 1593 13277 1627 13311
rect 4077 13277 4111 13311
rect 6377 13277 6411 13311
rect 17233 13277 17267 13311
rect 18613 13277 18647 13311
rect 18705 13277 18739 13311
rect 20637 13277 20671 13311
rect 22109 13277 22143 13311
rect 26249 13277 26283 13311
rect 34345 13277 34379 13311
rect 38025 13277 38059 13311
rect 4353 13209 4387 13243
rect 6653 13209 6687 13243
rect 11989 13209 12023 13243
rect 13737 13209 13771 13243
rect 14381 13209 14415 13243
rect 14473 13209 14507 13243
rect 15393 13209 15427 13243
rect 15853 13209 15887 13243
rect 18061 13209 18095 13243
rect 19533 13209 19567 13243
rect 19625 13209 19659 13243
rect 20177 13209 20211 13243
rect 34161 13141 34195 13175
rect 38209 13141 38243 13175
rect 9229 12937 9263 12971
rect 20913 12937 20947 12971
rect 27537 12937 27571 12971
rect 10609 12869 10643 12903
rect 15669 12869 15703 12903
rect 15761 12869 15795 12903
rect 17325 12869 17359 12903
rect 18153 12869 18187 12903
rect 18245 12869 18279 12903
rect 19809 12869 19843 12903
rect 22385 12869 22419 12903
rect 3893 12801 3927 12835
rect 6561 12801 6595 12835
rect 7481 12801 7515 12835
rect 9873 12801 9907 12835
rect 11713 12801 11747 12835
rect 12633 12801 12667 12835
rect 13277 12801 13311 12835
rect 16957 12801 16991 12835
rect 20821 12801 20855 12835
rect 22201 12801 22235 12835
rect 27721 12801 27755 12835
rect 28365 12801 28399 12835
rect 38117 12801 38151 12835
rect 1593 12733 1627 12767
rect 1869 12733 1903 12767
rect 4169 12733 4203 12767
rect 7757 12733 7791 12767
rect 13553 12733 13587 12767
rect 16313 12733 16347 12767
rect 18429 12733 18463 12767
rect 19717 12733 19751 12767
rect 20361 12733 20395 12767
rect 3341 12665 3375 12699
rect 5641 12665 5675 12699
rect 28181 12665 28215 12699
rect 6745 12597 6779 12631
rect 11805 12597 11839 12631
rect 12725 12597 12759 12631
rect 15025 12597 15059 12631
rect 38209 12597 38243 12631
rect 7297 12393 7331 12427
rect 9229 12393 9263 12427
rect 11529 12393 11563 12427
rect 12252 12393 12286 12427
rect 13737 12393 13771 12427
rect 16037 12393 16071 12427
rect 3341 12325 3375 12359
rect 7941 12325 7975 12359
rect 1869 12257 1903 12291
rect 4721 12257 4755 12291
rect 5549 12257 5583 12291
rect 11989 12257 12023 12291
rect 14289 12257 14323 12291
rect 16589 12257 16623 12291
rect 17785 12257 17819 12291
rect 19533 12257 19567 12291
rect 20913 12257 20947 12291
rect 24869 12257 24903 12291
rect 25053 12257 25087 12291
rect 26985 12257 27019 12291
rect 1593 12189 1627 12223
rect 7849 12189 7883 12223
rect 9137 12189 9171 12223
rect 9781 12189 9815 12223
rect 19441 12189 19475 12223
rect 22109 12189 22143 12223
rect 26893 12189 26927 12223
rect 3985 12121 4019 12155
rect 5825 12121 5859 12155
rect 10057 12121 10091 12155
rect 14565 12121 14599 12155
rect 16681 12121 16715 12155
rect 17233 12121 17267 12155
rect 17877 12121 17911 12155
rect 18429 12121 18463 12155
rect 20637 12121 20671 12155
rect 20729 12121 20763 12155
rect 22201 12053 22235 12087
rect 25513 12053 25547 12087
rect 6653 11849 6687 11883
rect 20545 11849 20579 11883
rect 7481 11781 7515 11815
rect 15025 11781 15059 11815
rect 15761 11781 15795 11815
rect 16313 11781 16347 11815
rect 17049 11781 17083 11815
rect 17601 11781 17635 11815
rect 21189 11781 21223 11815
rect 22201 11781 22235 11815
rect 2053 11713 2087 11747
rect 4261 11713 4295 11747
rect 6561 11713 6595 11747
rect 9413 11713 9447 11747
rect 11713 11713 11747 11747
rect 12357 11713 12391 11747
rect 12449 11713 12483 11747
rect 13001 11713 13035 11747
rect 18061 11713 18095 11747
rect 18981 11713 19015 11747
rect 20453 11713 20487 11747
rect 21097 11713 21131 11747
rect 23581 11713 23615 11747
rect 2329 11645 2363 11679
rect 4537 11645 4571 11679
rect 7205 11645 7239 11679
rect 9689 11645 9723 11679
rect 13277 11645 13311 11679
rect 15669 11645 15703 11679
rect 16957 11645 16991 11679
rect 18245 11645 18279 11679
rect 19165 11645 19199 11679
rect 22109 11645 22143 11679
rect 22385 11645 22419 11679
rect 11161 11577 11195 11611
rect 3801 11509 3835 11543
rect 6009 11509 6043 11543
rect 8953 11509 8987 11543
rect 11805 11509 11839 11543
rect 23673 11509 23707 11543
rect 3341 11305 3375 11339
rect 4616 11305 4650 11339
rect 6824 11305 6858 11339
rect 9229 11305 9263 11339
rect 16037 11305 16071 11339
rect 23305 11305 23339 11339
rect 11529 11237 11563 11271
rect 13737 11237 13771 11271
rect 20085 11237 20119 11271
rect 1593 11169 1627 11203
rect 1869 11169 1903 11203
rect 4353 11169 4387 11203
rect 6561 11169 6595 11203
rect 11989 11169 12023 11203
rect 16681 11169 16715 11203
rect 17693 11169 17727 11203
rect 37749 11169 37783 11203
rect 9137 11101 9171 11135
rect 9781 11101 9815 11135
rect 14289 11101 14323 11135
rect 18153 11101 18187 11135
rect 20637 11101 20671 11135
rect 21281 11101 21315 11135
rect 21925 11101 21959 11135
rect 22569 11101 22603 11135
rect 23213 11101 23247 11135
rect 26065 11101 26099 11135
rect 37473 11101 37507 11135
rect 8585 11033 8619 11067
rect 10057 11033 10091 11067
rect 12265 11033 12299 11067
rect 14565 11033 14599 11067
rect 16773 11033 16807 11067
rect 18429 11033 18463 11067
rect 19533 11033 19567 11067
rect 19625 11033 19659 11067
rect 22017 11033 22051 11067
rect 26157 11033 26191 11067
rect 6101 10965 6135 10999
rect 20729 10965 20763 10999
rect 21373 10965 21407 10999
rect 22661 10965 22695 10999
rect 1961 10761 1995 10795
rect 2605 10761 2639 10795
rect 3249 10761 3283 10795
rect 5549 10761 5583 10795
rect 11805 10761 11839 10795
rect 12449 10761 12483 10795
rect 17509 10761 17543 10795
rect 10701 10693 10735 10727
rect 13277 10693 13311 10727
rect 15761 10693 15795 10727
rect 18153 10693 18187 10727
rect 19717 10693 19751 10727
rect 20913 10693 20947 10727
rect 1869 10625 1903 10659
rect 2513 10625 2547 10659
rect 3157 10625 3191 10659
rect 3801 10625 3835 10659
rect 6745 10625 6779 10659
rect 8953 10625 8987 10659
rect 11705 10623 11739 10657
rect 12357 10625 12391 10659
rect 17049 10625 17083 10659
rect 22017 10625 22051 10659
rect 22661 10625 22695 10659
rect 23489 10625 23523 10659
rect 24685 10625 24719 10659
rect 4077 10557 4111 10591
rect 7021 10557 7055 10591
rect 13001 10557 13035 10591
rect 15025 10557 15059 10591
rect 15669 10557 15703 10591
rect 16865 10557 16899 10591
rect 18061 10557 18095 10591
rect 19073 10557 19107 10591
rect 19625 10557 19659 10591
rect 20821 10557 20855 10591
rect 23581 10557 23615 10591
rect 16221 10489 16255 10523
rect 20177 10489 20211 10523
rect 21373 10489 21407 10523
rect 22753 10489 22787 10523
rect 8493 10421 8527 10455
rect 22109 10421 22143 10455
rect 24501 10421 24535 10455
rect 2605 10217 2639 10251
rect 3341 10217 3375 10251
rect 5733 10217 5767 10251
rect 9689 10217 9723 10251
rect 10333 10217 10367 10251
rect 2053 10149 2087 10183
rect 21649 10149 21683 10183
rect 29837 10149 29871 10183
rect 4261 10081 4295 10115
rect 10885 10081 10919 10115
rect 14289 10081 14323 10115
rect 17325 10081 17359 10115
rect 19533 10081 19567 10115
rect 20545 10081 20579 10115
rect 22477 10081 22511 10115
rect 23489 10081 23523 10115
rect 1961 10013 1995 10047
rect 2789 10013 2823 10047
rect 3249 10013 3283 10047
rect 3985 10013 4019 10047
rect 6469 10013 6503 10047
rect 9597 10013 9631 10047
rect 10241 10013 10275 10047
rect 12909 10013 12943 10047
rect 13553 10013 13587 10047
rect 16589 10013 16623 10047
rect 17969 10013 18003 10047
rect 22293 10013 22327 10047
rect 23397 10013 23431 10047
rect 29745 10013 29779 10047
rect 38025 10013 38059 10047
rect 6745 9945 6779 9979
rect 11161 9945 11195 9979
rect 14565 9945 14599 9979
rect 18245 9945 18279 9979
rect 19625 9945 19659 9979
rect 21097 9945 21131 9979
rect 21189 9945 21223 9979
rect 22937 9945 22971 9979
rect 8217 9877 8251 9911
rect 13645 9877 13679 9911
rect 16037 9877 16071 9911
rect 25053 9877 25087 9911
rect 38209 9877 38243 9911
rect 6009 9673 6043 9707
rect 18337 9673 18371 9707
rect 22661 9673 22695 9707
rect 7665 9605 7699 9639
rect 8493 9605 8527 9639
rect 11713 9605 11747 9639
rect 12449 9605 12483 9639
rect 13277 9605 13311 9639
rect 19257 9605 19291 9639
rect 19901 9605 19935 9639
rect 20913 9605 20947 9639
rect 23489 9605 23523 9639
rect 24961 9605 24995 9639
rect 25053 9605 25087 9639
rect 6929 9537 6963 9571
rect 8393 9537 8427 9571
rect 13185 9537 13219 9571
rect 13829 9537 13863 9571
rect 16313 9537 16347 9571
rect 16865 9537 16899 9571
rect 17693 9537 17727 9571
rect 17877 9537 17911 9571
rect 19165 9537 19199 9571
rect 19809 9537 19843 9571
rect 21465 9537 21499 9571
rect 22017 9537 22051 9571
rect 22109 9537 22143 9571
rect 23397 9537 23431 9571
rect 24041 9537 24075 9571
rect 29929 9537 29963 9571
rect 1593 9469 1627 9503
rect 1869 9469 1903 9503
rect 4261 9469 4295 9503
rect 4537 9469 4571 9503
rect 9045 9469 9079 9503
rect 9321 9469 9355 9503
rect 14105 9469 14139 9503
rect 20821 9469 20855 9503
rect 25237 9469 25271 9503
rect 10793 9401 10827 9435
rect 3341 9333 3375 9367
rect 15577 9333 15611 9367
rect 16129 9333 16163 9367
rect 17049 9333 17083 9367
rect 24133 9333 24167 9367
rect 30021 9333 30055 9367
rect 2053 9129 2087 9163
rect 2605 9129 2639 9163
rect 3341 9129 3375 9163
rect 6653 9129 6687 9163
rect 12633 9129 12667 9163
rect 13277 9129 13311 9163
rect 23489 9129 23523 9163
rect 5457 9061 5491 9095
rect 11713 9061 11747 9095
rect 4721 8993 4755 9027
rect 9965 8993 9999 9027
rect 14289 8993 14323 9027
rect 16037 8993 16071 9027
rect 16589 8993 16623 9027
rect 1961 8925 1995 8959
rect 2789 8925 2823 8959
rect 3249 8925 3283 8959
rect 3985 8925 4019 8959
rect 5365 8925 5399 8959
rect 6561 8925 6595 8959
rect 8401 8925 8435 8959
rect 9321 8925 9355 8959
rect 12541 8925 12575 8959
rect 13185 8925 13219 8959
rect 19717 8925 19751 8959
rect 21649 8925 21683 8959
rect 22109 8925 22143 8959
rect 22753 8925 22787 8959
rect 23397 8925 23431 8959
rect 24593 8925 24627 8959
rect 7665 8857 7699 8891
rect 10241 8857 10275 8891
rect 14565 8857 14599 8891
rect 16681 8857 16715 8891
rect 17601 8857 17635 8891
rect 18153 8857 18187 8891
rect 18245 8857 18279 8891
rect 18797 8857 18831 8891
rect 21005 8857 21039 8891
rect 21097 8857 21131 8891
rect 9413 8789 9447 8823
rect 19809 8789 19843 8823
rect 22201 8789 22235 8823
rect 22845 8789 22879 8823
rect 24685 8789 24719 8823
rect 1593 8585 1627 8619
rect 5089 8585 5123 8619
rect 7205 8585 7239 8619
rect 9689 8517 9723 8551
rect 17049 8517 17083 8551
rect 17601 8517 17635 8551
rect 18337 8517 18371 8551
rect 19441 8517 19475 8551
rect 38301 8517 38335 8551
rect 1777 8449 1811 8483
rect 4445 8449 4479 8483
rect 4537 8449 4571 8483
rect 5273 8449 5307 8483
rect 6561 8449 6595 8483
rect 7389 8449 7423 8483
rect 8769 8449 8803 8483
rect 11713 8449 11747 8483
rect 13921 8449 13955 8483
rect 16129 8449 16163 8483
rect 18061 8449 18095 8483
rect 22661 8449 22695 8483
rect 23305 8449 23339 8483
rect 23949 8449 23983 8483
rect 24593 8449 24627 8483
rect 25237 8449 25271 8483
rect 38117 8449 38151 8483
rect 2237 8381 2271 8415
rect 2513 8381 2547 8415
rect 6653 8381 6687 8415
rect 9413 8381 9447 8415
rect 11161 8381 11195 8415
rect 11989 8381 12023 8415
rect 14197 8381 14231 8415
rect 16221 8381 16255 8415
rect 16957 8381 16991 8415
rect 19349 8381 19383 8415
rect 20361 8381 20395 8415
rect 21005 8381 21039 8415
rect 22017 8381 22051 8415
rect 22753 8381 22787 8415
rect 8861 8313 8895 8347
rect 13461 8313 13495 8347
rect 24041 8313 24075 8347
rect 25329 8313 25363 8347
rect 3985 8245 4019 8279
rect 15669 8245 15703 8279
rect 23397 8245 23431 8279
rect 24685 8245 24719 8279
rect 3433 8041 3467 8075
rect 6009 8041 6043 8075
rect 6837 8041 6871 8075
rect 11345 8041 11379 8075
rect 16037 8041 16071 8075
rect 11713 7973 11747 8007
rect 1685 7905 1719 7939
rect 1961 7905 1995 7939
rect 9873 7905 9907 7939
rect 11989 7905 12023 7939
rect 12265 7905 12299 7939
rect 14565 7905 14599 7939
rect 16589 7905 16623 7939
rect 17601 7905 17635 7939
rect 19533 7905 19567 7939
rect 20177 7905 20211 7939
rect 29837 7905 29871 7939
rect 37749 7905 37783 7939
rect 4077 7837 4111 7871
rect 5917 7837 5951 7871
rect 6745 7837 6779 7871
rect 9597 7837 9631 7871
rect 14289 7837 14323 7871
rect 19441 7837 19475 7871
rect 23213 7837 23247 7871
rect 23857 7837 23891 7871
rect 24777 7837 24811 7871
rect 29745 7837 29779 7871
rect 37473 7837 37507 7871
rect 16681 7769 16715 7803
rect 18245 7769 18279 7803
rect 18346 7769 18380 7803
rect 18889 7769 18923 7803
rect 20269 7769 20303 7803
rect 21189 7769 21223 7803
rect 21741 7769 21775 7803
rect 21833 7769 21867 7803
rect 22753 7769 22787 7803
rect 4169 7701 4203 7735
rect 13737 7701 13771 7735
rect 23305 7701 23339 7735
rect 23949 7701 23983 7735
rect 24593 7701 24627 7735
rect 4537 7497 4571 7531
rect 8401 7497 8435 7531
rect 25513 7497 25547 7531
rect 27261 7497 27295 7531
rect 1685 7429 1719 7463
rect 5917 7429 5951 7463
rect 9137 7429 9171 7463
rect 17417 7429 17451 7463
rect 18337 7429 18371 7463
rect 18889 7429 18923 7463
rect 18981 7429 19015 7463
rect 2789 7361 2823 7395
rect 5825 7361 5859 7395
rect 11713 7361 11747 7395
rect 20821 7361 20855 7395
rect 22017 7361 22051 7395
rect 22201 7361 22235 7395
rect 23121 7361 23155 7395
rect 23949 7361 23983 7395
rect 25421 7361 25455 7395
rect 27169 7361 27203 7395
rect 3065 7293 3099 7327
rect 6653 7293 6687 7327
rect 8861 7293 8895 7327
rect 11989 7293 12023 7327
rect 13461 7293 13495 7327
rect 14013 7293 14047 7327
rect 14289 7293 14323 7327
rect 15761 7293 15795 7327
rect 17325 7293 17359 7327
rect 19901 7293 19935 7327
rect 21005 7293 21039 7327
rect 23213 7293 23247 7327
rect 1869 7225 1903 7259
rect 21465 7225 21499 7259
rect 22385 7225 22419 7259
rect 23765 7225 23799 7259
rect 6916 7157 6950 7191
rect 10609 7157 10643 7191
rect 5536 6953 5570 6987
rect 9965 6953 9999 6987
rect 12909 6953 12943 6987
rect 14552 6953 14586 6987
rect 22661 6953 22695 6987
rect 1777 6885 1811 6919
rect 16037 6885 16071 6919
rect 17141 6885 17175 6919
rect 20085 6885 20119 6919
rect 4077 6817 4111 6851
rect 5273 6817 5307 6851
rect 7021 6817 7055 6851
rect 11161 6817 11195 6851
rect 13461 6817 13495 6851
rect 17785 6817 17819 6851
rect 18061 6817 18095 6851
rect 20637 6817 20671 6851
rect 21373 6817 21407 6851
rect 22017 6817 22051 6851
rect 1593 6749 1627 6783
rect 2513 6749 2547 6783
rect 3157 6749 3191 6783
rect 3985 6749 4019 6783
rect 7849 6749 7883 6783
rect 9229 6749 9263 6783
rect 9321 6749 9355 6783
rect 9865 6743 9899 6777
rect 10517 6749 10551 6783
rect 13369 6749 13403 6783
rect 14289 6749 14323 6783
rect 21281 6749 21315 6783
rect 21925 6749 21959 6783
rect 22569 6749 22603 6783
rect 23213 6749 23247 6783
rect 23305 6749 23339 6783
rect 23857 6749 23891 6783
rect 11437 6681 11471 6715
rect 16589 6681 16623 6715
rect 16681 6681 16715 6715
rect 17877 6681 17911 6715
rect 19533 6681 19567 6715
rect 19625 6681 19659 6715
rect 23949 6681 23983 6715
rect 2329 6613 2363 6647
rect 2973 6613 3007 6647
rect 7665 6613 7699 6647
rect 10609 6613 10643 6647
rect 1961 6409 1995 6443
rect 4537 6409 4571 6443
rect 8309 6409 8343 6443
rect 20361 6409 20395 6443
rect 38117 6409 38151 6443
rect 5089 6341 5123 6375
rect 11713 6341 11747 6375
rect 17785 6341 17819 6375
rect 21005 6341 21039 6375
rect 22661 6341 22695 6375
rect 1869 6273 1903 6307
rect 2697 6273 2731 6307
rect 3525 6273 3559 6307
rect 4445 6273 4479 6307
rect 6561 6273 6595 6307
rect 9045 6273 9079 6307
rect 12449 6273 12483 6307
rect 15853 6273 15887 6307
rect 16865 6273 16899 6307
rect 19165 6273 19199 6307
rect 20269 6273 20303 6307
rect 20913 6273 20947 6307
rect 30573 6273 30607 6307
rect 38301 6273 38335 6307
rect 5825 6205 5859 6239
rect 6837 6205 6871 6239
rect 9321 6205 9355 6239
rect 13461 6205 13495 6239
rect 13737 6205 13771 6239
rect 15669 6205 15703 6239
rect 17693 6205 17727 6239
rect 18153 6205 18187 6239
rect 19349 6205 19383 6239
rect 22569 6205 22603 6239
rect 23213 6205 23247 6239
rect 30665 6137 30699 6171
rect 2513 6069 2547 6103
rect 3341 6069 3375 6103
rect 8677 6069 8711 6103
rect 10793 6069 10827 6103
rect 15209 6069 15243 6103
rect 16313 6069 16347 6103
rect 16957 6069 16991 6103
rect 19533 6069 19567 6103
rect 3341 5865 3375 5899
rect 11069 5865 11103 5899
rect 11792 5865 11826 5899
rect 18429 5865 18463 5899
rect 20453 5865 20487 5899
rect 3985 5797 4019 5831
rect 7849 5797 7883 5831
rect 23673 5797 23707 5831
rect 1869 5729 1903 5763
rect 5273 5729 5307 5763
rect 9321 5729 9355 5763
rect 9597 5729 9631 5763
rect 11529 5729 11563 5763
rect 16589 5729 16623 5763
rect 17601 5729 17635 5763
rect 21741 5729 21775 5763
rect 22293 5729 22327 5763
rect 1593 5661 1627 5695
rect 4169 5661 4203 5695
rect 4813 5661 4847 5695
rect 7757 5661 7791 5695
rect 8401 5661 8435 5695
rect 14289 5661 14323 5695
rect 18061 5661 18095 5695
rect 18245 5661 18279 5695
rect 19441 5661 19475 5695
rect 20361 5661 20395 5695
rect 21005 5661 21039 5695
rect 21649 5661 21683 5695
rect 22937 5661 22971 5695
rect 23581 5661 23615 5695
rect 25697 5661 25731 5695
rect 5549 5593 5583 5627
rect 7297 5593 7331 5627
rect 14565 5593 14599 5627
rect 16681 5593 16715 5627
rect 19717 5593 19751 5627
rect 23029 5593 23063 5627
rect 4629 5525 4663 5559
rect 8493 5525 8527 5559
rect 13277 5525 13311 5559
rect 16037 5525 16071 5559
rect 21097 5525 21131 5559
rect 25789 5525 25823 5559
rect 3433 5321 3467 5355
rect 23857 5321 23891 5355
rect 6929 5253 6963 5287
rect 7757 5253 7791 5287
rect 12081 5253 12115 5287
rect 12909 5253 12943 5287
rect 16957 5253 16991 5287
rect 17049 5253 17083 5287
rect 18521 5253 18555 5287
rect 18613 5253 18647 5287
rect 20085 5253 20119 5287
rect 22109 5253 22143 5287
rect 22201 5253 22235 5287
rect 1593 5185 1627 5219
rect 3341 5185 3375 5219
rect 8309 5185 8343 5219
rect 10977 5185 11011 5219
rect 13461 5185 13495 5219
rect 15853 5185 15887 5219
rect 21097 5185 21131 5219
rect 22753 5185 22787 5219
rect 23213 5185 23247 5219
rect 24041 5185 24075 5219
rect 26433 5185 26467 5219
rect 29561 5185 29595 5219
rect 30389 5185 30423 5219
rect 38025 5185 38059 5219
rect 1869 5117 1903 5151
rect 3985 5117 4019 5151
rect 4261 5117 4295 5151
rect 8585 5117 8619 5151
rect 10057 5117 10091 5151
rect 13737 5117 13771 5151
rect 15669 5117 15703 5151
rect 17877 5117 17911 5151
rect 18797 5117 18831 5151
rect 19993 5117 20027 5151
rect 20637 5117 20671 5151
rect 15209 5049 15243 5083
rect 5733 4981 5767 5015
rect 11069 4981 11103 5015
rect 16313 4981 16347 5015
rect 21189 4981 21223 5015
rect 23305 4981 23339 5015
rect 26249 4981 26283 5015
rect 29653 4981 29687 5015
rect 30205 4981 30239 5015
rect 38209 4981 38243 5015
rect 1948 4777 1982 4811
rect 4077 4777 4111 4811
rect 9952 4777 9986 4811
rect 23213 4777 23247 4811
rect 23857 4777 23891 4811
rect 13737 4709 13771 4743
rect 16037 4709 16071 4743
rect 17141 4709 17175 4743
rect 24685 4709 24719 4743
rect 1685 4641 1719 4675
rect 6101 4641 6135 4675
rect 6377 4641 6411 4675
rect 9689 4641 9723 4675
rect 11989 4641 12023 4675
rect 16589 4641 16623 4675
rect 18245 4641 18279 4675
rect 18521 4641 18555 4675
rect 19625 4641 19659 4675
rect 21281 4641 21315 4675
rect 3985 4573 4019 4607
rect 4813 4573 4847 4607
rect 5457 4573 5491 4607
rect 14289 4573 14323 4607
rect 19441 4573 19475 4607
rect 20545 4573 20579 4607
rect 21189 4573 21223 4607
rect 21833 4573 21867 4607
rect 23121 4573 23155 4607
rect 23765 4573 23799 4607
rect 24593 4573 24627 4607
rect 25237 4573 25271 4607
rect 38025 4573 38059 4607
rect 4905 4505 4939 4539
rect 8125 4505 8159 4539
rect 12265 4505 12299 4539
rect 14565 4505 14599 4539
rect 16681 4505 16715 4539
rect 18337 4505 18371 4539
rect 20085 4505 20119 4539
rect 22477 4505 22511 4539
rect 25329 4505 25363 4539
rect 3433 4437 3467 4471
rect 5549 4437 5583 4471
rect 11437 4437 11471 4471
rect 20637 4437 20671 4471
rect 21925 4437 21959 4471
rect 37841 4437 37875 4471
rect 18613 4233 18647 4267
rect 20637 4233 20671 4267
rect 1685 4165 1719 4199
rect 3624 4165 3658 4199
rect 13553 4165 13587 4199
rect 1869 4097 1903 4131
rect 2881 4097 2915 4131
rect 3341 4097 3375 4131
rect 6009 4097 6043 4131
rect 6561 4097 6595 4131
rect 7205 4097 7239 4131
rect 9413 4097 9447 4131
rect 11989 4097 12023 4131
rect 12633 4097 12667 4131
rect 13277 4097 13311 4131
rect 16129 4097 16163 4131
rect 16221 4097 16255 4131
rect 19257 4097 19291 4131
rect 19901 4097 19935 4131
rect 19993 4097 20027 4131
rect 20545 4097 20579 4131
rect 21189 4097 21223 4131
rect 22017 4097 22051 4131
rect 22661 4097 22695 4131
rect 23305 4097 23339 4131
rect 23949 4097 23983 4131
rect 24593 4097 24627 4131
rect 24685 4097 24719 4131
rect 25237 4097 25271 4131
rect 26065 4097 26099 4131
rect 38301 4097 38335 4131
rect 7481 4029 7515 4063
rect 9689 4029 9723 4063
rect 12725 4029 12759 4063
rect 15301 4029 15335 4063
rect 16865 4029 16899 4063
rect 17141 4029 17175 4063
rect 21281 4029 21315 4063
rect 24041 4029 24075 4063
rect 5089 3961 5123 3995
rect 6653 3961 6687 3995
rect 12081 3961 12115 3995
rect 22753 3961 22787 3995
rect 38117 3961 38151 3995
rect 2697 3893 2731 3927
rect 5825 3893 5859 3927
rect 8953 3893 8987 3927
rect 11161 3893 11195 3927
rect 19349 3893 19383 3927
rect 22109 3893 22143 3927
rect 23397 3893 23431 3927
rect 25329 3893 25363 3927
rect 25881 3893 25915 3927
rect 1961 3689 1995 3723
rect 16037 3689 16071 3723
rect 18153 3689 18187 3723
rect 18797 3689 18831 3723
rect 20269 3689 20303 3723
rect 22845 3689 22879 3723
rect 24685 3689 24719 3723
rect 25329 3689 25363 3723
rect 37473 3689 37507 3723
rect 38117 3689 38151 3723
rect 6193 3553 6227 3587
rect 6837 3553 6871 3587
rect 8585 3553 8619 3587
rect 10057 3553 10091 3587
rect 11253 3553 11287 3587
rect 14289 3553 14323 3587
rect 26617 3553 26651 3587
rect 2145 3485 2179 3519
rect 2789 3485 2823 3519
rect 3433 3485 3467 3519
rect 4261 3485 4295 3519
rect 4905 3485 4939 3519
rect 9321 3485 9355 3519
rect 9965 3485 9999 3519
rect 10609 3485 10643 3519
rect 13277 3485 13311 3519
rect 18061 3485 18095 3519
rect 18705 3485 18739 3519
rect 19441 3485 19475 3519
rect 20177 3485 20211 3519
rect 20821 3485 20855 3519
rect 21465 3485 21499 3519
rect 22109 3485 22143 3519
rect 22753 3485 22787 3519
rect 23397 3485 23431 3519
rect 24593 3485 24627 3519
rect 25237 3485 25271 3519
rect 25881 3485 25915 3519
rect 26525 3485 26559 3519
rect 37657 3485 37691 3519
rect 38301 3485 38335 3519
rect 4353 3417 4387 3451
rect 7113 3417 7147 3451
rect 11529 3417 11563 3451
rect 14565 3417 14599 3451
rect 16589 3417 16623 3451
rect 16681 3417 16715 3451
rect 17601 3417 17635 3451
rect 19717 3417 19751 3451
rect 25973 3417 26007 3451
rect 2605 3349 2639 3383
rect 3249 3349 3283 3383
rect 4997 3349 5031 3383
rect 5549 3349 5583 3383
rect 9413 3349 9447 3383
rect 10701 3349 10735 3383
rect 20913 3349 20947 3383
rect 21557 3349 21591 3383
rect 22201 3349 22235 3383
rect 23489 3349 23523 3383
rect 3433 3145 3467 3179
rect 5457 3145 5491 3179
rect 22661 3145 22695 3179
rect 37473 3145 37507 3179
rect 12265 3077 12299 3111
rect 13461 3077 13495 3111
rect 15669 3077 15703 3111
rect 15761 3077 15795 3111
rect 17049 3077 17083 3111
rect 18153 3077 18187 3111
rect 18889 3077 18923 3111
rect 20361 3077 20395 3111
rect 20453 3077 20487 3111
rect 21005 3077 21039 3111
rect 27261 3077 27295 3111
rect 1593 3009 1627 3043
rect 2881 3009 2915 3043
rect 3341 3009 3375 3043
rect 3985 3009 4019 3043
rect 4629 3009 4663 3043
rect 5457 3009 5491 3043
rect 7021 3009 7055 3043
rect 7665 3009 7699 3043
rect 7757 3009 7791 3043
rect 8309 3009 8343 3043
rect 8953 3009 8987 3043
rect 12173 3009 12207 3043
rect 13185 3009 13219 3043
rect 16313 3009 16347 3043
rect 18061 3009 18095 3043
rect 22201 3009 22235 3043
rect 22845 3009 22879 3043
rect 23305 3009 23339 3043
rect 23949 3009 23983 3043
rect 24777 3009 24811 3043
rect 25421 3009 25455 3043
rect 25881 3009 25915 3043
rect 27169 3009 27203 3043
rect 33609 3009 33643 3043
rect 36921 3009 36955 3043
rect 37657 3009 37691 3043
rect 38301 3009 38335 3043
rect 9229 2941 9263 2975
rect 16957 2941 16991 2975
rect 17233 2941 17267 2975
rect 18797 2941 18831 2975
rect 19073 2941 19107 2975
rect 25973 2941 26007 2975
rect 4077 2873 4111 2907
rect 7113 2873 7147 2907
rect 10701 2873 10735 2907
rect 22017 2873 22051 2907
rect 24593 2873 24627 2907
rect 36737 2873 36771 2907
rect 38117 2873 38151 2907
rect 1777 2805 1811 2839
rect 2697 2805 2731 2839
rect 4721 2805 4755 2839
rect 8401 2805 8435 2839
rect 14933 2805 14967 2839
rect 23397 2805 23431 2839
rect 24041 2805 24075 2839
rect 25237 2805 25271 2839
rect 33793 2805 33827 2839
rect 1777 2601 1811 2635
rect 10333 2601 10367 2635
rect 11897 2601 11931 2635
rect 14552 2601 14586 2635
rect 16037 2601 16071 2635
rect 16957 2601 16991 2635
rect 19533 2601 19567 2635
rect 20453 2601 20487 2635
rect 21189 2601 21223 2635
rect 22017 2601 22051 2635
rect 27813 2601 27847 2635
rect 28641 2601 28675 2635
rect 30481 2601 30515 2635
rect 3249 2533 3283 2567
rect 9689 2533 9723 2567
rect 18429 2533 18463 2567
rect 23397 2533 23431 2567
rect 14289 2465 14323 2499
rect 20269 2465 20303 2499
rect 32597 2465 32631 2499
rect 2329 2397 2363 2431
rect 3065 2397 3099 2431
rect 4169 2397 4203 2431
rect 4629 2397 4663 2431
rect 5273 2397 5307 2431
rect 7113 2397 7147 2431
rect 7757 2397 7791 2431
rect 8401 2397 8435 2431
rect 9589 2399 9623 2433
rect 10241 2397 10275 2431
rect 10885 2397 10919 2431
rect 12817 2397 12851 2431
rect 13461 2397 13495 2431
rect 16865 2397 16899 2431
rect 17509 2397 17543 2431
rect 18245 2397 18279 2431
rect 19441 2397 19475 2431
rect 20085 2397 20119 2431
rect 21373 2397 21407 2431
rect 22201 2397 22235 2431
rect 22661 2397 22695 2431
rect 23581 2397 23615 2431
rect 24593 2397 24627 2431
rect 25237 2397 25271 2431
rect 25973 2397 26007 2431
rect 27353 2397 27387 2431
rect 27997 2397 28031 2431
rect 29745 2397 29779 2431
rect 30665 2397 30699 2431
rect 32321 2397 32355 2431
rect 33609 2397 33643 2431
rect 34897 2397 34931 2431
rect 36185 2397 36219 2431
rect 38025 2397 38059 2431
rect 1685 2329 1719 2363
rect 7205 2329 7239 2363
rect 11805 2329 11839 2363
rect 28549 2329 28583 2363
rect 2513 2261 2547 2295
rect 3985 2261 4019 2295
rect 4721 2261 4755 2295
rect 5457 2261 5491 2295
rect 7849 2261 7883 2295
rect 8493 2261 8527 2295
rect 11069 2261 11103 2295
rect 12909 2261 12943 2295
rect 13645 2261 13679 2295
rect 17693 2261 17727 2295
rect 22845 2261 22879 2295
rect 24685 2261 24719 2295
rect 25421 2261 25455 2295
rect 26157 2261 26191 2295
rect 27169 2261 27203 2295
rect 29929 2261 29963 2295
rect 33793 2261 33827 2295
rect 35081 2261 35115 2295
rect 36369 2261 36403 2295
rect 38209 2261 38243 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 1762 37448 1768 37460
rect 1723 37420 1768 37448
rect 1762 37408 1768 37420
rect 1820 37408 1826 37460
rect 18506 37272 18512 37324
rect 18564 37312 18570 37324
rect 18877 37315 18935 37321
rect 18877 37312 18889 37315
rect 18564 37284 18889 37312
rect 18564 37272 18570 37284
rect 18877 37281 18889 37284
rect 18923 37281 18935 37315
rect 18877 37275 18935 37281
rect 21266 37272 21272 37324
rect 21324 37312 21330 37324
rect 22005 37315 22063 37321
rect 22005 37312 22017 37315
rect 21324 37284 22017 37312
rect 21324 37272 21330 37284
rect 22005 37281 22017 37284
rect 22051 37281 22063 37315
rect 22005 37275 22063 37281
rect 27433 37315 27491 37321
rect 27433 37281 27445 37315
rect 27479 37312 27491 37315
rect 32766 37312 32772 37324
rect 27479 37284 32772 37312
rect 27479 37281 27491 37284
rect 27433 37275 27491 37281
rect 32766 37272 32772 37284
rect 32824 37272 32830 37324
rect 1581 37247 1639 37253
rect 1581 37213 1593 37247
rect 1627 37244 1639 37247
rect 2406 37244 2412 37256
rect 1627 37216 2412 37244
rect 1627 37213 1639 37216
rect 1581 37207 1639 37213
rect 2406 37204 2412 37216
rect 2464 37204 2470 37256
rect 2774 37204 2780 37256
rect 2832 37244 2838 37256
rect 2869 37247 2927 37253
rect 2869 37244 2881 37247
rect 2832 37216 2881 37244
rect 2832 37204 2838 37216
rect 2869 37213 2881 37216
rect 2915 37213 2927 37247
rect 3970 37244 3976 37256
rect 3931 37216 3976 37244
rect 2869 37207 2927 37213
rect 3970 37204 3976 37216
rect 4028 37204 4034 37256
rect 4614 37204 4620 37256
rect 4672 37244 4678 37256
rect 4893 37247 4951 37253
rect 4893 37244 4905 37247
rect 4672 37216 4905 37244
rect 4672 37204 4678 37216
rect 4893 37213 4905 37216
rect 4939 37213 4951 37247
rect 4893 37207 4951 37213
rect 5810 37204 5816 37256
rect 5868 37244 5874 37256
rect 5997 37247 6055 37253
rect 5997 37244 6009 37247
rect 5868 37216 6009 37244
rect 5868 37204 5874 37216
rect 5997 37213 6009 37216
rect 6043 37213 6055 37247
rect 5997 37207 6055 37213
rect 6454 37204 6460 37256
rect 6512 37244 6518 37256
rect 6733 37247 6791 37253
rect 6733 37244 6745 37247
rect 6512 37216 6745 37244
rect 6512 37204 6518 37216
rect 6733 37213 6745 37216
rect 6779 37213 6791 37247
rect 7834 37244 7840 37256
rect 7795 37216 7840 37244
rect 6733 37207 6791 37213
rect 7834 37204 7840 37216
rect 7892 37204 7898 37256
rect 9766 37244 9772 37256
rect 9727 37216 9772 37244
rect 9766 37204 9772 37216
rect 9824 37204 9830 37256
rect 11701 37247 11759 37253
rect 11701 37213 11713 37247
rect 11747 37213 11759 37247
rect 11701 37207 11759 37213
rect 6822 37176 6828 37188
rect 2700 37148 6828 37176
rect 2700 37117 2728 37148
rect 6822 37136 6828 37148
rect 6880 37136 6886 37188
rect 9490 37136 9496 37188
rect 9548 37176 9554 37188
rect 11716 37176 11744 37207
rect 12434 37204 12440 37256
rect 12492 37244 12498 37256
rect 12621 37247 12679 37253
rect 12621 37244 12633 37247
rect 12492 37216 12633 37244
rect 12492 37204 12498 37216
rect 12621 37213 12633 37216
rect 12667 37213 12679 37247
rect 12621 37207 12679 37213
rect 13725 37247 13783 37253
rect 13725 37213 13737 37247
rect 13771 37244 13783 37247
rect 14182 37244 14188 37256
rect 13771 37216 14188 37244
rect 13771 37213 13783 37216
rect 13725 37207 13783 37213
rect 14182 37204 14188 37216
rect 14240 37204 14246 37256
rect 14274 37204 14280 37256
rect 14332 37244 14338 37256
rect 14332 37216 14377 37244
rect 14332 37204 14338 37216
rect 14826 37204 14832 37256
rect 14884 37244 14890 37256
rect 15565 37247 15623 37253
rect 15565 37244 15577 37247
rect 14884 37216 15577 37244
rect 14884 37204 14890 37216
rect 15565 37213 15577 37216
rect 15611 37213 15623 37247
rect 15565 37207 15623 37213
rect 17497 37247 17555 37253
rect 17497 37213 17509 37247
rect 17543 37213 17555 37247
rect 18690 37244 18696 37256
rect 18651 37216 18696 37244
rect 17497 37207 17555 37213
rect 9548 37148 11744 37176
rect 17512 37176 17540 37207
rect 18690 37204 18696 37216
rect 18748 37204 18754 37256
rect 20070 37244 20076 37256
rect 20031 37216 20076 37244
rect 20070 37204 20076 37216
rect 20128 37204 20134 37256
rect 21450 37204 21456 37256
rect 21508 37244 21514 37256
rect 22281 37247 22339 37253
rect 22281 37244 22293 37247
rect 21508 37216 22293 37244
rect 21508 37204 21514 37216
rect 22281 37213 22293 37216
rect 22327 37213 22339 37247
rect 22281 37207 22339 37213
rect 24581 37247 24639 37253
rect 24581 37213 24593 37247
rect 24627 37213 24639 37247
rect 24581 37207 24639 37213
rect 19058 37176 19064 37188
rect 17512 37148 19064 37176
rect 9548 37136 9554 37148
rect 19058 37136 19064 37148
rect 19116 37136 19122 37188
rect 21818 37136 21824 37188
rect 21876 37176 21882 37188
rect 24596 37176 24624 37207
rect 25130 37204 25136 37256
rect 25188 37244 25194 37256
rect 25501 37247 25559 37253
rect 25501 37244 25513 37247
rect 25188 37216 25513 37244
rect 25188 37204 25194 37216
rect 25501 37213 25513 37216
rect 25547 37213 25559 37247
rect 25501 37207 25559 37213
rect 26418 37204 26424 37256
rect 26476 37244 26482 37256
rect 27249 37247 27307 37253
rect 27249 37244 27261 37247
rect 26476 37216 27261 37244
rect 26476 37204 26482 37216
rect 27249 37213 27261 37216
rect 27295 37213 27307 37247
rect 27890 37244 27896 37256
rect 27851 37216 27896 37244
rect 27249 37207 27307 37213
rect 27890 37204 27896 37216
rect 27948 37204 27954 37256
rect 28350 37204 28356 37256
rect 28408 37244 28414 37256
rect 28813 37247 28871 37253
rect 28813 37244 28825 37247
rect 28408 37216 28825 37244
rect 28408 37204 28414 37216
rect 28813 37213 28825 37216
rect 28859 37213 28871 37247
rect 28813 37207 28871 37213
rect 29638 37204 29644 37256
rect 29696 37244 29702 37256
rect 29917 37247 29975 37253
rect 29917 37244 29929 37247
rect 29696 37216 29929 37244
rect 29696 37204 29702 37216
rect 29917 37213 29929 37216
rect 29963 37213 29975 37247
rect 29917 37207 29975 37213
rect 30926 37204 30932 37256
rect 30984 37244 30990 37256
rect 31205 37247 31263 37253
rect 31205 37244 31217 37247
rect 30984 37216 31217 37244
rect 30984 37204 30990 37216
rect 31205 37213 31217 37216
rect 31251 37213 31263 37247
rect 32306 37244 32312 37256
rect 32267 37216 32312 37244
rect 31205 37207 31263 37213
rect 32306 37204 32312 37216
rect 32364 37204 32370 37256
rect 32398 37204 32404 37256
rect 32456 37244 32462 37256
rect 33045 37247 33103 37253
rect 33045 37244 33057 37247
rect 32456 37216 33057 37244
rect 32456 37204 32462 37216
rect 33045 37213 33057 37216
rect 33091 37213 33103 37247
rect 33045 37207 33103 37213
rect 34790 37204 34796 37256
rect 34848 37244 34854 37256
rect 34885 37247 34943 37253
rect 34885 37244 34897 37247
rect 34848 37216 34897 37244
rect 34848 37204 34854 37216
rect 34885 37213 34897 37216
rect 34931 37244 34943 37247
rect 35437 37247 35495 37253
rect 35437 37244 35449 37247
rect 34931 37216 35449 37244
rect 34931 37213 34943 37216
rect 34885 37207 34943 37213
rect 35437 37213 35449 37216
rect 35483 37244 35495 37247
rect 35805 37247 35863 37253
rect 35805 37244 35817 37247
rect 35483 37216 35817 37244
rect 35483 37213 35495 37216
rect 35437 37207 35495 37213
rect 35805 37213 35817 37216
rect 35851 37213 35863 37247
rect 35805 37207 35863 37213
rect 36078 37204 36084 37256
rect 36136 37244 36142 37256
rect 36265 37247 36323 37253
rect 36265 37244 36277 37247
rect 36136 37216 36277 37244
rect 36136 37204 36142 37216
rect 36265 37213 36277 37216
rect 36311 37213 36323 37247
rect 36265 37207 36323 37213
rect 37366 37204 37372 37256
rect 37424 37244 37430 37256
rect 37553 37247 37611 37253
rect 37553 37244 37565 37247
rect 37424 37216 37565 37244
rect 37424 37204 37430 37216
rect 37553 37213 37565 37216
rect 37599 37213 37611 37247
rect 37553 37207 37611 37213
rect 21876 37148 24624 37176
rect 21876 37136 21882 37148
rect 28258 37136 28264 37188
rect 28316 37176 28322 37188
rect 28316 37148 31064 37176
rect 28316 37136 28322 37148
rect 2685 37111 2743 37117
rect 2685 37077 2697 37111
rect 2731 37077 2743 37111
rect 2685 37071 2743 37077
rect 3234 37068 3240 37120
rect 3292 37108 3298 37120
rect 4157 37111 4215 37117
rect 4157 37108 4169 37111
rect 3292 37080 4169 37108
rect 3292 37068 3298 37080
rect 4157 37077 4169 37080
rect 4203 37077 4215 37111
rect 4706 37108 4712 37120
rect 4667 37080 4712 37108
rect 4157 37071 4215 37077
rect 4706 37068 4712 37080
rect 4764 37068 4770 37120
rect 5813 37111 5871 37117
rect 5813 37077 5825 37111
rect 5859 37108 5871 37111
rect 6362 37108 6368 37120
rect 5859 37080 6368 37108
rect 5859 37077 5871 37080
rect 5813 37071 5871 37077
rect 6362 37068 6368 37080
rect 6420 37068 6426 37120
rect 6546 37108 6552 37120
rect 6507 37080 6552 37108
rect 6546 37068 6552 37080
rect 6604 37068 6610 37120
rect 7742 37068 7748 37120
rect 7800 37108 7806 37120
rect 8021 37111 8079 37117
rect 8021 37108 8033 37111
rect 7800 37080 8033 37108
rect 7800 37068 7806 37080
rect 8021 37077 8033 37080
rect 8067 37077 8079 37111
rect 8021 37071 8079 37077
rect 9674 37068 9680 37120
rect 9732 37108 9738 37120
rect 9953 37111 10011 37117
rect 9953 37108 9965 37111
rect 9732 37080 9965 37108
rect 9732 37068 9738 37080
rect 9953 37077 9965 37080
rect 9999 37077 10011 37111
rect 9953 37071 10011 37077
rect 11054 37068 11060 37120
rect 11112 37108 11118 37120
rect 11885 37111 11943 37117
rect 11885 37108 11897 37111
rect 11112 37080 11897 37108
rect 11112 37068 11118 37080
rect 11885 37077 11897 37080
rect 11931 37077 11943 37111
rect 12434 37108 12440 37120
rect 12395 37080 12440 37108
rect 11885 37071 11943 37077
rect 12434 37068 12440 37080
rect 12492 37068 12498 37120
rect 12894 37068 12900 37120
rect 12952 37108 12958 37120
rect 13541 37111 13599 37117
rect 13541 37108 13553 37111
rect 12952 37080 13553 37108
rect 12952 37068 12958 37080
rect 13541 37077 13553 37080
rect 13587 37077 13599 37111
rect 13541 37071 13599 37077
rect 13814 37068 13820 37120
rect 13872 37108 13878 37120
rect 14461 37111 14519 37117
rect 14461 37108 14473 37111
rect 13872 37080 14473 37108
rect 13872 37068 13878 37080
rect 14461 37077 14473 37080
rect 14507 37077 14519 37111
rect 14461 37071 14519 37077
rect 15470 37068 15476 37120
rect 15528 37108 15534 37120
rect 15749 37111 15807 37117
rect 15749 37108 15761 37111
rect 15528 37080 15761 37108
rect 15528 37068 15534 37080
rect 15749 37077 15761 37080
rect 15795 37077 15807 37111
rect 15749 37071 15807 37077
rect 17402 37068 17408 37120
rect 17460 37108 17466 37120
rect 17681 37111 17739 37117
rect 17681 37108 17693 37111
rect 17460 37080 17693 37108
rect 17460 37068 17466 37080
rect 17681 37077 17693 37080
rect 17727 37077 17739 37111
rect 17681 37071 17739 37077
rect 19978 37068 19984 37120
rect 20036 37108 20042 37120
rect 20257 37111 20315 37117
rect 20257 37108 20269 37111
rect 20036 37080 20269 37108
rect 20036 37068 20042 37080
rect 20257 37077 20269 37080
rect 20303 37077 20315 37111
rect 20257 37071 20315 37077
rect 24486 37068 24492 37120
rect 24544 37108 24550 37120
rect 24765 37111 24823 37117
rect 24765 37108 24777 37111
rect 24544 37080 24777 37108
rect 24544 37068 24550 37080
rect 24765 37077 24777 37080
rect 24811 37077 24823 37111
rect 25314 37108 25320 37120
rect 25275 37080 25320 37108
rect 24765 37071 24823 37077
rect 25314 37068 25320 37080
rect 25372 37068 25378 37120
rect 27706 37068 27712 37120
rect 27764 37108 27770 37120
rect 28077 37111 28135 37117
rect 28077 37108 28089 37111
rect 27764 37080 28089 37108
rect 27764 37068 27770 37080
rect 28077 37077 28089 37080
rect 28123 37077 28135 37111
rect 28626 37108 28632 37120
rect 28587 37080 28632 37108
rect 28077 37071 28135 37077
rect 28626 37068 28632 37080
rect 28684 37068 28690 37120
rect 28718 37068 28724 37120
rect 28776 37108 28782 37120
rect 31036 37117 31064 37148
rect 29733 37111 29791 37117
rect 29733 37108 29745 37111
rect 28776 37080 29745 37108
rect 28776 37068 28782 37080
rect 29733 37077 29745 37080
rect 29779 37077 29791 37111
rect 29733 37071 29791 37077
rect 31021 37111 31079 37117
rect 31021 37077 31033 37111
rect 31067 37077 31079 37111
rect 31021 37071 31079 37077
rect 32214 37068 32220 37120
rect 32272 37108 32278 37120
rect 32493 37111 32551 37117
rect 32493 37108 32505 37111
rect 32272 37080 32505 37108
rect 32272 37068 32278 37080
rect 32493 37077 32505 37080
rect 32539 37077 32551 37111
rect 32493 37071 32551 37077
rect 33134 37068 33140 37120
rect 33192 37108 33198 37120
rect 33229 37111 33287 37117
rect 33229 37108 33241 37111
rect 33192 37080 33241 37108
rect 33192 37068 33198 37080
rect 33229 37077 33241 37080
rect 33275 37077 33287 37111
rect 33229 37071 33287 37077
rect 34514 37068 34520 37120
rect 34572 37108 34578 37120
rect 35069 37111 35127 37117
rect 35069 37108 35081 37111
rect 34572 37080 35081 37108
rect 34572 37068 34578 37080
rect 35069 37077 35081 37080
rect 35115 37077 35127 37111
rect 36354 37108 36360 37120
rect 36315 37080 36360 37108
rect 35069 37071 35127 37077
rect 36354 37068 36360 37080
rect 36412 37068 36418 37120
rect 37642 37108 37648 37120
rect 37603 37080 37648 37108
rect 37642 37068 37648 37080
rect 37700 37068 37706 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 1670 36864 1676 36916
rect 1728 36904 1734 36916
rect 1765 36907 1823 36913
rect 1765 36904 1777 36907
rect 1728 36876 1777 36904
rect 1728 36864 1734 36876
rect 1765 36873 1777 36876
rect 1811 36873 1823 36907
rect 1765 36867 1823 36873
rect 9030 36864 9036 36916
rect 9088 36904 9094 36916
rect 9309 36907 9367 36913
rect 9309 36904 9321 36907
rect 9088 36876 9321 36904
rect 9088 36864 9094 36876
rect 9309 36873 9321 36876
rect 9355 36873 9367 36907
rect 14826 36904 14832 36916
rect 14787 36876 14832 36904
rect 9309 36867 9367 36873
rect 14826 36864 14832 36876
rect 14884 36864 14890 36916
rect 16758 36864 16764 36916
rect 16816 36904 16822 36916
rect 17037 36907 17095 36913
rect 17037 36904 17049 36907
rect 16816 36876 17049 36904
rect 16816 36864 16822 36876
rect 17037 36873 17049 36876
rect 17083 36873 17095 36907
rect 22830 36904 22836 36916
rect 17037 36867 17095 36873
rect 17144 36876 22836 36904
rect 14 36796 20 36848
rect 72 36836 78 36848
rect 72 36808 3188 36836
rect 72 36796 78 36808
rect 1581 36771 1639 36777
rect 1581 36737 1593 36771
rect 1627 36737 1639 36771
rect 2498 36768 2504 36780
rect 2459 36740 2504 36768
rect 1581 36731 1639 36737
rect 1596 36700 1624 36731
rect 2498 36728 2504 36740
rect 2556 36728 2562 36780
rect 3160 36777 3188 36808
rect 7834 36796 7840 36848
rect 7892 36836 7898 36848
rect 17144 36836 17172 36876
rect 22830 36864 22836 36876
rect 22888 36864 22894 36916
rect 27157 36907 27215 36913
rect 27157 36873 27169 36907
rect 27203 36904 27215 36907
rect 32306 36904 32312 36916
rect 27203 36876 32312 36904
rect 27203 36873 27215 36876
rect 27157 36867 27215 36873
rect 32306 36864 32312 36876
rect 32364 36864 32370 36916
rect 7892 36808 17172 36836
rect 7892 36796 7898 36808
rect 19334 36796 19340 36848
rect 19392 36836 19398 36848
rect 38102 36836 38108 36848
rect 19392 36808 35894 36836
rect 38063 36808 38108 36836
rect 19392 36796 19398 36808
rect 3145 36771 3203 36777
rect 3145 36737 3157 36771
rect 3191 36737 3203 36771
rect 9122 36768 9128 36780
rect 9083 36740 9128 36768
rect 3145 36731 3203 36737
rect 9122 36728 9128 36740
rect 9180 36728 9186 36780
rect 14090 36768 14096 36780
rect 14051 36740 14096 36768
rect 14090 36728 14096 36740
rect 14148 36728 14154 36780
rect 14185 36771 14243 36777
rect 14185 36737 14197 36771
rect 14231 36768 14243 36771
rect 15013 36771 15071 36777
rect 15013 36768 15025 36771
rect 14231 36740 15025 36768
rect 14231 36737 14243 36740
rect 14185 36731 14243 36737
rect 15013 36737 15025 36740
rect 15059 36737 15071 36771
rect 16850 36768 16856 36780
rect 16811 36740 16856 36768
rect 15013 36731 15071 36737
rect 16850 36728 16856 36740
rect 16908 36728 16914 36780
rect 17865 36771 17923 36777
rect 17865 36737 17877 36771
rect 17911 36768 17923 36771
rect 19352 36768 19380 36796
rect 17911 36740 19380 36768
rect 17911 36737 17923 36740
rect 17865 36731 17923 36737
rect 22094 36728 22100 36780
rect 22152 36768 22158 36780
rect 22189 36771 22247 36777
rect 22189 36768 22201 36771
rect 22152 36740 22201 36768
rect 22152 36728 22158 36740
rect 22189 36737 22201 36740
rect 22235 36737 22247 36771
rect 22189 36731 22247 36737
rect 23198 36728 23204 36780
rect 23256 36768 23262 36780
rect 23293 36771 23351 36777
rect 23293 36768 23305 36771
rect 23256 36740 23305 36768
rect 23256 36728 23262 36740
rect 23293 36737 23305 36740
rect 23339 36737 23351 36771
rect 27341 36771 27399 36777
rect 27341 36768 27353 36771
rect 23293 36731 23351 36737
rect 26206 36740 27353 36768
rect 4062 36700 4068 36712
rect 1596 36672 4068 36700
rect 4062 36660 4068 36672
rect 4120 36660 4126 36712
rect 23569 36703 23627 36709
rect 23569 36700 23581 36703
rect 22112 36672 23581 36700
rect 22112 36644 22140 36672
rect 23569 36669 23581 36672
rect 23615 36700 23627 36703
rect 26206 36700 26234 36740
rect 27341 36737 27353 36740
rect 27387 36737 27399 36771
rect 27341 36731 27399 36737
rect 35434 36728 35440 36780
rect 35492 36768 35498 36780
rect 35713 36771 35771 36777
rect 35713 36768 35725 36771
rect 35492 36740 35725 36768
rect 35492 36728 35498 36740
rect 35713 36737 35725 36740
rect 35759 36737 35771 36771
rect 35713 36731 35771 36737
rect 23615 36672 26234 36700
rect 35866 36700 35894 36808
rect 38102 36796 38108 36808
rect 38160 36796 38166 36848
rect 36909 36771 36967 36777
rect 36909 36737 36921 36771
rect 36955 36768 36967 36771
rect 39298 36768 39304 36780
rect 36955 36740 39304 36768
rect 36955 36737 36967 36740
rect 36909 36731 36967 36737
rect 39298 36728 39304 36740
rect 39356 36728 39362 36780
rect 37642 36700 37648 36712
rect 35866 36672 37648 36700
rect 23615 36669 23627 36672
rect 23569 36663 23627 36669
rect 37642 36660 37648 36672
rect 37700 36660 37706 36712
rect 14274 36592 14280 36644
rect 14332 36632 14338 36644
rect 17681 36635 17739 36641
rect 17681 36632 17693 36635
rect 14332 36604 17693 36632
rect 14332 36592 14338 36604
rect 17681 36601 17693 36604
rect 17727 36601 17739 36635
rect 17681 36595 17739 36601
rect 22094 36592 22100 36644
rect 22152 36592 22158 36644
rect 33134 36592 33140 36644
rect 33192 36632 33198 36644
rect 36725 36635 36783 36641
rect 36725 36632 36737 36635
rect 33192 36604 36737 36632
rect 33192 36592 33198 36604
rect 36725 36601 36737 36604
rect 36771 36601 36783 36635
rect 36725 36595 36783 36601
rect 38289 36635 38347 36641
rect 38289 36601 38301 36635
rect 38335 36632 38347 36635
rect 38378 36632 38384 36644
rect 38335 36604 38384 36632
rect 38335 36601 38347 36604
rect 38289 36595 38347 36601
rect 38378 36592 38384 36604
rect 38436 36592 38442 36644
rect 2314 36564 2320 36576
rect 2275 36536 2320 36564
rect 2314 36524 2320 36536
rect 2372 36524 2378 36576
rect 2961 36567 3019 36573
rect 2961 36533 2973 36567
rect 3007 36564 3019 36567
rect 5810 36564 5816 36576
rect 3007 36536 5816 36564
rect 3007 36533 3019 36536
rect 2961 36527 3019 36533
rect 5810 36524 5816 36536
rect 5868 36524 5874 36576
rect 20714 36524 20720 36576
rect 20772 36564 20778 36576
rect 22005 36567 22063 36573
rect 22005 36564 22017 36567
rect 20772 36536 22017 36564
rect 20772 36524 20778 36536
rect 22005 36533 22017 36536
rect 22051 36533 22063 36567
rect 35526 36564 35532 36576
rect 35487 36536 35532 36564
rect 22005 36527 22063 36533
rect 35526 36524 35532 36536
rect 35584 36524 35590 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 19705 36363 19763 36369
rect 19705 36329 19717 36363
rect 19751 36360 19763 36363
rect 20070 36360 20076 36372
rect 19751 36332 20076 36360
rect 19751 36329 19763 36332
rect 19705 36323 19763 36329
rect 20070 36320 20076 36332
rect 20128 36320 20134 36372
rect 37182 36320 37188 36372
rect 37240 36360 37246 36372
rect 37461 36363 37519 36369
rect 37461 36360 37473 36363
rect 37240 36332 37473 36360
rect 37240 36320 37246 36332
rect 37461 36329 37473 36332
rect 37507 36329 37519 36363
rect 37461 36323 37519 36329
rect 27614 36184 27620 36236
rect 27672 36224 27678 36236
rect 28718 36224 28724 36236
rect 27672 36196 28724 36224
rect 27672 36184 27678 36196
rect 28718 36184 28724 36196
rect 28776 36184 28782 36236
rect 38470 36224 38476 36236
rect 37292 36196 38476 36224
rect 1302 36116 1308 36168
rect 1360 36156 1366 36168
rect 1765 36159 1823 36165
rect 1765 36156 1777 36159
rect 1360 36128 1777 36156
rect 1360 36116 1366 36128
rect 1765 36125 1777 36128
rect 1811 36125 1823 36159
rect 1765 36119 1823 36125
rect 19889 36159 19947 36165
rect 19889 36125 19901 36159
rect 19935 36156 19947 36159
rect 19978 36156 19984 36168
rect 19935 36128 19984 36156
rect 19935 36125 19947 36128
rect 19889 36119 19947 36125
rect 19978 36116 19984 36128
rect 20036 36116 20042 36168
rect 37292 36165 37320 36196
rect 38470 36184 38476 36196
rect 38528 36184 38534 36236
rect 37277 36159 37335 36165
rect 37277 36125 37289 36159
rect 37323 36125 37335 36159
rect 37277 36119 37335 36125
rect 38013 36159 38071 36165
rect 38013 36125 38025 36159
rect 38059 36125 38071 36159
rect 38013 36119 38071 36125
rect 33226 36048 33232 36100
rect 33284 36088 33290 36100
rect 38028 36088 38056 36119
rect 33284 36060 38056 36088
rect 33284 36048 33290 36060
rect 1581 36023 1639 36029
rect 1581 35989 1593 36023
rect 1627 36020 1639 36023
rect 2590 36020 2596 36032
rect 1627 35992 2596 36020
rect 1627 35989 1639 35992
rect 1581 35983 1639 35989
rect 2590 35980 2596 35992
rect 2648 35980 2654 36032
rect 38194 36020 38200 36032
rect 38155 35992 38200 36020
rect 38194 35980 38200 35992
rect 38252 35980 38258 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 38102 35680 38108 35692
rect 38063 35652 38108 35680
rect 38102 35640 38108 35652
rect 38160 35640 38166 35692
rect 1578 35612 1584 35624
rect 1539 35584 1584 35612
rect 1578 35572 1584 35584
rect 1636 35572 1642 35624
rect 1857 35615 1915 35621
rect 1857 35581 1869 35615
rect 1903 35612 1915 35615
rect 7466 35612 7472 35624
rect 1903 35584 7472 35612
rect 1903 35581 1915 35584
rect 1857 35575 1915 35581
rect 7466 35572 7472 35584
rect 7524 35572 7530 35624
rect 37642 35436 37648 35488
rect 37700 35476 37706 35488
rect 38197 35479 38255 35485
rect 38197 35476 38209 35479
rect 37700 35448 38209 35476
rect 37700 35436 37706 35448
rect 38197 35445 38209 35448
rect 38243 35445 38255 35479
rect 38197 35439 38255 35445
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 3145 35275 3203 35281
rect 3145 35241 3157 35275
rect 3191 35272 3203 35275
rect 3970 35272 3976 35284
rect 3191 35244 3976 35272
rect 3191 35241 3203 35244
rect 3145 35235 3203 35241
rect 3970 35232 3976 35244
rect 4028 35232 4034 35284
rect 19521 35275 19579 35281
rect 19521 35241 19533 35275
rect 19567 35272 19579 35275
rect 19978 35272 19984 35284
rect 19567 35244 19984 35272
rect 19567 35241 19579 35244
rect 19521 35235 19579 35241
rect 19978 35232 19984 35244
rect 20036 35232 20042 35284
rect 1762 35068 1768 35080
rect 1723 35040 1768 35068
rect 1762 35028 1768 35040
rect 1820 35028 1826 35080
rect 1854 35028 1860 35080
rect 1912 35068 1918 35080
rect 3329 35071 3387 35077
rect 3329 35068 3341 35071
rect 1912 35040 3341 35068
rect 1912 35028 1918 35040
rect 3329 35037 3341 35040
rect 3375 35037 3387 35071
rect 19426 35068 19432 35080
rect 19387 35040 19432 35068
rect 3329 35031 3387 35037
rect 19426 35028 19432 35040
rect 19484 35028 19490 35080
rect 38289 35071 38347 35077
rect 38289 35037 38301 35071
rect 38335 35068 38347 35071
rect 38654 35068 38660 35080
rect 38335 35040 38660 35068
rect 38335 35037 38347 35040
rect 38289 35031 38347 35037
rect 38654 35028 38660 35040
rect 38712 35028 38718 35080
rect 1581 34935 1639 34941
rect 1581 34901 1593 34935
rect 1627 34932 1639 34935
rect 2682 34932 2688 34944
rect 1627 34904 2688 34932
rect 1627 34901 1639 34904
rect 1581 34895 1639 34901
rect 2682 34892 2688 34904
rect 2740 34892 2746 34944
rect 37274 34892 37280 34944
rect 37332 34932 37338 34944
rect 38105 34935 38163 34941
rect 38105 34932 38117 34935
rect 37332 34904 38117 34932
rect 37332 34892 37338 34904
rect 38105 34901 38117 34904
rect 38151 34901 38163 34935
rect 38105 34895 38163 34901
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 4062 34688 4068 34740
rect 4120 34728 4126 34740
rect 4341 34731 4399 34737
rect 4341 34728 4353 34731
rect 4120 34700 4353 34728
rect 4120 34688 4126 34700
rect 4341 34697 4353 34700
rect 4387 34697 4399 34731
rect 4341 34691 4399 34697
rect 4525 34595 4583 34601
rect 4525 34561 4537 34595
rect 4571 34592 4583 34595
rect 5718 34592 5724 34604
rect 4571 34564 5724 34592
rect 4571 34561 4583 34564
rect 4525 34555 4583 34561
rect 5718 34552 5724 34564
rect 5776 34552 5782 34604
rect 38013 34595 38071 34601
rect 38013 34561 38025 34595
rect 38059 34592 38071 34595
rect 38562 34592 38568 34604
rect 38059 34564 38568 34592
rect 38059 34561 38071 34564
rect 38013 34555 38071 34561
rect 38562 34552 38568 34564
rect 38620 34552 38626 34604
rect 38194 34388 38200 34400
rect 38155 34360 38200 34388
rect 38194 34348 38200 34360
rect 38252 34348 38258 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 21818 34144 21824 34196
rect 21876 34184 21882 34196
rect 22005 34187 22063 34193
rect 22005 34184 22017 34187
rect 21876 34156 22017 34184
rect 21876 34144 21882 34156
rect 22005 34153 22017 34156
rect 22051 34153 22063 34187
rect 22005 34147 22063 34153
rect 21358 33940 21364 33992
rect 21416 33980 21422 33992
rect 22189 33983 22247 33989
rect 22189 33980 22201 33983
rect 21416 33952 22201 33980
rect 21416 33940 21422 33952
rect 22189 33949 22201 33952
rect 22235 33949 22247 33983
rect 22189 33943 22247 33949
rect 2406 33804 2412 33856
rect 2464 33844 2470 33856
rect 17402 33844 17408 33856
rect 2464 33816 17408 33844
rect 2464 33804 2470 33816
rect 17402 33804 17408 33816
rect 17460 33804 17466 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 1581 33507 1639 33513
rect 1581 33473 1593 33507
rect 1627 33504 1639 33507
rect 4062 33504 4068 33516
rect 1627 33476 4068 33504
rect 1627 33473 1639 33476
rect 1581 33467 1639 33473
rect 4062 33464 4068 33476
rect 4120 33464 4126 33516
rect 4706 33464 4712 33516
rect 4764 33504 4770 33516
rect 8573 33507 8631 33513
rect 8573 33504 8585 33507
rect 4764 33476 8585 33504
rect 4764 33464 4770 33476
rect 8573 33473 8585 33476
rect 8619 33473 8631 33507
rect 8573 33467 8631 33473
rect 1762 33368 1768 33380
rect 1723 33340 1768 33368
rect 1762 33328 1768 33340
rect 1820 33328 1826 33380
rect 8665 33303 8723 33309
rect 8665 33269 8677 33303
rect 8711 33300 8723 33303
rect 9306 33300 9312 33312
rect 8711 33272 9312 33300
rect 8711 33269 8723 33272
rect 8665 33263 8723 33269
rect 9306 33260 9312 33272
rect 9364 33260 9370 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 33226 33096 33232 33108
rect 33187 33068 33232 33096
rect 33226 33056 33232 33068
rect 33284 33056 33290 33108
rect 6546 32852 6552 32904
rect 6604 32892 6610 32904
rect 9585 32895 9643 32901
rect 9585 32892 9597 32895
rect 6604 32864 9597 32892
rect 6604 32852 6610 32864
rect 9585 32861 9597 32864
rect 9631 32861 9643 32895
rect 9585 32855 9643 32861
rect 11057 32895 11115 32901
rect 11057 32861 11069 32895
rect 11103 32892 11115 32895
rect 13630 32892 13636 32904
rect 11103 32864 13636 32892
rect 11103 32861 11115 32864
rect 11057 32855 11115 32861
rect 13630 32852 13636 32864
rect 13688 32852 13694 32904
rect 28258 32892 28264 32904
rect 28219 32864 28264 32892
rect 28258 32852 28264 32864
rect 28316 32852 28322 32904
rect 30466 32852 30472 32904
rect 30524 32892 30530 32904
rect 33413 32895 33471 32901
rect 33413 32892 33425 32895
rect 30524 32864 33425 32892
rect 30524 32852 30530 32864
rect 33413 32861 33425 32864
rect 33459 32861 33471 32895
rect 33413 32855 33471 32861
rect 38102 32824 38108 32836
rect 38063 32796 38108 32824
rect 38102 32784 38108 32796
rect 38160 32784 38166 32836
rect 9677 32759 9735 32765
rect 9677 32725 9689 32759
rect 9723 32756 9735 32759
rect 10134 32756 10140 32768
rect 9723 32728 10140 32756
rect 9723 32725 9735 32728
rect 9677 32719 9735 32725
rect 10134 32716 10140 32728
rect 10192 32716 10198 32768
rect 10778 32716 10784 32768
rect 10836 32756 10842 32768
rect 11149 32759 11207 32765
rect 11149 32756 11161 32759
rect 10836 32728 11161 32756
rect 10836 32716 10842 32728
rect 11149 32725 11161 32728
rect 11195 32725 11207 32759
rect 28350 32756 28356 32768
rect 28311 32728 28356 32756
rect 11149 32719 11207 32725
rect 28350 32716 28356 32728
rect 28408 32716 28414 32768
rect 38194 32756 38200 32768
rect 38155 32728 38200 32756
rect 38194 32716 38200 32728
rect 38252 32716 38258 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 9033 32555 9091 32561
rect 9033 32521 9045 32555
rect 9079 32552 9091 32555
rect 9490 32552 9496 32564
rect 9079 32524 9496 32552
rect 9079 32521 9091 32524
rect 9033 32515 9091 32521
rect 9490 32512 9496 32524
rect 9548 32512 9554 32564
rect 9766 32512 9772 32564
rect 9824 32552 9830 32564
rect 10597 32555 10655 32561
rect 10597 32552 10609 32555
rect 9824 32524 10609 32552
rect 9824 32512 9830 32524
rect 10597 32521 10609 32524
rect 10643 32521 10655 32555
rect 10597 32515 10655 32521
rect 1581 32419 1639 32425
rect 1581 32385 1593 32419
rect 1627 32416 1639 32419
rect 9214 32416 9220 32428
rect 1627 32388 2268 32416
rect 9175 32388 9220 32416
rect 1627 32385 1639 32388
rect 1581 32379 1639 32385
rect 2240 32224 2268 32388
rect 9214 32376 9220 32388
rect 9272 32376 9278 32428
rect 10778 32416 10784 32428
rect 10739 32388 10784 32416
rect 10778 32376 10784 32388
rect 10836 32376 10842 32428
rect 20714 32416 20720 32428
rect 20675 32388 20720 32416
rect 20714 32376 20720 32388
rect 20772 32376 20778 32428
rect 23477 32419 23535 32425
rect 23477 32385 23489 32419
rect 23523 32416 23535 32419
rect 28626 32416 28632 32428
rect 23523 32388 28632 32416
rect 23523 32385 23535 32388
rect 23477 32379 23535 32385
rect 28626 32376 28632 32388
rect 28684 32376 28690 32428
rect 38102 32416 38108 32428
rect 38063 32388 38108 32416
rect 38102 32376 38108 32388
rect 38160 32376 38166 32428
rect 1762 32212 1768 32224
rect 1723 32184 1768 32212
rect 1762 32172 1768 32184
rect 1820 32172 1826 32224
rect 2222 32212 2228 32224
rect 2183 32184 2228 32212
rect 2222 32172 2228 32184
rect 2280 32172 2286 32224
rect 20622 32172 20628 32224
rect 20680 32212 20686 32224
rect 20809 32215 20867 32221
rect 20809 32212 20821 32215
rect 20680 32184 20821 32212
rect 20680 32172 20686 32184
rect 20809 32181 20821 32184
rect 20855 32181 20867 32215
rect 23566 32212 23572 32224
rect 23527 32184 23572 32212
rect 20809 32175 20867 32181
rect 23566 32172 23572 32184
rect 23624 32172 23630 32224
rect 37918 32172 37924 32224
rect 37976 32212 37982 32224
rect 38197 32215 38255 32221
rect 38197 32212 38209 32215
rect 37976 32184 38209 32212
rect 37976 32172 37982 32184
rect 38197 32181 38209 32184
rect 38243 32181 38255 32215
rect 38197 32175 38255 32181
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 2222 31968 2228 32020
rect 2280 32008 2286 32020
rect 17218 32008 17224 32020
rect 2280 31980 17224 32008
rect 2280 31968 2286 31980
rect 17218 31968 17224 31980
rect 17276 31968 17282 32020
rect 18782 31968 18788 32020
rect 18840 32008 18846 32020
rect 24673 32011 24731 32017
rect 24673 32008 24685 32011
rect 18840 31980 24685 32008
rect 18840 31968 18846 31980
rect 24673 31977 24685 31980
rect 24719 31977 24731 32011
rect 24673 31971 24731 31977
rect 15378 31900 15384 31952
rect 15436 31940 15442 31952
rect 23566 31940 23572 31952
rect 15436 31912 23572 31940
rect 15436 31900 15442 31912
rect 23566 31900 23572 31912
rect 23624 31900 23630 31952
rect 1854 31872 1860 31884
rect 1815 31844 1860 31872
rect 1854 31832 1860 31844
rect 1912 31872 1918 31884
rect 2958 31872 2964 31884
rect 1912 31844 2964 31872
rect 1912 31832 1918 31844
rect 2958 31832 2964 31844
rect 3016 31832 3022 31884
rect 20714 31832 20720 31884
rect 20772 31872 20778 31884
rect 21453 31875 21511 31881
rect 21453 31872 21465 31875
rect 20772 31844 21465 31872
rect 20772 31832 20778 31844
rect 21453 31841 21465 31844
rect 21499 31841 21511 31875
rect 25314 31872 25320 31884
rect 21453 31835 21511 31841
rect 24504 31844 25320 31872
rect 1578 31804 1584 31816
rect 1539 31776 1584 31804
rect 1578 31764 1584 31776
rect 1636 31764 1642 31816
rect 21361 31807 21419 31813
rect 21361 31773 21373 31807
rect 21407 31804 21419 31807
rect 24504 31804 24532 31844
rect 25314 31832 25320 31844
rect 25372 31832 25378 31884
rect 27798 31832 27804 31884
rect 27856 31872 27862 31884
rect 28077 31875 28135 31881
rect 28077 31872 28089 31875
rect 27856 31844 28089 31872
rect 27856 31832 27862 31844
rect 28077 31841 28089 31844
rect 28123 31841 28135 31875
rect 28077 31835 28135 31841
rect 21407 31776 24532 31804
rect 24581 31807 24639 31813
rect 21407 31773 21419 31776
rect 21361 31767 21419 31773
rect 24581 31773 24593 31807
rect 24627 31804 24639 31807
rect 27614 31804 27620 31816
rect 24627 31776 27620 31804
rect 24627 31773 24639 31776
rect 24581 31767 24639 31773
rect 27614 31764 27620 31776
rect 27672 31764 27678 31816
rect 27985 31807 28043 31813
rect 27985 31773 27997 31807
rect 28031 31804 28043 31807
rect 35526 31804 35532 31816
rect 28031 31776 35532 31804
rect 28031 31773 28043 31776
rect 27985 31767 28043 31773
rect 35526 31764 35532 31776
rect 35584 31764 35590 31816
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 29273 31331 29331 31337
rect 29273 31297 29285 31331
rect 29319 31328 29331 31331
rect 33134 31328 33140 31340
rect 29319 31300 33140 31328
rect 29319 31297 29331 31300
rect 29273 31291 29331 31297
rect 33134 31288 33140 31300
rect 33192 31288 33198 31340
rect 17586 31084 17592 31136
rect 17644 31124 17650 31136
rect 29365 31127 29423 31133
rect 29365 31124 29377 31127
rect 17644 31096 29377 31124
rect 17644 31084 17650 31096
rect 29365 31093 29377 31096
rect 29411 31093 29423 31127
rect 29365 31087 29423 31093
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 8389 30923 8447 30929
rect 8389 30889 8401 30923
rect 8435 30920 8447 30923
rect 9214 30920 9220 30932
rect 8435 30892 9220 30920
rect 8435 30889 8447 30892
rect 8389 30883 8447 30889
rect 9214 30880 9220 30892
rect 9272 30880 9278 30932
rect 25961 30923 26019 30929
rect 25961 30889 25973 30923
rect 26007 30920 26019 30923
rect 27890 30920 27896 30932
rect 26007 30892 27896 30920
rect 26007 30889 26019 30892
rect 25961 30883 26019 30889
rect 27890 30880 27896 30892
rect 27948 30880 27954 30932
rect 5905 30855 5963 30861
rect 5905 30821 5917 30855
rect 5951 30852 5963 30855
rect 9766 30852 9772 30864
rect 5951 30824 9772 30852
rect 5951 30821 5963 30824
rect 5905 30815 5963 30821
rect 9766 30812 9772 30824
rect 9824 30812 9830 30864
rect 37274 30852 37280 30864
rect 31726 30824 37280 30852
rect 2590 30744 2596 30796
rect 2648 30784 2654 30796
rect 2648 30756 7144 30784
rect 2648 30744 2654 30756
rect 2314 30676 2320 30728
rect 2372 30716 2378 30728
rect 3973 30719 4031 30725
rect 3973 30716 3985 30719
rect 2372 30688 3985 30716
rect 2372 30676 2378 30688
rect 3973 30685 3985 30688
rect 4019 30685 4031 30719
rect 5810 30716 5816 30728
rect 5771 30688 5816 30716
rect 3973 30679 4031 30685
rect 5810 30676 5816 30688
rect 5868 30676 5874 30728
rect 6362 30676 6368 30728
rect 6420 30716 6426 30728
rect 7116 30725 7144 30756
rect 6457 30719 6515 30725
rect 6457 30716 6469 30719
rect 6420 30688 6469 30716
rect 6420 30676 6426 30688
rect 6457 30685 6469 30688
rect 6503 30685 6515 30719
rect 6457 30679 6515 30685
rect 7101 30719 7159 30725
rect 7101 30685 7113 30719
rect 7147 30685 7159 30719
rect 7101 30679 7159 30685
rect 7650 30676 7656 30728
rect 7708 30716 7714 30728
rect 8297 30719 8355 30725
rect 8297 30716 8309 30719
rect 7708 30688 8309 30716
rect 7708 30676 7714 30688
rect 8297 30685 8309 30688
rect 8343 30685 8355 30719
rect 8297 30679 8355 30685
rect 9677 30719 9735 30725
rect 9677 30685 9689 30719
rect 9723 30716 9735 30719
rect 12434 30716 12440 30728
rect 9723 30688 12440 30716
rect 9723 30685 9735 30688
rect 9677 30679 9735 30685
rect 12434 30676 12440 30688
rect 12492 30676 12498 30728
rect 12894 30716 12900 30728
rect 12855 30688 12900 30716
rect 12894 30676 12900 30688
rect 12952 30676 12958 30728
rect 26142 30716 26148 30728
rect 26103 30688 26148 30716
rect 26142 30676 26148 30688
rect 26200 30676 26206 30728
rect 27985 30719 28043 30725
rect 27985 30685 27997 30719
rect 28031 30716 28043 30719
rect 31726 30716 31754 30824
rect 37274 30812 37280 30824
rect 37332 30812 37338 30864
rect 37737 30787 37795 30793
rect 37737 30784 37749 30787
rect 28031 30688 31754 30716
rect 35866 30756 37749 30784
rect 28031 30685 28043 30688
rect 27985 30679 28043 30685
rect 7193 30651 7251 30657
rect 7193 30617 7205 30651
rect 7239 30648 7251 30651
rect 9858 30648 9864 30660
rect 7239 30620 9864 30648
rect 7239 30617 7251 30620
rect 7193 30611 7251 30617
rect 9858 30608 9864 30620
rect 9916 30608 9922 30660
rect 26160 30648 26188 30676
rect 35866 30648 35894 30756
rect 37737 30753 37749 30756
rect 37783 30753 37795 30787
rect 37737 30747 37795 30753
rect 37458 30716 37464 30728
rect 37419 30688 37464 30716
rect 37458 30676 37464 30688
rect 37516 30676 37522 30728
rect 26160 30620 35894 30648
rect 4065 30583 4123 30589
rect 4065 30549 4077 30583
rect 4111 30580 4123 30583
rect 5350 30580 5356 30592
rect 4111 30552 5356 30580
rect 4111 30549 4123 30552
rect 4065 30543 4123 30549
rect 5350 30540 5356 30552
rect 5408 30540 5414 30592
rect 6546 30580 6552 30592
rect 6507 30552 6552 30580
rect 6546 30540 6552 30552
rect 6604 30540 6610 30592
rect 9769 30583 9827 30589
rect 9769 30549 9781 30583
rect 9815 30580 9827 30583
rect 10318 30580 10324 30592
rect 9815 30552 10324 30580
rect 9815 30549 9827 30552
rect 9769 30543 9827 30549
rect 10318 30540 10324 30552
rect 10376 30540 10382 30592
rect 12989 30583 13047 30589
rect 12989 30549 13001 30583
rect 13035 30580 13047 30583
rect 13354 30580 13360 30592
rect 13035 30552 13360 30580
rect 13035 30549 13047 30552
rect 12989 30543 13047 30549
rect 13354 30540 13360 30552
rect 13412 30540 13418 30592
rect 28074 30580 28080 30592
rect 28035 30552 28080 30580
rect 28074 30540 28080 30552
rect 28132 30540 28138 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 13262 30336 13268 30388
rect 13320 30376 13326 30388
rect 14090 30376 14096 30388
rect 13320 30348 14096 30376
rect 13320 30336 13326 30348
rect 14090 30336 14096 30348
rect 14148 30336 14154 30388
rect 1581 30243 1639 30249
rect 1581 30209 1593 30243
rect 1627 30209 1639 30243
rect 1581 30203 1639 30209
rect 1596 30172 1624 30203
rect 2682 30200 2688 30252
rect 2740 30240 2746 30252
rect 4341 30243 4399 30249
rect 4341 30240 4353 30243
rect 2740 30212 4353 30240
rect 2740 30200 2746 30212
rect 4341 30209 4353 30212
rect 4387 30209 4399 30243
rect 4341 30203 4399 30209
rect 5166 30172 5172 30184
rect 1596 30144 5172 30172
rect 5166 30132 5172 30144
rect 5224 30132 5230 30184
rect 1762 30036 1768 30048
rect 1723 30008 1768 30036
rect 1762 29996 1768 30008
rect 1820 29996 1826 30048
rect 4433 30039 4491 30045
rect 4433 30005 4445 30039
rect 4479 30036 4491 30039
rect 4982 30036 4988 30048
rect 4479 30008 4988 30036
rect 4479 30005 4491 30008
rect 4433 29999 4491 30005
rect 4982 29996 4988 30008
rect 5040 29996 5046 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 4062 29792 4068 29844
rect 4120 29832 4126 29844
rect 4893 29835 4951 29841
rect 4893 29832 4905 29835
rect 4120 29804 4905 29832
rect 4120 29792 4126 29804
rect 4893 29801 4905 29804
rect 4939 29801 4951 29835
rect 4893 29795 4951 29801
rect 27433 29835 27491 29841
rect 27433 29801 27445 29835
rect 27479 29832 27491 29835
rect 30466 29832 30472 29844
rect 27479 29804 30472 29832
rect 27479 29801 27491 29804
rect 27433 29795 27491 29801
rect 30466 29792 30472 29804
rect 30524 29792 30530 29844
rect 16758 29656 16764 29708
rect 16816 29696 16822 29708
rect 32398 29696 32404 29708
rect 16816 29668 32404 29696
rect 16816 29656 16822 29668
rect 32398 29656 32404 29668
rect 32456 29656 32462 29708
rect 1762 29628 1768 29640
rect 1723 29600 1768 29628
rect 1762 29588 1768 29600
rect 1820 29588 1826 29640
rect 5077 29631 5135 29637
rect 5077 29597 5089 29631
rect 5123 29628 5135 29631
rect 5810 29628 5816 29640
rect 5123 29600 5816 29628
rect 5123 29597 5135 29600
rect 5077 29591 5135 29597
rect 5810 29588 5816 29600
rect 5868 29588 5874 29640
rect 6822 29588 6828 29640
rect 6880 29628 6886 29640
rect 9125 29631 9183 29637
rect 9125 29628 9137 29631
rect 6880 29600 9137 29628
rect 6880 29588 6886 29600
rect 9125 29597 9137 29600
rect 9171 29597 9183 29631
rect 9125 29591 9183 29597
rect 11793 29631 11851 29637
rect 11793 29597 11805 29631
rect 11839 29628 11851 29631
rect 16206 29628 16212 29640
rect 11839 29600 16212 29628
rect 11839 29597 11851 29600
rect 11793 29591 11851 29597
rect 16206 29588 16212 29600
rect 16264 29628 16270 29640
rect 17865 29631 17923 29637
rect 17865 29628 17877 29631
rect 16264 29600 17877 29628
rect 16264 29588 16270 29600
rect 17865 29597 17877 29600
rect 17911 29597 17923 29631
rect 17865 29591 17923 29597
rect 17954 29588 17960 29640
rect 18012 29628 18018 29640
rect 27341 29631 27399 29637
rect 27341 29628 27353 29631
rect 18012 29600 27353 29628
rect 18012 29588 18018 29600
rect 27341 29597 27353 29600
rect 27387 29597 27399 29631
rect 27341 29591 27399 29597
rect 37366 29588 37372 29640
rect 37424 29628 37430 29640
rect 38013 29631 38071 29637
rect 38013 29628 38025 29631
rect 37424 29600 38025 29628
rect 37424 29588 37430 29600
rect 38013 29597 38025 29600
rect 38059 29597 38071 29631
rect 38013 29591 38071 29597
rect 9217 29563 9275 29569
rect 9217 29529 9229 29563
rect 9263 29560 9275 29563
rect 14274 29560 14280 29572
rect 9263 29532 14280 29560
rect 9263 29529 9275 29532
rect 9217 29523 9275 29529
rect 14274 29520 14280 29532
rect 14332 29520 14338 29572
rect 1581 29495 1639 29501
rect 1581 29461 1593 29495
rect 1627 29492 1639 29495
rect 4706 29492 4712 29504
rect 1627 29464 4712 29492
rect 1627 29461 1639 29464
rect 1581 29455 1639 29461
rect 4706 29452 4712 29464
rect 4764 29452 4770 29504
rect 11609 29495 11667 29501
rect 11609 29461 11621 29495
rect 11655 29492 11667 29495
rect 11882 29492 11888 29504
rect 11655 29464 11888 29492
rect 11655 29461 11667 29464
rect 11609 29455 11667 29461
rect 11882 29452 11888 29464
rect 11940 29452 11946 29504
rect 17678 29492 17684 29504
rect 17639 29464 17684 29492
rect 17678 29452 17684 29464
rect 17736 29452 17742 29504
rect 38194 29492 38200 29504
rect 38155 29464 38200 29492
rect 38194 29452 38200 29464
rect 38252 29452 38258 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 5718 29248 5724 29300
rect 5776 29288 5782 29300
rect 8205 29291 8263 29297
rect 8205 29288 8217 29291
rect 5776 29260 8217 29288
rect 5776 29248 5782 29260
rect 8205 29257 8217 29260
rect 8251 29257 8263 29291
rect 16850 29288 16856 29300
rect 16811 29260 16856 29288
rect 8205 29251 8263 29257
rect 16850 29248 16856 29260
rect 16908 29248 16914 29300
rect 1765 29155 1823 29161
rect 1765 29121 1777 29155
rect 1811 29152 1823 29155
rect 2774 29152 2780 29164
rect 1811 29124 2780 29152
rect 1811 29121 1823 29124
rect 1765 29115 1823 29121
rect 2774 29112 2780 29124
rect 2832 29112 2838 29164
rect 8113 29155 8171 29161
rect 8113 29121 8125 29155
rect 8159 29152 8171 29155
rect 8294 29152 8300 29164
rect 8159 29124 8300 29152
rect 8159 29121 8171 29124
rect 8113 29115 8171 29121
rect 8294 29112 8300 29124
rect 8352 29112 8358 29164
rect 11882 29152 11888 29164
rect 11843 29124 11888 29152
rect 11882 29112 11888 29124
rect 11940 29112 11946 29164
rect 16666 29112 16672 29164
rect 16724 29152 16730 29164
rect 17037 29155 17095 29161
rect 17037 29152 17049 29155
rect 16724 29124 17049 29152
rect 16724 29112 16730 29124
rect 17037 29121 17049 29124
rect 17083 29121 17095 29155
rect 17678 29152 17684 29164
rect 17639 29124 17684 29152
rect 17037 29115 17095 29121
rect 17678 29112 17684 29124
rect 17736 29112 17742 29164
rect 1578 29016 1584 29028
rect 1539 28988 1584 29016
rect 1578 28976 1584 28988
rect 1636 28976 1642 29028
rect 10594 28976 10600 29028
rect 10652 29016 10658 29028
rect 11701 29019 11759 29025
rect 11701 29016 11713 29019
rect 10652 28988 11713 29016
rect 10652 28976 10658 28988
rect 11701 28985 11713 28988
rect 11747 28985 11759 29019
rect 11701 28979 11759 28985
rect 17494 28948 17500 28960
rect 17455 28920 17500 28948
rect 17494 28908 17500 28920
rect 17552 28908 17558 28960
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 16850 28636 16856 28688
rect 16908 28676 16914 28688
rect 17221 28679 17279 28685
rect 17221 28676 17233 28679
rect 16908 28648 17233 28676
rect 16908 28636 16914 28648
rect 17221 28645 17233 28648
rect 17267 28645 17279 28679
rect 17221 28639 17279 28645
rect 750 28568 756 28620
rect 808 28608 814 28620
rect 17037 28611 17095 28617
rect 808 28580 2544 28608
rect 808 28568 814 28580
rect 1854 28540 1860 28552
rect 1815 28512 1860 28540
rect 1854 28500 1860 28512
rect 1912 28500 1918 28552
rect 2516 28549 2544 28580
rect 17037 28577 17049 28611
rect 17083 28608 17095 28611
rect 17494 28608 17500 28620
rect 17083 28580 17500 28608
rect 17083 28577 17095 28580
rect 17037 28571 17095 28577
rect 17494 28568 17500 28580
rect 17552 28568 17558 28620
rect 2501 28543 2559 28549
rect 2501 28509 2513 28543
rect 2547 28509 2559 28543
rect 2501 28503 2559 28509
rect 15746 28500 15752 28552
rect 15804 28540 15810 28552
rect 16206 28540 16212 28552
rect 15804 28512 16212 28540
rect 15804 28500 15810 28512
rect 16206 28500 16212 28512
rect 16264 28500 16270 28552
rect 16853 28543 16911 28549
rect 16853 28509 16865 28543
rect 16899 28540 16911 28543
rect 16942 28540 16948 28552
rect 16899 28512 16948 28540
rect 16899 28509 16911 28512
rect 16853 28503 16911 28509
rect 16942 28500 16948 28512
rect 17000 28500 17006 28552
rect 1949 28475 2007 28481
rect 1949 28441 1961 28475
rect 1995 28472 2007 28475
rect 2866 28472 2872 28484
rect 1995 28444 2872 28472
rect 1995 28441 2007 28444
rect 1949 28435 2007 28441
rect 2866 28432 2872 28444
rect 2924 28432 2930 28484
rect 2314 28364 2320 28416
rect 2372 28404 2378 28416
rect 2593 28407 2651 28413
rect 2593 28404 2605 28407
rect 2372 28376 2605 28404
rect 2372 28364 2378 28376
rect 2593 28373 2605 28376
rect 2639 28373 2651 28407
rect 2593 28367 2651 28373
rect 16301 28407 16359 28413
rect 16301 28373 16313 28407
rect 16347 28404 16359 28407
rect 17494 28404 17500 28416
rect 16347 28376 17500 28404
rect 16347 28373 16359 28376
rect 16301 28367 16359 28373
rect 17494 28364 17500 28376
rect 17552 28364 17558 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 5810 28200 5816 28212
rect 5771 28172 5816 28200
rect 5810 28160 5816 28172
rect 5868 28160 5874 28212
rect 16942 28200 16948 28212
rect 16903 28172 16948 28200
rect 16942 28160 16948 28172
rect 17000 28160 17006 28212
rect 21358 28200 21364 28212
rect 21319 28172 21364 28200
rect 21358 28160 21364 28172
rect 21416 28160 21422 28212
rect 1946 28064 1952 28076
rect 1907 28036 1952 28064
rect 1946 28024 1952 28036
rect 2004 28024 2010 28076
rect 2590 28064 2596 28076
rect 2551 28036 2596 28064
rect 2590 28024 2596 28036
rect 2648 28024 2654 28076
rect 3418 28064 3424 28076
rect 3379 28036 3424 28064
rect 3418 28024 3424 28036
rect 3476 28024 3482 28076
rect 4062 28064 4068 28076
rect 4023 28036 4068 28064
rect 4062 28024 4068 28036
rect 4120 28024 4126 28076
rect 5721 28067 5779 28073
rect 5721 28033 5733 28067
rect 5767 28064 5779 28067
rect 6454 28064 6460 28076
rect 5767 28036 6460 28064
rect 5767 28033 5779 28036
rect 5721 28027 5779 28033
rect 6454 28024 6460 28036
rect 6512 28024 6518 28076
rect 8297 28067 8355 28073
rect 8297 28033 8309 28067
rect 8343 28064 8355 28067
rect 8386 28064 8392 28076
rect 8343 28036 8392 28064
rect 8343 28033 8355 28036
rect 8297 28027 8355 28033
rect 8386 28024 8392 28036
rect 8444 28024 8450 28076
rect 8941 28067 8999 28073
rect 8941 28033 8953 28067
rect 8987 28033 8999 28067
rect 12618 28064 12624 28076
rect 12579 28036 12624 28064
rect 8941 28027 8999 28033
rect 8956 27996 8984 28027
rect 12618 28024 12624 28036
rect 12676 28024 12682 28076
rect 17678 28064 17684 28076
rect 17639 28036 17684 28064
rect 17678 28024 17684 28036
rect 17736 28024 17742 28076
rect 19242 28064 19248 28076
rect 19203 28036 19248 28064
rect 19242 28024 19248 28036
rect 19300 28024 19306 28076
rect 21269 28067 21327 28073
rect 21269 28033 21281 28067
rect 21315 28033 21327 28067
rect 21269 28027 21327 28033
rect 8128 27968 8984 27996
rect 1578 27888 1584 27940
rect 1636 27928 1642 27940
rect 8128 27937 8156 27968
rect 9674 27956 9680 28008
rect 9732 27996 9738 28008
rect 10413 27999 10471 28005
rect 10413 27996 10425 27999
rect 9732 27968 10425 27996
rect 9732 27956 9738 27968
rect 10413 27965 10425 27968
rect 10459 27965 10471 27999
rect 10413 27959 10471 27965
rect 10597 27999 10655 28005
rect 10597 27965 10609 27999
rect 10643 27996 10655 27999
rect 12713 27999 12771 28005
rect 12713 27996 12725 27999
rect 10643 27968 12725 27996
rect 10643 27965 10655 27968
rect 10597 27959 10655 27965
rect 12713 27965 12725 27968
rect 12759 27965 12771 27999
rect 12713 27959 12771 27965
rect 16942 27956 16948 28008
rect 17000 27996 17006 28008
rect 21284 27996 21312 28027
rect 37458 27996 37464 28008
rect 17000 27968 21312 27996
rect 37419 27968 37464 27996
rect 17000 27956 17006 27968
rect 37458 27956 37464 27968
rect 37516 27956 37522 28008
rect 37737 27999 37795 28005
rect 37737 27965 37749 27999
rect 37783 27996 37795 27999
rect 37826 27996 37832 28008
rect 37783 27968 37832 27996
rect 37783 27965 37795 27968
rect 37737 27959 37795 27965
rect 37826 27956 37832 27968
rect 37884 27956 37890 28008
rect 2685 27931 2743 27937
rect 2685 27928 2697 27931
rect 1636 27900 2697 27928
rect 1636 27888 1642 27900
rect 2685 27897 2697 27900
rect 2731 27897 2743 27931
rect 2685 27891 2743 27897
rect 8113 27931 8171 27937
rect 8113 27897 8125 27931
rect 8159 27897 8171 27931
rect 8113 27891 8171 27897
rect 2038 27860 2044 27872
rect 1999 27832 2044 27860
rect 2038 27820 2044 27832
rect 2096 27820 2102 27872
rect 3234 27860 3240 27872
rect 3195 27832 3240 27860
rect 3234 27820 3240 27832
rect 3292 27820 3298 27872
rect 3881 27863 3939 27869
rect 3881 27829 3893 27863
rect 3927 27860 3939 27863
rect 5074 27860 5080 27872
rect 3927 27832 5080 27860
rect 3927 27829 3939 27832
rect 3881 27823 3939 27829
rect 5074 27820 5080 27832
rect 5132 27820 5138 27872
rect 8202 27820 8208 27872
rect 8260 27860 8266 27872
rect 8757 27863 8815 27869
rect 8757 27860 8769 27863
rect 8260 27832 8769 27860
rect 8260 27820 8266 27832
rect 8757 27829 8769 27832
rect 8803 27829 8815 27863
rect 8757 27823 8815 27829
rect 11057 27863 11115 27869
rect 11057 27829 11069 27863
rect 11103 27860 11115 27863
rect 11146 27860 11152 27872
rect 11103 27832 11152 27860
rect 11103 27829 11115 27832
rect 11057 27823 11115 27829
rect 11146 27820 11152 27832
rect 11204 27820 11210 27872
rect 17034 27820 17040 27872
rect 17092 27860 17098 27872
rect 17773 27863 17831 27869
rect 17773 27860 17785 27863
rect 17092 27832 17785 27860
rect 17092 27820 17098 27832
rect 17773 27829 17785 27832
rect 17819 27829 17831 27863
rect 17773 27823 17831 27829
rect 17862 27820 17868 27872
rect 17920 27860 17926 27872
rect 19061 27863 19119 27869
rect 19061 27860 19073 27863
rect 17920 27832 19073 27860
rect 17920 27820 17926 27832
rect 19061 27829 19073 27832
rect 19107 27829 19119 27863
rect 19061 27823 19119 27829
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 17678 27616 17684 27668
rect 17736 27656 17742 27668
rect 18693 27659 18751 27665
rect 17736 27628 18184 27656
rect 17736 27616 17742 27628
rect 11057 27591 11115 27597
rect 11057 27557 11069 27591
rect 11103 27588 11115 27591
rect 12066 27588 12072 27600
rect 11103 27560 12072 27588
rect 11103 27557 11115 27560
rect 11057 27551 11115 27557
rect 12066 27548 12072 27560
rect 12124 27588 12130 27600
rect 17313 27591 17371 27597
rect 17313 27588 17325 27591
rect 12124 27560 17325 27588
rect 12124 27548 12130 27560
rect 17313 27557 17325 27560
rect 17359 27557 17371 27591
rect 17313 27551 17371 27557
rect 6546 27480 6552 27532
rect 6604 27520 6610 27532
rect 10413 27523 10471 27529
rect 10413 27520 10425 27523
rect 6604 27492 10425 27520
rect 6604 27480 6610 27492
rect 10413 27489 10425 27492
rect 10459 27489 10471 27523
rect 10594 27520 10600 27532
rect 10555 27492 10600 27520
rect 10413 27483 10471 27489
rect 10594 27480 10600 27492
rect 10652 27480 10658 27532
rect 15746 27480 15752 27532
rect 15804 27520 15810 27532
rect 17129 27523 17187 27529
rect 15804 27492 17080 27520
rect 15804 27480 15810 27492
rect 1854 27452 1860 27464
rect 1815 27424 1860 27452
rect 1854 27412 1860 27424
rect 1912 27412 1918 27464
rect 2498 27452 2504 27464
rect 2459 27424 2504 27452
rect 2498 27412 2504 27424
rect 2556 27412 2562 27464
rect 3145 27455 3203 27461
rect 3145 27421 3157 27455
rect 3191 27421 3203 27455
rect 3145 27415 3203 27421
rect 3160 27384 3188 27415
rect 3234 27412 3240 27464
rect 3292 27452 3298 27464
rect 3973 27455 4031 27461
rect 3973 27452 3985 27455
rect 3292 27424 3985 27452
rect 3292 27412 3298 27424
rect 3973 27421 3985 27424
rect 4019 27421 4031 27455
rect 3973 27415 4031 27421
rect 7745 27455 7803 27461
rect 7745 27421 7757 27455
rect 7791 27452 7803 27455
rect 8386 27452 8392 27464
rect 7791 27424 8392 27452
rect 7791 27421 7803 27424
rect 7745 27415 7803 27421
rect 8386 27412 8392 27424
rect 8444 27452 8450 27464
rect 8938 27452 8944 27464
rect 8444 27424 8944 27452
rect 8444 27412 8450 27424
rect 8938 27412 8944 27424
rect 8996 27412 9002 27464
rect 9953 27455 10011 27461
rect 9953 27421 9965 27455
rect 9999 27421 10011 27455
rect 9953 27415 10011 27421
rect 12989 27455 13047 27461
rect 12989 27421 13001 27455
rect 13035 27452 13047 27455
rect 13170 27452 13176 27464
rect 13035 27424 13176 27452
rect 13035 27421 13047 27424
rect 12989 27415 13047 27421
rect 3878 27384 3884 27396
rect 3160 27356 3884 27384
rect 3878 27344 3884 27356
rect 3936 27344 3942 27396
rect 9968 27384 9996 27415
rect 13170 27412 13176 27424
rect 13228 27412 13234 27464
rect 16945 27455 17003 27461
rect 16945 27421 16957 27455
rect 16991 27421 17003 27455
rect 17052 27452 17080 27492
rect 17129 27489 17141 27523
rect 17175 27520 17187 27523
rect 17494 27520 17500 27532
rect 17175 27492 17500 27520
rect 17175 27489 17187 27492
rect 17129 27483 17187 27489
rect 17494 27480 17500 27492
rect 17552 27480 17558 27532
rect 18049 27455 18107 27461
rect 18049 27452 18061 27455
rect 17052 27424 18061 27452
rect 16945 27415 17003 27421
rect 18049 27421 18061 27424
rect 18095 27421 18107 27455
rect 18156 27452 18184 27628
rect 18693 27625 18705 27659
rect 18739 27656 18751 27659
rect 19242 27656 19248 27668
rect 18739 27628 19248 27656
rect 18739 27625 18751 27628
rect 18693 27619 18751 27625
rect 19242 27616 19248 27628
rect 19300 27616 19306 27668
rect 37366 27588 37372 27600
rect 37327 27560 37372 27588
rect 37366 27548 37372 27560
rect 37424 27548 37430 27600
rect 18877 27455 18935 27461
rect 18877 27452 18889 27455
rect 18156 27424 18889 27452
rect 18049 27415 18107 27421
rect 18877 27421 18889 27424
rect 18923 27421 18935 27455
rect 18877 27415 18935 27421
rect 16960 27384 16988 27415
rect 19334 27412 19340 27464
rect 19392 27452 19398 27464
rect 19429 27455 19487 27461
rect 19429 27452 19441 27455
rect 19392 27424 19441 27452
rect 19392 27412 19398 27424
rect 19429 27421 19441 27424
rect 19475 27421 19487 27455
rect 19429 27415 19487 27421
rect 22094 27412 22100 27464
rect 22152 27452 22158 27464
rect 37550 27452 37556 27464
rect 22152 27424 22197 27452
rect 37511 27424 37556 27452
rect 22152 27412 22158 27424
rect 37550 27412 37556 27424
rect 37608 27412 37614 27464
rect 38010 27452 38016 27464
rect 37971 27424 38016 27452
rect 38010 27412 38016 27424
rect 38068 27412 38074 27464
rect 20346 27384 20352 27396
rect 9968 27356 12020 27384
rect 16960 27356 20352 27384
rect 11992 27328 12020 27356
rect 20346 27344 20352 27356
rect 20404 27344 20410 27396
rect 1946 27316 1952 27328
rect 1907 27288 1952 27316
rect 1946 27276 1952 27288
rect 2004 27276 2010 27328
rect 2130 27276 2136 27328
rect 2188 27316 2194 27328
rect 2593 27319 2651 27325
rect 2593 27316 2605 27319
rect 2188 27288 2605 27316
rect 2188 27276 2194 27288
rect 2593 27285 2605 27288
rect 2639 27285 2651 27319
rect 2593 27279 2651 27285
rect 3237 27319 3295 27325
rect 3237 27285 3249 27319
rect 3283 27316 3295 27319
rect 3694 27316 3700 27328
rect 3283 27288 3700 27316
rect 3283 27285 3295 27288
rect 3237 27279 3295 27285
rect 3694 27276 3700 27288
rect 3752 27276 3758 27328
rect 7834 27316 7840 27328
rect 7795 27288 7840 27316
rect 7834 27276 7840 27288
rect 7892 27276 7898 27328
rect 9769 27319 9827 27325
rect 9769 27285 9781 27319
rect 9815 27316 9827 27319
rect 10042 27316 10048 27328
rect 9815 27288 10048 27316
rect 9815 27285 9827 27288
rect 9769 27279 9827 27285
rect 10042 27276 10048 27288
rect 10100 27276 10106 27328
rect 11974 27276 11980 27328
rect 12032 27316 12038 27328
rect 12618 27316 12624 27328
rect 12032 27288 12624 27316
rect 12032 27276 12038 27288
rect 12618 27276 12624 27288
rect 12676 27276 12682 27328
rect 12710 27276 12716 27328
rect 12768 27316 12774 27328
rect 12805 27319 12863 27325
rect 12805 27316 12817 27319
rect 12768 27288 12817 27316
rect 12768 27276 12774 27288
rect 12805 27285 12817 27288
rect 12851 27285 12863 27319
rect 18138 27316 18144 27328
rect 18099 27288 18144 27316
rect 12805 27279 12863 27285
rect 18138 27276 18144 27288
rect 18196 27276 18202 27328
rect 18782 27276 18788 27328
rect 18840 27316 18846 27328
rect 19521 27319 19579 27325
rect 19521 27316 19533 27319
rect 18840 27288 19533 27316
rect 18840 27276 18846 27288
rect 19521 27285 19533 27288
rect 19567 27285 19579 27319
rect 19521 27279 19579 27285
rect 22189 27319 22247 27325
rect 22189 27285 22201 27319
rect 22235 27316 22247 27319
rect 22554 27316 22560 27328
rect 22235 27288 22560 27316
rect 22235 27285 22247 27288
rect 22189 27279 22247 27285
rect 22554 27276 22560 27288
rect 22612 27276 22618 27328
rect 38194 27316 38200 27328
rect 38155 27288 38200 27316
rect 38194 27276 38200 27288
rect 38252 27276 38258 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 2958 27072 2964 27124
rect 3016 27112 3022 27124
rect 5166 27112 5172 27124
rect 3016 27084 4568 27112
rect 5127 27084 5172 27112
rect 3016 27072 3022 27084
rect 1210 27004 1216 27056
rect 1268 27044 1274 27056
rect 4540 27044 4568 27084
rect 5166 27072 5172 27084
rect 5224 27072 5230 27124
rect 11146 27072 11152 27124
rect 11204 27112 11210 27124
rect 11204 27084 14688 27112
rect 11204 27072 11210 27084
rect 12710 27044 12716 27056
rect 1268 27016 4476 27044
rect 4540 27016 7144 27044
rect 12671 27016 12716 27044
rect 1268 27004 1274 27016
rect 566 26936 572 26988
rect 624 26976 630 26988
rect 1854 26976 1860 26988
rect 624 26948 1860 26976
rect 624 26936 630 26948
rect 1854 26936 1860 26948
rect 1912 26976 1918 26988
rect 2501 26979 2559 26985
rect 2501 26976 2513 26979
rect 1912 26948 2513 26976
rect 1912 26936 1918 26948
rect 2501 26945 2513 26948
rect 2547 26976 2559 26979
rect 2958 26976 2964 26988
rect 2547 26948 2964 26976
rect 2547 26945 2559 26948
rect 2501 26939 2559 26945
rect 2958 26936 2964 26948
rect 3016 26936 3022 26988
rect 4448 26985 4476 27016
rect 3789 26979 3847 26985
rect 3789 26945 3801 26979
rect 3835 26945 3847 26979
rect 3789 26939 3847 26945
rect 4433 26979 4491 26985
rect 4433 26945 4445 26979
rect 4479 26945 4491 26979
rect 4433 26939 4491 26945
rect 5353 26979 5411 26985
rect 5353 26945 5365 26979
rect 5399 26976 5411 26979
rect 6822 26976 6828 26988
rect 5399 26948 6828 26976
rect 5399 26945 5411 26948
rect 5353 26939 5411 26945
rect 3050 26868 3056 26920
rect 3108 26908 3114 26920
rect 3145 26911 3203 26917
rect 3145 26908 3157 26911
rect 3108 26880 3157 26908
rect 3108 26868 3114 26880
rect 3145 26877 3157 26880
rect 3191 26877 3203 26911
rect 3804 26908 3832 26939
rect 6822 26936 6828 26948
rect 6880 26936 6886 26988
rect 7116 26985 7144 27016
rect 12710 27004 12716 27016
rect 12768 27004 12774 27056
rect 7101 26979 7159 26985
rect 7101 26945 7113 26979
rect 7147 26945 7159 26979
rect 7101 26939 7159 26945
rect 11238 26936 11244 26988
rect 11296 26976 11302 26988
rect 11885 26979 11943 26985
rect 11885 26976 11897 26979
rect 11296 26948 11897 26976
rect 11296 26936 11302 26948
rect 11885 26945 11897 26948
rect 11931 26945 11943 26979
rect 11885 26939 11943 26945
rect 5258 26908 5264 26920
rect 3804 26880 5264 26908
rect 3145 26871 3203 26877
rect 5258 26868 5264 26880
rect 5316 26868 5322 26920
rect 12621 26911 12679 26917
rect 12621 26877 12633 26911
rect 12667 26877 12679 26911
rect 12621 26871 12679 26877
rect 842 26800 848 26852
rect 900 26840 906 26852
rect 2593 26843 2651 26849
rect 2593 26840 2605 26843
rect 900 26812 2605 26840
rect 900 26800 906 26812
rect 2593 26809 2605 26812
rect 2639 26809 2651 26843
rect 2593 26803 2651 26809
rect 1118 26732 1124 26784
rect 1176 26772 1182 26784
rect 1949 26775 2007 26781
rect 1949 26772 1961 26775
rect 1176 26744 1961 26772
rect 1176 26732 1182 26744
rect 1949 26741 1961 26744
rect 1995 26741 2007 26775
rect 1949 26735 2007 26741
rect 3142 26732 3148 26784
rect 3200 26772 3206 26784
rect 3881 26775 3939 26781
rect 3881 26772 3893 26775
rect 3200 26744 3893 26772
rect 3200 26732 3206 26744
rect 3881 26741 3893 26744
rect 3927 26741 3939 26775
rect 3881 26735 3939 26741
rect 4525 26775 4583 26781
rect 4525 26741 4537 26775
rect 4571 26772 4583 26775
rect 4614 26772 4620 26784
rect 4571 26744 4620 26772
rect 4571 26741 4583 26744
rect 4525 26735 4583 26741
rect 4614 26732 4620 26744
rect 4672 26732 4678 26784
rect 7193 26775 7251 26781
rect 7193 26741 7205 26775
rect 7239 26772 7251 26775
rect 7282 26772 7288 26784
rect 7239 26744 7288 26772
rect 7239 26741 7251 26744
rect 7193 26735 7251 26741
rect 7282 26732 7288 26744
rect 7340 26732 7346 26784
rect 11977 26775 12035 26781
rect 11977 26741 11989 26775
rect 12023 26772 12035 26775
rect 12158 26772 12164 26784
rect 12023 26744 12164 26772
rect 12023 26741 12035 26744
rect 11977 26735 12035 26741
rect 12158 26732 12164 26744
rect 12216 26732 12222 26784
rect 12636 26772 12664 26871
rect 12710 26868 12716 26920
rect 12768 26908 12774 26920
rect 12897 26911 12955 26917
rect 12897 26908 12909 26911
rect 12768 26880 12909 26908
rect 12768 26868 12774 26880
rect 12897 26877 12909 26880
rect 12943 26877 12955 26911
rect 14660 26908 14688 27084
rect 17494 27072 17500 27124
rect 17552 27112 17558 27124
rect 28074 27112 28080 27124
rect 17552 27084 28080 27112
rect 17552 27072 17558 27084
rect 28074 27072 28080 27084
rect 28132 27072 28138 27124
rect 37550 27112 37556 27124
rect 37511 27084 37556 27112
rect 37550 27072 37556 27084
rect 37608 27072 37614 27124
rect 17034 27044 17040 27056
rect 16995 27016 17040 27044
rect 17034 27004 17040 27016
rect 17092 27004 17098 27056
rect 17589 27047 17647 27053
rect 17589 27013 17601 27047
rect 17635 27044 17647 27047
rect 17954 27044 17960 27056
rect 17635 27016 17960 27044
rect 17635 27013 17647 27016
rect 17589 27007 17647 27013
rect 17954 27004 17960 27016
rect 18012 27004 18018 27056
rect 18785 26979 18843 26985
rect 18785 26945 18797 26979
rect 18831 26976 18843 26979
rect 22094 26976 22100 26988
rect 18831 26948 22100 26976
rect 18831 26945 18843 26948
rect 18785 26939 18843 26945
rect 22094 26936 22100 26948
rect 22152 26936 22158 26988
rect 37274 26936 37280 26988
rect 37332 26976 37338 26988
rect 37461 26979 37519 26985
rect 37461 26976 37473 26979
rect 37332 26948 37473 26976
rect 37332 26936 37338 26948
rect 37461 26945 37473 26948
rect 37507 26945 37519 26979
rect 37461 26939 37519 26945
rect 16945 26911 17003 26917
rect 16945 26908 16957 26911
rect 14660 26880 16957 26908
rect 12897 26871 12955 26877
rect 16945 26877 16957 26880
rect 16991 26877 17003 26911
rect 16945 26871 17003 26877
rect 18138 26868 18144 26920
rect 18196 26908 18202 26920
rect 18969 26911 19027 26917
rect 18969 26908 18981 26911
rect 18196 26880 18981 26908
rect 18196 26868 18202 26880
rect 18969 26877 18981 26880
rect 19015 26877 19027 26911
rect 18969 26871 19027 26877
rect 22462 26868 22468 26920
rect 22520 26908 22526 26920
rect 28350 26908 28356 26920
rect 22520 26880 28356 26908
rect 22520 26868 22526 26880
rect 28350 26868 28356 26880
rect 28408 26868 28414 26920
rect 16850 26772 16856 26784
rect 12636 26744 16856 26772
rect 16850 26732 16856 26744
rect 16908 26772 16914 26784
rect 19337 26775 19395 26781
rect 19337 26772 19349 26775
rect 16908 26744 19349 26772
rect 16908 26732 16914 26744
rect 19337 26741 19349 26744
rect 19383 26741 19395 26775
rect 19337 26735 19395 26741
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 8294 26568 8300 26580
rect 8255 26540 8300 26568
rect 8294 26528 8300 26540
rect 8352 26528 8358 26580
rect 11238 26528 11244 26580
rect 11296 26568 11302 26580
rect 12986 26568 12992 26580
rect 11296 26540 12992 26568
rect 11296 26528 11302 26540
rect 12986 26528 12992 26540
rect 13044 26528 13050 26580
rect 13170 26568 13176 26580
rect 13131 26540 13176 26568
rect 13170 26528 13176 26540
rect 13228 26528 13234 26580
rect 14826 26528 14832 26580
rect 14884 26568 14890 26580
rect 15838 26568 15844 26580
rect 14884 26540 15844 26568
rect 14884 26528 14890 26540
rect 15838 26528 15844 26540
rect 15896 26568 15902 26580
rect 15896 26540 20944 26568
rect 15896 26528 15902 26540
rect 5813 26503 5871 26509
rect 5813 26469 5825 26503
rect 5859 26469 5871 26503
rect 5813 26463 5871 26469
rect 7009 26503 7067 26509
rect 7009 26469 7021 26503
rect 7055 26500 7067 26503
rect 9582 26500 9588 26512
rect 7055 26472 9588 26500
rect 7055 26469 7067 26472
rect 7009 26463 7067 26469
rect 658 26392 664 26444
rect 716 26432 722 26444
rect 3237 26435 3295 26441
rect 3237 26432 3249 26435
rect 716 26404 3249 26432
rect 716 26392 722 26404
rect 3237 26401 3249 26404
rect 3283 26401 3295 26435
rect 5828 26432 5856 26463
rect 9582 26460 9588 26472
rect 9640 26460 9646 26512
rect 12250 26460 12256 26512
rect 12308 26500 12314 26512
rect 14461 26503 14519 26509
rect 14461 26500 14473 26503
rect 12308 26472 14473 26500
rect 12308 26460 12314 26472
rect 14461 26469 14473 26472
rect 14507 26469 14519 26503
rect 14461 26463 14519 26469
rect 15933 26503 15991 26509
rect 15933 26469 15945 26503
rect 15979 26469 15991 26503
rect 15933 26463 15991 26469
rect 7834 26432 7840 26444
rect 3237 26395 3295 26401
rect 4080 26404 5856 26432
rect 7795 26404 7840 26432
rect 1854 26364 1860 26376
rect 1815 26336 1860 26364
rect 1854 26324 1860 26336
rect 1912 26324 1918 26376
rect 2498 26364 2504 26376
rect 2459 26336 2504 26364
rect 2498 26324 2504 26336
rect 2556 26324 2562 26376
rect 2958 26324 2964 26376
rect 3016 26364 3022 26376
rect 4080 26373 4108 26404
rect 7834 26392 7840 26404
rect 7892 26392 7898 26444
rect 12066 26432 12072 26444
rect 12027 26404 12072 26432
rect 12066 26392 12072 26404
rect 12124 26392 12130 26444
rect 12434 26392 12440 26444
rect 12492 26432 12498 26444
rect 15948 26432 15976 26463
rect 20622 26432 20628 26444
rect 12492 26404 12537 26432
rect 15948 26404 16804 26432
rect 20583 26404 20628 26432
rect 12492 26392 12498 26404
rect 3145 26367 3203 26373
rect 3145 26364 3157 26367
rect 3016 26336 3157 26364
rect 3016 26324 3022 26336
rect 3145 26333 3157 26336
rect 3191 26333 3203 26367
rect 3145 26327 3203 26333
rect 4065 26367 4123 26373
rect 4065 26333 4077 26367
rect 4111 26333 4123 26367
rect 5166 26364 5172 26376
rect 5127 26336 5172 26364
rect 4065 26327 4123 26333
rect 5166 26324 5172 26336
rect 5224 26324 5230 26376
rect 5261 26367 5319 26373
rect 5261 26333 5273 26367
rect 5307 26364 5319 26367
rect 5442 26364 5448 26376
rect 5307 26336 5448 26364
rect 5307 26333 5319 26336
rect 5261 26327 5319 26333
rect 5442 26324 5448 26336
rect 5500 26324 5506 26376
rect 5997 26367 6055 26373
rect 5997 26333 6009 26367
rect 6043 26364 6055 26367
rect 6086 26364 6092 26376
rect 6043 26336 6092 26364
rect 6043 26333 6055 26336
rect 5997 26327 6055 26333
rect 6086 26324 6092 26336
rect 6144 26324 6150 26376
rect 6914 26364 6920 26376
rect 6875 26336 6920 26364
rect 6914 26324 6920 26336
rect 6972 26324 6978 26376
rect 7653 26367 7711 26373
rect 7653 26333 7665 26367
rect 7699 26364 7711 26367
rect 11054 26364 11060 26376
rect 7699 26336 11060 26364
rect 7699 26333 7711 26336
rect 7653 26327 7711 26333
rect 11054 26324 11060 26336
rect 11112 26324 11118 26376
rect 12986 26324 12992 26376
rect 13044 26364 13050 26376
rect 13357 26367 13415 26373
rect 13357 26364 13369 26367
rect 13044 26336 13369 26364
rect 13044 26324 13050 26336
rect 13357 26333 13369 26336
rect 13403 26333 13415 26367
rect 14366 26364 14372 26376
rect 14327 26336 14372 26364
rect 13357 26327 13415 26333
rect 14366 26324 14372 26336
rect 14424 26324 14430 26376
rect 16114 26364 16120 26376
rect 16075 26336 16120 26364
rect 16114 26324 16120 26336
rect 16172 26324 16178 26376
rect 16776 26373 16804 26404
rect 20622 26392 20628 26404
rect 20680 26392 20686 26444
rect 20916 26441 20944 26540
rect 34514 26460 34520 26512
rect 34572 26500 34578 26512
rect 38105 26503 38163 26509
rect 38105 26500 38117 26503
rect 34572 26472 38117 26500
rect 34572 26460 34578 26472
rect 38105 26469 38117 26472
rect 38151 26469 38163 26503
rect 38105 26463 38163 26469
rect 20901 26435 20959 26441
rect 20901 26401 20913 26435
rect 20947 26401 20959 26435
rect 20901 26395 20959 26401
rect 16761 26367 16819 26373
rect 16761 26333 16773 26367
rect 16807 26333 16819 26367
rect 38286 26364 38292 26376
rect 38247 26336 38292 26364
rect 16761 26327 16819 26333
rect 38286 26324 38292 26336
rect 38344 26324 38350 26376
rect 1946 26296 1952 26308
rect 1907 26268 1952 26296
rect 1946 26256 1952 26268
rect 2004 26256 2010 26308
rect 2593 26299 2651 26305
rect 2593 26265 2605 26299
rect 2639 26296 2651 26299
rect 2682 26296 2688 26308
rect 2639 26268 2688 26296
rect 2639 26265 2651 26268
rect 2593 26259 2651 26265
rect 2682 26256 2688 26268
rect 2740 26256 2746 26308
rect 4157 26299 4215 26305
rect 4157 26265 4169 26299
rect 4203 26296 4215 26299
rect 11422 26296 11428 26308
rect 4203 26268 11428 26296
rect 4203 26265 4215 26268
rect 4157 26259 4215 26265
rect 11422 26256 11428 26268
rect 11480 26256 11486 26308
rect 12158 26256 12164 26308
rect 12216 26296 12222 26308
rect 20717 26299 20775 26305
rect 12216 26268 12261 26296
rect 12216 26256 12222 26268
rect 20717 26265 20729 26299
rect 20763 26296 20775 26299
rect 20806 26296 20812 26308
rect 20763 26268 20812 26296
rect 20763 26265 20775 26268
rect 20717 26259 20775 26265
rect 20806 26256 20812 26268
rect 20864 26256 20870 26308
rect 16574 26228 16580 26240
rect 16535 26200 16580 26228
rect 16574 26188 16580 26200
rect 16632 26188 16638 26240
rect 17770 26228 17776 26240
rect 17731 26200 17776 26228
rect 17770 26188 17776 26200
rect 17828 26188 17834 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 6822 25984 6828 26036
rect 6880 26024 6886 26036
rect 7837 26027 7895 26033
rect 7837 26024 7849 26027
rect 6880 25996 7849 26024
rect 6880 25984 6886 25996
rect 7837 25993 7849 25996
rect 7883 25993 7895 26027
rect 7837 25987 7895 25993
rect 13357 26027 13415 26033
rect 13357 25993 13369 26027
rect 13403 25993 13415 26027
rect 13357 25987 13415 25993
rect 2038 25916 2044 25968
rect 2096 25956 2102 25968
rect 2682 25956 2688 25968
rect 2096 25928 2688 25956
rect 2096 25916 2102 25928
rect 2682 25916 2688 25928
rect 2740 25916 2746 25968
rect 5994 25956 6000 25968
rect 3252 25928 6000 25956
rect 1394 25848 1400 25900
rect 1452 25888 1458 25900
rect 3252 25897 3280 25928
rect 5994 25916 6000 25928
rect 6052 25916 6058 25968
rect 13372 25956 13400 25987
rect 17770 25956 17776 25968
rect 13372 25928 15516 25956
rect 17731 25928 17776 25956
rect 2133 25891 2191 25897
rect 2133 25888 2145 25891
rect 1452 25860 2145 25888
rect 1452 25848 1458 25860
rect 2133 25857 2145 25860
rect 2179 25857 2191 25891
rect 2133 25851 2191 25857
rect 3237 25891 3295 25897
rect 3237 25857 3249 25891
rect 3283 25857 3295 25891
rect 3237 25851 3295 25857
rect 3970 25848 3976 25900
rect 4028 25888 4034 25900
rect 4157 25891 4215 25897
rect 4157 25888 4169 25891
rect 4028 25860 4169 25888
rect 4028 25848 4034 25860
rect 4157 25857 4169 25860
rect 4203 25857 4215 25891
rect 4798 25888 4804 25900
rect 4759 25860 4804 25888
rect 4157 25851 4215 25857
rect 4798 25848 4804 25860
rect 4856 25848 4862 25900
rect 5626 25888 5632 25900
rect 5587 25860 5632 25888
rect 5626 25848 5632 25860
rect 5684 25848 5690 25900
rect 6549 25891 6607 25897
rect 6549 25857 6561 25891
rect 6595 25888 6607 25891
rect 6914 25888 6920 25900
rect 6595 25860 6920 25888
rect 6595 25857 6607 25860
rect 6549 25851 6607 25857
rect 6914 25848 6920 25860
rect 6972 25888 6978 25900
rect 7742 25888 7748 25900
rect 6972 25860 7144 25888
rect 7703 25860 7748 25888
rect 6972 25848 6978 25860
rect 5718 25780 5724 25832
rect 5776 25820 5782 25832
rect 6641 25823 6699 25829
rect 6641 25820 6653 25823
rect 5776 25792 6653 25820
rect 5776 25780 5782 25792
rect 6641 25789 6653 25792
rect 6687 25789 6699 25823
rect 7116 25820 7144 25860
rect 7742 25848 7748 25860
rect 7800 25848 7806 25900
rect 10686 25848 10692 25900
rect 10744 25888 10750 25900
rect 10965 25891 11023 25897
rect 10965 25888 10977 25891
rect 10744 25860 10977 25888
rect 10744 25848 10750 25860
rect 10965 25857 10977 25860
rect 11011 25857 11023 25891
rect 10965 25851 11023 25857
rect 13541 25891 13599 25897
rect 13541 25857 13553 25891
rect 13587 25888 13599 25891
rect 14001 25891 14059 25897
rect 14001 25888 14013 25891
rect 13587 25860 14013 25888
rect 13587 25857 13599 25860
rect 13541 25851 13599 25857
rect 14001 25857 14013 25860
rect 14047 25888 14059 25891
rect 14182 25888 14188 25900
rect 14047 25860 14188 25888
rect 14047 25857 14059 25860
rect 14001 25851 14059 25857
rect 14182 25848 14188 25860
rect 14240 25848 14246 25900
rect 14645 25891 14703 25897
rect 14645 25857 14657 25891
rect 14691 25888 14703 25891
rect 15010 25888 15016 25900
rect 14691 25860 15016 25888
rect 14691 25857 14703 25860
rect 14645 25851 14703 25857
rect 15010 25848 15016 25860
rect 15068 25848 15074 25900
rect 15488 25897 15516 25928
rect 17770 25916 17776 25928
rect 17828 25916 17834 25968
rect 17862 25916 17868 25968
rect 17920 25956 17926 25968
rect 17920 25928 17965 25956
rect 17920 25916 17926 25928
rect 15473 25891 15531 25897
rect 15473 25857 15485 25891
rect 15519 25857 15531 25891
rect 15473 25851 15531 25857
rect 7834 25820 7840 25832
rect 7116 25792 7840 25820
rect 6641 25783 6699 25789
rect 7834 25780 7840 25792
rect 7892 25780 7898 25832
rect 9674 25820 9680 25832
rect 9635 25792 9680 25820
rect 9674 25780 9680 25792
rect 9732 25780 9738 25832
rect 9861 25823 9919 25829
rect 9861 25789 9873 25823
rect 9907 25789 9919 25823
rect 9861 25783 9919 25789
rect 4893 25755 4951 25761
rect 4893 25721 4905 25755
rect 4939 25752 4951 25755
rect 7006 25752 7012 25764
rect 4939 25724 7012 25752
rect 4939 25721 4951 25724
rect 4893 25715 4951 25721
rect 7006 25712 7012 25724
rect 7064 25712 7070 25764
rect 9876 25752 9904 25783
rect 16298 25780 16304 25832
rect 16356 25820 16362 25832
rect 16853 25823 16911 25829
rect 16853 25820 16865 25823
rect 16356 25792 16865 25820
rect 16356 25780 16362 25792
rect 16853 25789 16865 25792
rect 16899 25789 16911 25823
rect 16853 25783 16911 25789
rect 17954 25780 17960 25832
rect 18012 25820 18018 25832
rect 18049 25823 18107 25829
rect 18049 25820 18061 25823
rect 18012 25792 18061 25820
rect 18012 25780 18018 25792
rect 18049 25789 18061 25792
rect 18095 25789 18107 25823
rect 18049 25783 18107 25789
rect 10781 25755 10839 25761
rect 10781 25752 10793 25755
rect 9876 25724 10793 25752
rect 10781 25721 10793 25724
rect 10827 25721 10839 25755
rect 10781 25715 10839 25721
rect 2225 25687 2283 25693
rect 2225 25653 2237 25687
rect 2271 25684 2283 25687
rect 2590 25684 2596 25696
rect 2271 25656 2596 25684
rect 2271 25653 2283 25656
rect 2225 25647 2283 25653
rect 2590 25644 2596 25656
rect 2648 25644 2654 25696
rect 3326 25684 3332 25696
rect 3287 25656 3332 25684
rect 3326 25644 3332 25656
rect 3384 25644 3390 25696
rect 3786 25644 3792 25696
rect 3844 25684 3850 25696
rect 4249 25687 4307 25693
rect 4249 25684 4261 25687
rect 3844 25656 4261 25684
rect 3844 25644 3850 25656
rect 4249 25653 4261 25656
rect 4295 25653 4307 25687
rect 4249 25647 4307 25653
rect 5721 25687 5779 25693
rect 5721 25653 5733 25687
rect 5767 25684 5779 25687
rect 6178 25684 6184 25696
rect 5767 25656 6184 25684
rect 5767 25653 5779 25656
rect 5721 25647 5779 25653
rect 6178 25644 6184 25656
rect 6236 25644 6242 25696
rect 6270 25644 6276 25696
rect 6328 25684 6334 25696
rect 10045 25687 10103 25693
rect 10045 25684 10057 25687
rect 6328 25656 10057 25684
rect 6328 25644 6334 25656
rect 10045 25653 10057 25656
rect 10091 25653 10103 25687
rect 14090 25684 14096 25696
rect 14051 25656 14096 25684
rect 10045 25647 10103 25653
rect 14090 25644 14096 25656
rect 14148 25644 14154 25696
rect 14734 25684 14740 25696
rect 14695 25656 14740 25684
rect 14734 25644 14740 25656
rect 14792 25644 14798 25696
rect 15286 25684 15292 25696
rect 15247 25656 15292 25684
rect 15286 25644 15292 25656
rect 15344 25644 15350 25696
rect 18874 25644 18880 25696
rect 18932 25684 18938 25696
rect 27798 25684 27804 25696
rect 18932 25656 27804 25684
rect 18932 25644 18938 25656
rect 27798 25644 27804 25656
rect 27856 25644 27862 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 7190 25480 7196 25492
rect 4540 25452 7196 25480
rect 1581 25279 1639 25285
rect 1581 25245 1593 25279
rect 1627 25276 1639 25279
rect 2222 25276 2228 25288
rect 1627 25248 2228 25276
rect 1627 25245 1639 25248
rect 1581 25239 1639 25245
rect 2222 25236 2228 25248
rect 2280 25236 2286 25288
rect 2317 25279 2375 25285
rect 2317 25245 2329 25279
rect 2363 25276 2375 25279
rect 3602 25276 3608 25288
rect 2363 25248 3608 25276
rect 2363 25245 2375 25248
rect 2317 25239 2375 25245
rect 3602 25236 3608 25248
rect 3660 25236 3666 25288
rect 4540 25285 4568 25452
rect 7190 25440 7196 25452
rect 7248 25440 7254 25492
rect 10686 25480 10692 25492
rect 10647 25452 10692 25480
rect 10686 25440 10692 25452
rect 10744 25440 10750 25492
rect 20073 25483 20131 25489
rect 20073 25449 20085 25483
rect 20119 25480 20131 25483
rect 20806 25480 20812 25492
rect 20119 25452 20812 25480
rect 20119 25449 20131 25452
rect 20073 25443 20131 25449
rect 20806 25440 20812 25452
rect 20864 25440 20870 25492
rect 29917 25483 29975 25489
rect 29917 25449 29929 25483
rect 29963 25480 29975 25483
rect 38010 25480 38016 25492
rect 29963 25452 38016 25480
rect 29963 25449 29975 25452
rect 29917 25443 29975 25449
rect 38010 25440 38016 25452
rect 38068 25440 38074 25492
rect 5353 25415 5411 25421
rect 5353 25381 5365 25415
rect 5399 25412 5411 25415
rect 7926 25412 7932 25424
rect 5399 25384 7932 25412
rect 5399 25381 5411 25384
rect 5353 25375 5411 25381
rect 7926 25372 7932 25384
rect 7984 25372 7990 25424
rect 11422 25372 11428 25424
rect 11480 25412 11486 25424
rect 11480 25384 15516 25412
rect 11480 25372 11486 25384
rect 6178 25344 6184 25356
rect 6139 25316 6184 25344
rect 6178 25304 6184 25316
rect 6236 25304 6242 25356
rect 13630 25344 13636 25356
rect 13591 25316 13636 25344
rect 13630 25304 13636 25316
rect 13688 25304 13694 25356
rect 15488 25344 15516 25384
rect 16114 25344 16120 25356
rect 15488 25316 16120 25344
rect 4525 25279 4583 25285
rect 4525 25245 4537 25279
rect 4571 25245 4583 25279
rect 4525 25239 4583 25245
rect 5537 25279 5595 25285
rect 5537 25245 5549 25279
rect 5583 25276 5595 25279
rect 5626 25276 5632 25288
rect 5583 25248 5632 25276
rect 5583 25245 5595 25248
rect 5537 25239 5595 25245
rect 1302 25168 1308 25220
rect 1360 25208 1366 25220
rect 5552 25208 5580 25239
rect 5626 25236 5632 25248
rect 5684 25236 5690 25288
rect 5997 25279 6055 25285
rect 5997 25245 6009 25279
rect 6043 25276 6055 25279
rect 6270 25276 6276 25288
rect 6043 25248 6276 25276
rect 6043 25245 6055 25248
rect 5997 25239 6055 25245
rect 6270 25236 6276 25248
rect 6328 25236 6334 25288
rect 6362 25236 6368 25288
rect 6420 25276 6426 25288
rect 7101 25279 7159 25285
rect 7101 25276 7113 25279
rect 6420 25248 7113 25276
rect 6420 25236 6426 25248
rect 7101 25245 7113 25248
rect 7147 25245 7159 25279
rect 9122 25276 9128 25288
rect 9083 25248 9128 25276
rect 7101 25239 7159 25245
rect 9122 25236 9128 25248
rect 9180 25236 9186 25288
rect 10870 25276 10876 25288
rect 10831 25248 10876 25276
rect 10870 25236 10876 25248
rect 10928 25236 10934 25288
rect 15105 25279 15163 25285
rect 15105 25245 15117 25279
rect 15151 25276 15163 25279
rect 15470 25276 15476 25288
rect 15151 25248 15476 25276
rect 15151 25245 15163 25248
rect 15105 25239 15163 25245
rect 15470 25236 15476 25248
rect 15528 25236 15534 25288
rect 15580 25285 15608 25316
rect 16114 25304 16120 25316
rect 16172 25304 16178 25356
rect 16298 25344 16304 25356
rect 16259 25316 16304 25344
rect 16298 25304 16304 25316
rect 16356 25304 16362 25356
rect 16942 25344 16948 25356
rect 16903 25316 16948 25344
rect 16942 25304 16948 25316
rect 17000 25304 17006 25356
rect 15565 25279 15623 25285
rect 15565 25245 15577 25279
rect 15611 25245 15623 25279
rect 15565 25239 15623 25245
rect 18693 25279 18751 25285
rect 18693 25245 18705 25279
rect 18739 25276 18751 25279
rect 19242 25276 19248 25288
rect 18739 25248 19248 25276
rect 18739 25245 18751 25248
rect 18693 25239 18751 25245
rect 19242 25236 19248 25248
rect 19300 25276 19306 25288
rect 19981 25279 20039 25285
rect 19981 25276 19993 25279
rect 19300 25248 19993 25276
rect 19300 25236 19306 25248
rect 19981 25245 19993 25248
rect 20027 25245 20039 25279
rect 19981 25239 20039 25245
rect 21453 25279 21511 25285
rect 21453 25245 21465 25279
rect 21499 25276 21511 25279
rect 26142 25276 26148 25288
rect 21499 25248 26148 25276
rect 21499 25245 21511 25248
rect 21453 25239 21511 25245
rect 26142 25236 26148 25248
rect 26200 25236 26206 25288
rect 30098 25276 30104 25288
rect 30059 25248 30104 25276
rect 30098 25236 30104 25248
rect 30156 25236 30162 25288
rect 1360 25180 5580 25208
rect 6641 25211 6699 25217
rect 1360 25168 1366 25180
rect 6641 25177 6653 25211
rect 6687 25208 6699 25211
rect 7742 25208 7748 25220
rect 6687 25180 7748 25208
rect 6687 25177 6699 25180
rect 6641 25171 6699 25177
rect 7742 25168 7748 25180
rect 7800 25168 7806 25220
rect 8018 25168 8024 25220
rect 8076 25208 8082 25220
rect 9217 25211 9275 25217
rect 9217 25208 9229 25211
rect 8076 25180 9229 25208
rect 8076 25168 8082 25180
rect 9217 25177 9229 25180
rect 9263 25177 9275 25211
rect 9217 25171 9275 25177
rect 12253 25211 12311 25217
rect 12253 25177 12265 25211
rect 12299 25208 12311 25211
rect 12989 25211 13047 25217
rect 12989 25208 13001 25211
rect 12299 25180 13001 25208
rect 12299 25177 12311 25180
rect 12253 25171 12311 25177
rect 12989 25177 13001 25180
rect 13035 25177 13047 25211
rect 12989 25171 13047 25177
rect 13081 25211 13139 25217
rect 13081 25177 13093 25211
rect 13127 25208 13139 25211
rect 15286 25208 15292 25220
rect 13127 25180 15292 25208
rect 13127 25177 13139 25180
rect 13081 25171 13139 25177
rect 15286 25168 15292 25180
rect 15344 25168 15350 25220
rect 16393 25211 16451 25217
rect 16393 25177 16405 25211
rect 16439 25208 16451 25211
rect 16574 25208 16580 25220
rect 16439 25180 16580 25208
rect 16439 25177 16451 25180
rect 16393 25171 16451 25177
rect 16574 25168 16580 25180
rect 16632 25168 16638 25220
rect 1762 25140 1768 25152
rect 1723 25112 1768 25140
rect 1762 25100 1768 25112
rect 1820 25100 1826 25152
rect 1854 25100 1860 25152
rect 1912 25140 1918 25152
rect 2409 25143 2467 25149
rect 2409 25140 2421 25143
rect 1912 25112 2421 25140
rect 1912 25100 1918 25112
rect 2409 25109 2421 25112
rect 2455 25109 2467 25143
rect 2409 25103 2467 25109
rect 2866 25100 2872 25152
rect 2924 25140 2930 25152
rect 2961 25143 3019 25149
rect 2961 25140 2973 25143
rect 2924 25112 2973 25140
rect 2924 25100 2930 25112
rect 2961 25109 2973 25112
rect 3007 25109 3019 25143
rect 2961 25103 3019 25109
rect 4617 25143 4675 25149
rect 4617 25109 4629 25143
rect 4663 25140 4675 25143
rect 4890 25140 4896 25152
rect 4663 25112 4896 25140
rect 4663 25109 4675 25112
rect 4617 25103 4675 25109
rect 4890 25100 4896 25112
rect 4948 25100 4954 25152
rect 6730 25100 6736 25152
rect 6788 25140 6794 25152
rect 7193 25143 7251 25149
rect 7193 25140 7205 25143
rect 6788 25112 7205 25140
rect 6788 25100 6794 25112
rect 7193 25109 7205 25112
rect 7239 25109 7251 25143
rect 8110 25140 8116 25152
rect 8071 25112 8116 25140
rect 7193 25103 7251 25109
rect 8110 25100 8116 25112
rect 8168 25100 8174 25152
rect 14277 25143 14335 25149
rect 14277 25109 14289 25143
rect 14323 25140 14335 25143
rect 14366 25140 14372 25152
rect 14323 25112 14372 25140
rect 14323 25109 14335 25112
rect 14277 25103 14335 25109
rect 14366 25100 14372 25112
rect 14424 25100 14430 25152
rect 14458 25100 14464 25152
rect 14516 25140 14522 25152
rect 14921 25143 14979 25149
rect 14921 25140 14933 25143
rect 14516 25112 14933 25140
rect 14516 25100 14522 25112
rect 14921 25109 14933 25112
rect 14967 25109 14979 25143
rect 14921 25103 14979 25109
rect 15194 25100 15200 25152
rect 15252 25140 15258 25152
rect 15657 25143 15715 25149
rect 15657 25140 15669 25143
rect 15252 25112 15669 25140
rect 15252 25100 15258 25112
rect 15657 25109 15669 25112
rect 15703 25109 15715 25143
rect 15657 25103 15715 25109
rect 17954 25100 17960 25152
rect 18012 25140 18018 25152
rect 18785 25143 18843 25149
rect 18785 25140 18797 25143
rect 18012 25112 18797 25140
rect 18012 25100 18018 25112
rect 18785 25109 18797 25112
rect 18831 25109 18843 25143
rect 18785 25103 18843 25109
rect 20806 25100 20812 25152
rect 20864 25140 20870 25152
rect 21545 25143 21603 25149
rect 21545 25140 21557 25143
rect 20864 25112 21557 25140
rect 20864 25100 20870 25112
rect 21545 25109 21557 25112
rect 21591 25109 21603 25143
rect 21545 25103 21603 25109
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 4798 24936 4804 24948
rect 4632 24908 4804 24936
rect 1949 24803 2007 24809
rect 1949 24769 1961 24803
rect 1995 24800 2007 24803
rect 2038 24800 2044 24812
rect 1995 24772 2044 24800
rect 1995 24769 2007 24772
rect 1949 24763 2007 24769
rect 2038 24760 2044 24772
rect 2096 24760 2102 24812
rect 3329 24803 3387 24809
rect 3329 24769 3341 24803
rect 3375 24800 3387 24803
rect 3878 24800 3884 24812
rect 3375 24772 3884 24800
rect 3375 24769 3387 24772
rect 3329 24763 3387 24769
rect 3878 24760 3884 24772
rect 3936 24800 3942 24812
rect 4632 24809 4660 24908
rect 4798 24896 4804 24908
rect 4856 24936 4862 24948
rect 4856 24908 9674 24936
rect 4856 24896 4862 24908
rect 4709 24871 4767 24877
rect 4709 24837 4721 24871
rect 4755 24868 4767 24871
rect 4755 24840 5396 24868
rect 4755 24837 4767 24840
rect 4709 24831 4767 24837
rect 3973 24803 4031 24809
rect 3973 24800 3985 24803
rect 3936 24772 3985 24800
rect 3936 24760 3942 24772
rect 3973 24769 3985 24772
rect 4019 24769 4031 24803
rect 3973 24763 4031 24769
rect 4617 24803 4675 24809
rect 4617 24769 4629 24803
rect 4663 24769 4675 24803
rect 5261 24803 5319 24809
rect 5261 24800 5273 24803
rect 4617 24763 4675 24769
rect 4724 24772 5273 24800
rect 2406 24692 2412 24744
rect 2464 24732 2470 24744
rect 2501 24735 2559 24741
rect 2501 24732 2513 24735
rect 2464 24704 2513 24732
rect 2464 24692 2470 24704
rect 2501 24701 2513 24704
rect 2547 24701 2559 24735
rect 2501 24695 2559 24701
rect 2958 24692 2964 24744
rect 3016 24732 3022 24744
rect 4724 24732 4752 24772
rect 5261 24769 5273 24772
rect 5307 24769 5319 24803
rect 5368 24800 5396 24840
rect 5534 24800 5540 24812
rect 5368 24772 5540 24800
rect 5261 24763 5319 24769
rect 5534 24760 5540 24772
rect 5592 24760 5598 24812
rect 8021 24803 8079 24809
rect 8021 24769 8033 24803
rect 8067 24800 8079 24803
rect 8110 24800 8116 24812
rect 8067 24772 8116 24800
rect 8067 24769 8079 24772
rect 8021 24763 8079 24769
rect 8110 24760 8116 24772
rect 8168 24760 8174 24812
rect 8202 24760 8208 24812
rect 8260 24800 8266 24812
rect 9309 24803 9367 24809
rect 8260 24772 8305 24800
rect 8260 24760 8266 24772
rect 9309 24769 9321 24803
rect 9355 24769 9367 24803
rect 9309 24763 9367 24769
rect 3016 24704 4752 24732
rect 5353 24735 5411 24741
rect 3016 24692 3022 24704
rect 5353 24701 5365 24735
rect 5399 24732 5411 24735
rect 6822 24732 6828 24744
rect 5399 24704 6828 24732
rect 5399 24701 5411 24704
rect 5353 24695 5411 24701
rect 6822 24692 6828 24704
rect 6880 24692 6886 24744
rect 7006 24732 7012 24744
rect 6967 24704 7012 24732
rect 7006 24692 7012 24704
rect 7064 24692 7070 24744
rect 7926 24692 7932 24744
rect 7984 24732 7990 24744
rect 9324 24732 9352 24763
rect 7984 24704 9352 24732
rect 9646 24732 9674 24908
rect 10134 24896 10140 24948
rect 10192 24936 10198 24948
rect 10778 24936 10784 24948
rect 10192 24908 10784 24936
rect 10192 24896 10198 24908
rect 10778 24896 10784 24908
rect 10836 24896 10842 24948
rect 15286 24936 15292 24948
rect 13188 24908 15292 24936
rect 10042 24800 10048 24812
rect 10003 24772 10048 24800
rect 10042 24760 10048 24772
rect 10100 24760 10106 24812
rect 10870 24760 10876 24812
rect 10928 24800 10934 24812
rect 13188 24800 13216 24908
rect 15286 24896 15292 24908
rect 15344 24896 15350 24948
rect 13449 24871 13507 24877
rect 13449 24837 13461 24871
rect 13495 24868 13507 24871
rect 14734 24868 14740 24880
rect 13495 24840 14740 24868
rect 13495 24837 13507 24840
rect 13449 24831 13507 24837
rect 14734 24828 14740 24840
rect 14792 24828 14798 24880
rect 15194 24868 15200 24880
rect 15155 24840 15200 24868
rect 15194 24828 15200 24840
rect 15252 24828 15258 24880
rect 17954 24868 17960 24880
rect 17915 24840 17960 24868
rect 17954 24828 17960 24840
rect 18012 24828 18018 24880
rect 10928 24772 13216 24800
rect 15749 24803 15807 24809
rect 10928 24760 10934 24772
rect 15749 24769 15761 24803
rect 15795 24800 15807 24803
rect 16942 24800 16948 24812
rect 15795 24772 16948 24800
rect 15795 24769 15807 24772
rect 15749 24763 15807 24769
rect 16942 24760 16948 24772
rect 17000 24760 17006 24812
rect 17037 24803 17095 24809
rect 17037 24769 17049 24803
rect 17083 24769 17095 24803
rect 17037 24763 17095 24769
rect 11514 24732 11520 24744
rect 9646 24704 11520 24732
rect 7984 24692 7990 24704
rect 11514 24692 11520 24704
rect 11572 24692 11578 24744
rect 13354 24732 13360 24744
rect 13315 24704 13360 24732
rect 13354 24692 13360 24704
rect 13412 24692 13418 24744
rect 14369 24735 14427 24741
rect 14369 24701 14381 24735
rect 14415 24732 14427 24735
rect 14826 24732 14832 24744
rect 14415 24704 14832 24732
rect 14415 24701 14427 24704
rect 14369 24695 14427 24701
rect 14826 24692 14832 24704
rect 14884 24692 14890 24744
rect 14918 24692 14924 24744
rect 14976 24732 14982 24744
rect 15105 24735 15163 24741
rect 15105 24732 15117 24735
rect 14976 24704 15117 24732
rect 14976 24692 14982 24704
rect 15105 24701 15117 24704
rect 15151 24701 15163 24735
rect 15105 24695 15163 24701
rect 15286 24692 15292 24744
rect 15344 24732 15350 24744
rect 16206 24732 16212 24744
rect 15344 24704 16212 24732
rect 15344 24692 15350 24704
rect 16206 24692 16212 24704
rect 16264 24732 16270 24744
rect 17052 24732 17080 24763
rect 32674 24760 32680 24812
rect 32732 24800 32738 24812
rect 38013 24803 38071 24809
rect 38013 24800 38025 24803
rect 32732 24772 38025 24800
rect 32732 24760 32738 24772
rect 38013 24769 38025 24772
rect 38059 24769 38071 24803
rect 38013 24763 38071 24769
rect 16264 24704 17080 24732
rect 16264 24692 16270 24704
rect 17586 24692 17592 24744
rect 17644 24732 17650 24744
rect 17862 24732 17868 24744
rect 17644 24704 17868 24732
rect 17644 24692 17650 24704
rect 17862 24692 17868 24704
rect 17920 24692 17926 24744
rect 18690 24732 18696 24744
rect 18651 24704 18696 24732
rect 18690 24692 18696 24704
rect 18748 24692 18754 24744
rect 8202 24664 8208 24676
rect 6748 24636 8208 24664
rect 934 24556 940 24608
rect 992 24596 998 24608
rect 1765 24599 1823 24605
rect 1765 24596 1777 24599
rect 992 24568 1777 24596
rect 992 24556 998 24568
rect 1765 24565 1777 24568
rect 1811 24565 1823 24599
rect 3418 24596 3424 24608
rect 3379 24568 3424 24596
rect 1765 24559 1823 24565
rect 3418 24556 3424 24568
rect 3476 24556 3482 24608
rect 4065 24599 4123 24605
rect 4065 24565 4077 24599
rect 4111 24596 4123 24599
rect 6748 24596 6776 24636
rect 8202 24624 8208 24636
rect 8260 24624 8266 24676
rect 8294 24624 8300 24676
rect 8352 24664 8358 24676
rect 8389 24667 8447 24673
rect 8389 24664 8401 24667
rect 8352 24636 8401 24664
rect 8352 24624 8358 24636
rect 8389 24633 8401 24636
rect 8435 24633 8447 24667
rect 8389 24627 8447 24633
rect 8846 24624 8852 24676
rect 8904 24664 8910 24676
rect 10686 24664 10692 24676
rect 8904 24636 10692 24664
rect 8904 24624 8910 24636
rect 10686 24624 10692 24636
rect 10744 24664 10750 24676
rect 10870 24664 10876 24676
rect 10744 24636 10876 24664
rect 10744 24624 10750 24636
rect 10870 24624 10876 24636
rect 10928 24624 10934 24676
rect 12710 24624 12716 24676
rect 12768 24664 12774 24676
rect 17954 24664 17960 24676
rect 12768 24636 17960 24664
rect 12768 24624 12774 24636
rect 17954 24624 17960 24636
rect 18012 24624 18018 24676
rect 9122 24596 9128 24608
rect 4111 24568 6776 24596
rect 9083 24568 9128 24596
rect 4111 24565 4123 24568
rect 4065 24559 4123 24565
rect 9122 24556 9128 24568
rect 9180 24556 9186 24608
rect 9490 24556 9496 24608
rect 9548 24596 9554 24608
rect 9861 24599 9919 24605
rect 9861 24596 9873 24599
rect 9548 24568 9873 24596
rect 9548 24556 9554 24568
rect 9861 24565 9873 24568
rect 9907 24565 9919 24599
rect 9861 24559 9919 24565
rect 11054 24556 11060 24608
rect 11112 24596 11118 24608
rect 12066 24596 12072 24608
rect 11112 24568 12072 24596
rect 11112 24556 11118 24568
rect 12066 24556 12072 24568
rect 12124 24596 12130 24608
rect 15286 24596 15292 24608
rect 12124 24568 15292 24596
rect 12124 24556 12130 24568
rect 15286 24556 15292 24568
rect 15344 24556 15350 24608
rect 15470 24556 15476 24608
rect 15528 24596 15534 24608
rect 16853 24599 16911 24605
rect 16853 24596 16865 24599
rect 15528 24568 16865 24596
rect 15528 24556 15534 24568
rect 16853 24565 16865 24568
rect 16899 24565 16911 24599
rect 38194 24596 38200 24608
rect 38155 24568 38200 24596
rect 16853 24559 16911 24565
rect 38194 24556 38200 24568
rect 38252 24556 38258 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 5905 24395 5963 24401
rect 5905 24392 5917 24395
rect 1596 24364 5917 24392
rect 1596 24197 1624 24364
rect 5905 24361 5917 24364
rect 5951 24361 5963 24395
rect 5905 24355 5963 24361
rect 6454 24352 6460 24404
rect 6512 24392 6518 24404
rect 8846 24392 8852 24404
rect 6512 24364 8852 24392
rect 6512 24352 6518 24364
rect 8846 24352 8852 24364
rect 8904 24352 8910 24404
rect 9030 24352 9036 24404
rect 9088 24392 9094 24404
rect 9125 24395 9183 24401
rect 9125 24392 9137 24395
rect 9088 24364 9137 24392
rect 9088 24352 9094 24364
rect 9125 24361 9137 24364
rect 9171 24361 9183 24395
rect 12710 24392 12716 24404
rect 9125 24355 9183 24361
rect 9646 24364 12716 24392
rect 3970 24284 3976 24336
rect 4028 24284 4034 24336
rect 4065 24327 4123 24333
rect 4065 24293 4077 24327
rect 4111 24324 4123 24327
rect 4111 24296 6040 24324
rect 4111 24293 4123 24296
rect 4065 24287 4123 24293
rect 3988 24256 4016 24284
rect 2516 24228 4292 24256
rect 2516 24197 2544 24228
rect 1581 24191 1639 24197
rect 1581 24157 1593 24191
rect 1627 24157 1639 24191
rect 1581 24151 1639 24157
rect 2501 24191 2559 24197
rect 2501 24157 2513 24191
rect 2547 24157 2559 24191
rect 2501 24151 2559 24157
rect 3145 24191 3203 24197
rect 3145 24157 3157 24191
rect 3191 24188 3203 24191
rect 3510 24188 3516 24200
rect 3191 24160 3516 24188
rect 3191 24157 3203 24160
rect 3145 24151 3203 24157
rect 1026 24080 1032 24132
rect 1084 24120 1090 24132
rect 2516 24120 2544 24151
rect 3510 24148 3516 24160
rect 3568 24148 3574 24200
rect 3970 24188 3976 24200
rect 3931 24160 3976 24188
rect 3970 24148 3976 24160
rect 4028 24148 4034 24200
rect 4264 24188 4292 24228
rect 4617 24191 4675 24197
rect 4617 24188 4629 24191
rect 4264 24160 4629 24188
rect 4617 24157 4629 24160
rect 4663 24157 4675 24191
rect 4617 24151 4675 24157
rect 4798 24148 4804 24200
rect 4856 24188 4862 24200
rect 5261 24191 5319 24197
rect 5261 24188 5273 24191
rect 4856 24160 5273 24188
rect 4856 24148 4862 24160
rect 5261 24157 5273 24160
rect 5307 24157 5319 24191
rect 5261 24151 5319 24157
rect 1084 24092 2544 24120
rect 4709 24123 4767 24129
rect 1084 24080 1090 24092
rect 4709 24089 4721 24123
rect 4755 24120 4767 24123
rect 5626 24120 5632 24132
rect 4755 24092 5632 24120
rect 4755 24089 4767 24092
rect 4709 24083 4767 24089
rect 5626 24080 5632 24092
rect 5684 24080 5690 24132
rect 1762 24052 1768 24064
rect 1723 24024 1768 24052
rect 1762 24012 1768 24024
rect 1820 24012 1826 24064
rect 2498 24012 2504 24064
rect 2556 24052 2562 24064
rect 2593 24055 2651 24061
rect 2593 24052 2605 24055
rect 2556 24024 2605 24052
rect 2556 24012 2562 24024
rect 2593 24021 2605 24024
rect 2639 24021 2651 24055
rect 2593 24015 2651 24021
rect 2958 24012 2964 24064
rect 3016 24052 3022 24064
rect 3237 24055 3295 24061
rect 3237 24052 3249 24055
rect 3016 24024 3249 24052
rect 3016 24012 3022 24024
rect 3237 24021 3249 24024
rect 3283 24021 3295 24055
rect 3237 24015 3295 24021
rect 5353 24055 5411 24061
rect 5353 24021 5365 24055
rect 5399 24052 5411 24055
rect 5810 24052 5816 24064
rect 5399 24024 5816 24052
rect 5399 24021 5411 24024
rect 5353 24015 5411 24021
rect 5810 24012 5816 24024
rect 5868 24012 5874 24064
rect 6012 24052 6040 24296
rect 6822 24284 6828 24336
rect 6880 24324 6886 24336
rect 7374 24324 7380 24336
rect 6880 24296 7380 24324
rect 6880 24284 6886 24296
rect 7374 24284 7380 24296
rect 7432 24284 7438 24336
rect 7558 24284 7564 24336
rect 7616 24324 7622 24336
rect 9646 24324 9674 24364
rect 12710 24352 12716 24364
rect 12768 24352 12774 24404
rect 19058 24352 19064 24404
rect 19116 24392 19122 24404
rect 19429 24395 19487 24401
rect 19429 24392 19441 24395
rect 19116 24364 19441 24392
rect 19116 24352 19122 24364
rect 19429 24361 19441 24364
rect 19475 24361 19487 24395
rect 20346 24392 20352 24404
rect 20307 24364 20352 24392
rect 19429 24355 19487 24361
rect 20346 24352 20352 24364
rect 20404 24352 20410 24404
rect 15654 24324 15660 24336
rect 7616 24296 9674 24324
rect 13372 24296 15660 24324
rect 7616 24284 7622 24296
rect 7006 24256 7012 24268
rect 6967 24228 7012 24256
rect 7006 24216 7012 24228
rect 7064 24216 7070 24268
rect 7466 24216 7472 24268
rect 7524 24256 7530 24268
rect 7524 24228 8248 24256
rect 7524 24216 7530 24228
rect 8220 24200 8248 24228
rect 8754 24216 8760 24268
rect 8812 24256 8818 24268
rect 13372 24256 13400 24296
rect 15654 24284 15660 24296
rect 15712 24284 15718 24336
rect 16482 24284 16488 24336
rect 16540 24324 16546 24336
rect 18601 24327 18659 24333
rect 18601 24324 18613 24327
rect 16540 24296 18613 24324
rect 16540 24284 16546 24296
rect 18601 24293 18613 24296
rect 18647 24324 18659 24327
rect 23290 24324 23296 24336
rect 18647 24296 23296 24324
rect 18647 24293 18659 24296
rect 18601 24287 18659 24293
rect 23290 24284 23296 24296
rect 23348 24284 23354 24336
rect 8812 24228 13400 24256
rect 13449 24259 13507 24265
rect 8812 24216 8818 24228
rect 13449 24225 13461 24259
rect 13495 24256 13507 24259
rect 13630 24256 13636 24268
rect 13495 24228 13636 24256
rect 13495 24225 13507 24228
rect 13449 24219 13507 24225
rect 13630 24216 13636 24228
rect 13688 24216 13694 24268
rect 14366 24256 14372 24268
rect 14327 24228 14372 24256
rect 14366 24216 14372 24228
rect 14424 24216 14430 24268
rect 14826 24256 14832 24268
rect 14787 24228 14832 24256
rect 14826 24216 14832 24228
rect 14884 24216 14890 24268
rect 15286 24216 15292 24268
rect 15344 24256 15350 24268
rect 16669 24259 16727 24265
rect 16669 24256 16681 24259
rect 15344 24228 16681 24256
rect 15344 24216 15350 24228
rect 16669 24225 16681 24228
rect 16715 24225 16727 24259
rect 30098 24256 30104 24268
rect 16669 24219 16727 24225
rect 18524 24228 30104 24256
rect 18524 24200 18552 24228
rect 30098 24216 30104 24228
rect 30156 24216 30162 24268
rect 6089 24191 6147 24197
rect 6089 24157 6101 24191
rect 6135 24188 6147 24191
rect 6822 24188 6828 24200
rect 6135 24160 6828 24188
rect 6135 24157 6147 24160
rect 6089 24151 6147 24157
rect 6822 24148 6828 24160
rect 6880 24148 6886 24200
rect 7650 24148 7656 24200
rect 7708 24188 7714 24200
rect 8202 24188 8208 24200
rect 7708 24160 7753 24188
rect 8115 24160 8208 24188
rect 7708 24148 7714 24160
rect 8202 24148 8208 24160
rect 8260 24148 8266 24200
rect 8662 24148 8668 24200
rect 8720 24188 8726 24200
rect 9309 24191 9367 24197
rect 9309 24188 9321 24191
rect 8720 24160 9321 24188
rect 8720 24148 8726 24160
rect 9309 24157 9321 24160
rect 9355 24157 9367 24191
rect 9309 24151 9367 24157
rect 10045 24191 10103 24197
rect 10045 24157 10057 24191
rect 10091 24188 10103 24191
rect 10410 24188 10416 24200
rect 10091 24160 10416 24188
rect 10091 24157 10103 24160
rect 10045 24151 10103 24157
rect 10410 24148 10416 24160
rect 10468 24148 10474 24200
rect 11057 24191 11115 24197
rect 11057 24157 11069 24191
rect 11103 24188 11115 24191
rect 12526 24188 12532 24200
rect 11103 24160 12532 24188
rect 11103 24157 11115 24160
rect 11057 24151 11115 24157
rect 12526 24148 12532 24160
rect 12584 24148 12590 24200
rect 15841 24191 15899 24197
rect 15841 24157 15853 24191
rect 15887 24157 15899 24191
rect 15841 24151 15899 24157
rect 17497 24191 17555 24197
rect 17497 24157 17509 24191
rect 17543 24188 17555 24191
rect 18414 24188 18420 24200
rect 17543 24160 18420 24188
rect 17543 24157 17555 24160
rect 17497 24151 17555 24157
rect 6638 24080 6644 24132
rect 6696 24120 6702 24132
rect 7101 24123 7159 24129
rect 7101 24120 7113 24123
rect 6696 24092 7113 24120
rect 6696 24080 6702 24092
rect 7101 24089 7113 24092
rect 7147 24089 7159 24123
rect 7101 24083 7159 24089
rect 7190 24080 7196 24132
rect 7248 24120 7254 24132
rect 7668 24120 7696 24148
rect 8386 24120 8392 24132
rect 7248 24092 7696 24120
rect 8347 24092 8392 24120
rect 7248 24080 7254 24092
rect 8386 24080 8392 24092
rect 8444 24080 8450 24132
rect 9214 24080 9220 24132
rect 9272 24120 9278 24132
rect 12618 24120 12624 24132
rect 9272 24092 12624 24120
rect 9272 24080 9278 24092
rect 12618 24080 12624 24092
rect 12676 24080 12682 24132
rect 12802 24120 12808 24132
rect 12763 24092 12808 24120
rect 12802 24080 12808 24092
rect 12860 24080 12866 24132
rect 12897 24123 12955 24129
rect 12897 24089 12909 24123
rect 12943 24120 12955 24123
rect 14090 24120 14096 24132
rect 12943 24092 14096 24120
rect 12943 24089 12955 24092
rect 12897 24083 12955 24089
rect 14090 24080 14096 24092
rect 14148 24080 14154 24132
rect 14458 24080 14464 24132
rect 14516 24120 14522 24132
rect 15856 24120 15884 24151
rect 18414 24148 18420 24160
rect 18472 24148 18478 24200
rect 18506 24148 18512 24200
rect 18564 24188 18570 24200
rect 19613 24191 19671 24197
rect 18564 24160 18609 24188
rect 18564 24148 18570 24160
rect 19613 24157 19625 24191
rect 19659 24157 19671 24191
rect 19613 24151 19671 24157
rect 20257 24191 20315 24197
rect 20257 24157 20269 24191
rect 20303 24188 20315 24191
rect 21450 24188 21456 24200
rect 20303 24160 21456 24188
rect 20303 24157 20315 24160
rect 20257 24151 20315 24157
rect 16390 24120 16396 24132
rect 14516 24092 14561 24120
rect 14660 24092 15884 24120
rect 16351 24092 16396 24120
rect 14516 24080 14522 24092
rect 7466 24052 7472 24064
rect 6012 24024 7472 24052
rect 7466 24012 7472 24024
rect 7524 24012 7530 24064
rect 10137 24055 10195 24061
rect 10137 24021 10149 24055
rect 10183 24052 10195 24055
rect 10226 24052 10232 24064
rect 10183 24024 10232 24052
rect 10183 24021 10195 24024
rect 10137 24015 10195 24021
rect 10226 24012 10232 24024
rect 10284 24012 10290 24064
rect 11054 24012 11060 24064
rect 11112 24052 11118 24064
rect 11149 24055 11207 24061
rect 11149 24052 11161 24055
rect 11112 24024 11161 24052
rect 11112 24012 11118 24024
rect 11149 24021 11161 24024
rect 11195 24021 11207 24055
rect 11149 24015 11207 24021
rect 13906 24012 13912 24064
rect 13964 24052 13970 24064
rect 14660 24052 14688 24092
rect 16390 24080 16396 24092
rect 16448 24080 16454 24132
rect 16485 24123 16543 24129
rect 16485 24089 16497 24123
rect 16531 24089 16543 24123
rect 16485 24083 16543 24089
rect 13964 24024 14688 24052
rect 15657 24055 15715 24061
rect 13964 24012 13970 24024
rect 15657 24021 15669 24055
rect 15703 24052 15715 24055
rect 16500 24052 16528 24083
rect 17770 24080 17776 24132
rect 17828 24120 17834 24132
rect 19628 24120 19656 24151
rect 21450 24148 21456 24160
rect 21508 24148 21514 24200
rect 31021 24191 31079 24197
rect 31021 24157 31033 24191
rect 31067 24188 31079 24191
rect 34514 24188 34520 24200
rect 31067 24160 34520 24188
rect 31067 24157 31079 24160
rect 31021 24151 31079 24157
rect 34514 24148 34520 24160
rect 34572 24148 34578 24200
rect 37734 24148 37740 24200
rect 37792 24188 37798 24200
rect 38013 24191 38071 24197
rect 38013 24188 38025 24191
rect 37792 24160 38025 24188
rect 37792 24148 37798 24160
rect 38013 24157 38025 24160
rect 38059 24157 38071 24191
rect 38013 24151 38071 24157
rect 17828 24092 19656 24120
rect 17828 24080 17834 24092
rect 15703 24024 16528 24052
rect 15703 24021 15715 24024
rect 15657 24015 15715 24021
rect 16574 24012 16580 24064
rect 16632 24052 16638 24064
rect 17589 24055 17647 24061
rect 17589 24052 17601 24055
rect 16632 24024 17601 24052
rect 16632 24012 16638 24024
rect 17589 24021 17601 24024
rect 17635 24021 17647 24055
rect 31110 24052 31116 24064
rect 31071 24024 31116 24052
rect 17589 24015 17647 24021
rect 31110 24012 31116 24024
rect 31168 24012 31174 24064
rect 38194 24052 38200 24064
rect 38155 24024 38200 24052
rect 38194 24012 38200 24024
rect 38252 24012 38258 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 3878 23848 3884 23860
rect 2608 23820 3884 23848
rect 1670 23712 1676 23724
rect 1631 23684 1676 23712
rect 1670 23672 1676 23684
rect 1728 23672 1734 23724
rect 2608 23721 2636 23820
rect 3878 23808 3884 23820
rect 3936 23808 3942 23860
rect 3973 23851 4031 23857
rect 3973 23817 3985 23851
rect 4019 23848 4031 23851
rect 6638 23848 6644 23860
rect 4019 23820 6500 23848
rect 6599 23820 6644 23848
rect 4019 23817 4031 23820
rect 3973 23811 4031 23817
rect 6086 23780 6092 23792
rect 3988 23752 6092 23780
rect 2593 23715 2651 23721
rect 2593 23681 2605 23715
rect 2639 23681 2651 23715
rect 2593 23675 2651 23681
rect 3237 23715 3295 23721
rect 3237 23681 3249 23715
rect 3283 23712 3295 23715
rect 3602 23712 3608 23724
rect 3283 23684 3608 23712
rect 3283 23681 3295 23684
rect 3237 23675 3295 23681
rect 3602 23672 3608 23684
rect 3660 23672 3666 23724
rect 3881 23715 3939 23721
rect 3881 23681 3893 23715
rect 3927 23710 3939 23715
rect 3988 23710 4016 23752
rect 6086 23740 6092 23752
rect 6144 23740 6150 23792
rect 6472 23780 6500 23820
rect 6638 23808 6644 23820
rect 6696 23808 6702 23860
rect 6822 23808 6828 23860
rect 6880 23848 6886 23860
rect 7469 23851 7527 23857
rect 7469 23848 7481 23851
rect 6880 23820 7481 23848
rect 6880 23808 6886 23820
rect 7469 23817 7481 23820
rect 7515 23817 7527 23851
rect 7469 23811 7527 23817
rect 7742 23808 7748 23860
rect 7800 23848 7806 23860
rect 8849 23851 8907 23857
rect 8849 23848 8861 23851
rect 7800 23820 8861 23848
rect 7800 23808 7806 23820
rect 8849 23817 8861 23820
rect 8895 23817 8907 23851
rect 8849 23811 8907 23817
rect 9953 23851 10011 23857
rect 9953 23817 9965 23851
rect 9999 23848 10011 23851
rect 11146 23848 11152 23860
rect 9999 23820 11152 23848
rect 9999 23817 10011 23820
rect 9953 23811 10011 23817
rect 11146 23808 11152 23820
rect 11204 23808 11210 23860
rect 13357 23851 13415 23857
rect 13357 23817 13369 23851
rect 13403 23848 13415 23851
rect 13403 23820 17264 23848
rect 13403 23817 13415 23820
rect 13357 23811 13415 23817
rect 7006 23780 7012 23792
rect 6472 23752 7012 23780
rect 7006 23740 7012 23752
rect 7064 23740 7070 23792
rect 12434 23780 12440 23792
rect 7392 23752 12440 23780
rect 3927 23682 4016 23710
rect 3927 23681 3939 23682
rect 3881 23675 3939 23681
rect 4706 23672 4712 23724
rect 4764 23712 4770 23724
rect 5166 23712 5172 23724
rect 4764 23684 4809 23712
rect 5127 23684 5172 23712
rect 4764 23672 4770 23684
rect 5166 23672 5172 23684
rect 5224 23672 5230 23724
rect 5813 23715 5871 23721
rect 5813 23681 5825 23715
rect 5859 23712 5871 23715
rect 6454 23712 6460 23724
rect 5859 23684 6460 23712
rect 5859 23681 5871 23684
rect 5813 23675 5871 23681
rect 6454 23672 6460 23684
rect 6512 23672 6518 23724
rect 6549 23715 6607 23721
rect 6549 23681 6561 23715
rect 6595 23712 6607 23715
rect 7282 23712 7288 23724
rect 6595 23684 7288 23712
rect 6595 23681 6607 23684
rect 6549 23675 6607 23681
rect 7282 23672 7288 23684
rect 7340 23672 7346 23724
rect 7392 23721 7420 23752
rect 12434 23740 12440 23752
rect 12492 23740 12498 23792
rect 12526 23740 12532 23792
rect 12584 23780 12590 23792
rect 12894 23780 12900 23792
rect 12584 23752 12900 23780
rect 12584 23740 12590 23752
rect 12894 23740 12900 23752
rect 12952 23780 12958 23792
rect 15378 23780 15384 23792
rect 12952 23752 14596 23780
rect 15339 23752 15384 23780
rect 12952 23740 12958 23752
rect 7377 23715 7435 23721
rect 7377 23681 7389 23715
rect 7423 23681 7435 23715
rect 7377 23675 7435 23681
rect 7650 23672 7656 23724
rect 7708 23712 7714 23724
rect 8389 23715 8447 23721
rect 7708 23684 8340 23712
rect 7708 23672 7714 23684
rect 1857 23647 1915 23653
rect 1857 23613 1869 23647
rect 1903 23644 1915 23647
rect 7558 23644 7564 23656
rect 1903 23616 7564 23644
rect 1903 23613 1915 23616
rect 1857 23607 1915 23613
rect 7558 23604 7564 23616
rect 7616 23604 7622 23656
rect 8205 23647 8263 23653
rect 8205 23613 8217 23647
rect 8251 23613 8263 23647
rect 8312 23644 8340 23684
rect 8389 23681 8401 23715
rect 8435 23712 8447 23715
rect 9122 23712 9128 23724
rect 8435 23684 9128 23712
rect 8435 23681 8447 23684
rect 8389 23675 8447 23681
rect 9122 23672 9128 23684
rect 9180 23672 9186 23724
rect 9306 23712 9312 23724
rect 9267 23684 9312 23712
rect 9306 23672 9312 23684
rect 9364 23672 9370 23724
rect 9490 23712 9496 23724
rect 9451 23684 9496 23712
rect 9490 23672 9496 23684
rect 9548 23672 9554 23724
rect 10505 23715 10563 23721
rect 10505 23681 10517 23715
rect 10551 23712 10563 23715
rect 10594 23712 10600 23724
rect 10551 23684 10600 23712
rect 10551 23681 10563 23684
rect 10505 23675 10563 23681
rect 10594 23672 10600 23684
rect 10652 23672 10658 23724
rect 11698 23712 11704 23724
rect 11659 23684 11704 23712
rect 11698 23672 11704 23684
rect 11756 23712 11762 23724
rect 11756 23684 12434 23712
rect 11756 23672 11762 23684
rect 10870 23644 10876 23656
rect 8312 23616 10876 23644
rect 8205 23607 8263 23613
rect 3329 23579 3387 23585
rect 3329 23545 3341 23579
rect 3375 23576 3387 23579
rect 3375 23548 4752 23576
rect 3375 23545 3387 23548
rect 3329 23539 3387 23545
rect 4724 23520 4752 23548
rect 5810 23536 5816 23588
rect 5868 23576 5874 23588
rect 8220 23576 8248 23607
rect 10870 23604 10876 23616
rect 10928 23604 10934 23656
rect 12406 23644 12434 23684
rect 12618 23672 12624 23724
rect 12676 23712 12682 23724
rect 14568 23721 14596 23752
rect 15378 23740 15384 23752
rect 15436 23740 15442 23792
rect 15473 23783 15531 23789
rect 15473 23749 15485 23783
rect 15519 23780 15531 23783
rect 16574 23780 16580 23792
rect 15519 23752 16580 23780
rect 15519 23749 15531 23752
rect 15473 23743 15531 23749
rect 16574 23740 16580 23752
rect 16632 23740 16638 23792
rect 17236 23789 17264 23820
rect 22094 23808 22100 23860
rect 22152 23848 22158 23860
rect 32674 23848 32680 23860
rect 22152 23820 22197 23848
rect 32635 23820 32680 23848
rect 22152 23808 22158 23820
rect 32674 23808 32680 23820
rect 32732 23808 32738 23860
rect 17221 23783 17279 23789
rect 17221 23749 17233 23783
rect 17267 23749 17279 23783
rect 18966 23780 18972 23792
rect 18927 23752 18972 23780
rect 17221 23743 17279 23749
rect 18966 23740 18972 23752
rect 19024 23740 19030 23792
rect 22020 23752 31754 23780
rect 22020 23721 22048 23752
rect 13265 23715 13323 23721
rect 13265 23712 13277 23715
rect 12676 23684 13277 23712
rect 12676 23672 12682 23684
rect 13265 23681 13277 23684
rect 13311 23681 13323 23715
rect 13265 23675 13323 23681
rect 14093 23715 14151 23721
rect 14093 23681 14105 23715
rect 14139 23681 14151 23715
rect 14093 23675 14151 23681
rect 14553 23715 14611 23721
rect 14553 23681 14565 23715
rect 14599 23681 14611 23715
rect 14553 23675 14611 23681
rect 22005 23715 22063 23721
rect 22005 23681 22017 23715
rect 22051 23681 22063 23715
rect 23290 23712 23296 23724
rect 23251 23684 23296 23712
rect 22005 23675 22063 23681
rect 14108 23644 14136 23675
rect 23290 23672 23296 23684
rect 23348 23672 23354 23724
rect 24489 23715 24547 23721
rect 24489 23681 24501 23715
rect 24535 23712 24547 23715
rect 25406 23712 25412 23724
rect 24535 23684 25412 23712
rect 24535 23681 24547 23684
rect 24489 23675 24547 23681
rect 25406 23672 25412 23684
rect 25464 23672 25470 23724
rect 31726 23712 31754 23752
rect 32858 23712 32864 23724
rect 31726 23684 32864 23712
rect 32858 23672 32864 23684
rect 32916 23672 32922 23724
rect 14826 23644 14832 23656
rect 12406 23616 14136 23644
rect 14200 23616 14832 23644
rect 13906 23576 13912 23588
rect 5868 23548 7604 23576
rect 8220 23548 12434 23576
rect 13867 23548 13912 23576
rect 5868 23536 5874 23548
rect 2498 23468 2504 23520
rect 2556 23508 2562 23520
rect 2685 23511 2743 23517
rect 2685 23508 2697 23511
rect 2556 23480 2697 23508
rect 2556 23468 2562 23480
rect 2685 23477 2697 23480
rect 2731 23477 2743 23511
rect 2685 23471 2743 23477
rect 3878 23468 3884 23520
rect 3936 23508 3942 23520
rect 4525 23511 4583 23517
rect 4525 23508 4537 23511
rect 3936 23480 4537 23508
rect 3936 23468 3942 23480
rect 4525 23477 4537 23480
rect 4571 23477 4583 23511
rect 4525 23471 4583 23477
rect 4706 23468 4712 23520
rect 4764 23468 4770 23520
rect 5258 23508 5264 23520
rect 5219 23480 5264 23508
rect 5258 23468 5264 23480
rect 5316 23468 5322 23520
rect 5905 23511 5963 23517
rect 5905 23477 5917 23511
rect 5951 23508 5963 23511
rect 6638 23508 6644 23520
rect 5951 23480 6644 23508
rect 5951 23477 5963 23480
rect 5905 23471 5963 23477
rect 6638 23468 6644 23480
rect 6696 23468 6702 23520
rect 7576 23508 7604 23548
rect 9766 23508 9772 23520
rect 7576 23480 9772 23508
rect 9766 23468 9772 23480
rect 9824 23468 9830 23520
rect 10597 23511 10655 23517
rect 10597 23477 10609 23511
rect 10643 23508 10655 23511
rect 11606 23508 11612 23520
rect 10643 23480 11612 23508
rect 10643 23477 10655 23480
rect 10597 23471 10655 23477
rect 11606 23468 11612 23480
rect 11664 23468 11670 23520
rect 11790 23508 11796 23520
rect 11751 23480 11796 23508
rect 11790 23468 11796 23480
rect 11848 23468 11854 23520
rect 12406 23508 12434 23548
rect 13906 23536 13912 23548
rect 13964 23536 13970 23588
rect 14200 23508 14228 23616
rect 14826 23604 14832 23616
rect 14884 23604 14890 23656
rect 15654 23644 15660 23656
rect 15615 23616 15660 23644
rect 15654 23604 15660 23616
rect 15712 23604 15718 23656
rect 17129 23647 17187 23653
rect 17129 23613 17141 23647
rect 17175 23613 17187 23647
rect 18046 23644 18052 23656
rect 18007 23616 18052 23644
rect 17129 23607 17187 23613
rect 17144 23576 17172 23607
rect 18046 23604 18052 23616
rect 18104 23604 18110 23656
rect 18874 23644 18880 23656
rect 18835 23616 18880 23644
rect 18874 23604 18880 23616
rect 18932 23604 18938 23656
rect 19337 23647 19395 23653
rect 19337 23613 19349 23647
rect 19383 23613 19395 23647
rect 19337 23607 19395 23613
rect 23477 23647 23535 23653
rect 23477 23613 23489 23647
rect 23523 23644 23535 23647
rect 24581 23647 24639 23653
rect 24581 23644 24593 23647
rect 23523 23616 24593 23644
rect 23523 23613 23535 23616
rect 23477 23607 23535 23613
rect 24581 23613 24593 23616
rect 24627 23613 24639 23647
rect 24581 23607 24639 23613
rect 18598 23576 18604 23588
rect 17144 23548 18604 23576
rect 18598 23536 18604 23548
rect 18656 23536 18662 23588
rect 12406 23480 14228 23508
rect 14458 23468 14464 23520
rect 14516 23508 14522 23520
rect 14645 23511 14703 23517
rect 14645 23508 14657 23511
rect 14516 23480 14657 23508
rect 14516 23468 14522 23480
rect 14645 23477 14657 23480
rect 14691 23477 14703 23511
rect 14645 23471 14703 23477
rect 16390 23468 16396 23520
rect 16448 23508 16454 23520
rect 17310 23508 17316 23520
rect 16448 23480 17316 23508
rect 16448 23468 16454 23480
rect 17310 23468 17316 23480
rect 17368 23468 17374 23520
rect 18506 23468 18512 23520
rect 18564 23508 18570 23520
rect 19352 23508 19380 23607
rect 23934 23508 23940 23520
rect 18564 23480 19380 23508
rect 23895 23480 23940 23508
rect 18564 23468 18570 23480
rect 23934 23468 23940 23480
rect 23992 23468 23998 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 6089 23307 6147 23313
rect 6089 23273 6101 23307
rect 6135 23304 6147 23307
rect 6270 23304 6276 23316
rect 6135 23276 6276 23304
rect 6135 23273 6147 23276
rect 6089 23267 6147 23273
rect 6270 23264 6276 23276
rect 6328 23264 6334 23316
rect 10520 23276 17264 23304
rect 5629 23171 5687 23177
rect 4172 23140 5580 23168
rect 3237 23103 3295 23109
rect 3237 23069 3249 23103
rect 3283 23100 3295 23103
rect 3510 23100 3516 23112
rect 3283 23072 3516 23100
rect 3283 23069 3295 23072
rect 3237 23063 3295 23069
rect 3510 23060 3516 23072
rect 3568 23060 3574 23112
rect 4172 23109 4200 23140
rect 4157 23103 4215 23109
rect 4157 23069 4169 23103
rect 4203 23069 4215 23103
rect 4157 23063 4215 23069
rect 4614 23060 4620 23112
rect 4672 23100 4678 23112
rect 4801 23103 4859 23109
rect 4801 23100 4813 23103
rect 4672 23072 4813 23100
rect 4672 23060 4678 23072
rect 4801 23069 4813 23072
rect 4847 23069 4859 23103
rect 4801 23063 4859 23069
rect 5445 23103 5503 23109
rect 5445 23069 5457 23103
rect 5491 23069 5503 23103
rect 5552 23100 5580 23140
rect 5629 23137 5641 23171
rect 5675 23168 5687 23171
rect 6638 23168 6644 23180
rect 5675 23140 6644 23168
rect 5675 23137 5687 23140
rect 5629 23131 5687 23137
rect 6638 23128 6644 23140
rect 6696 23128 6702 23180
rect 9493 23171 9551 23177
rect 9493 23137 9505 23171
rect 9539 23168 9551 23171
rect 9674 23168 9680 23180
rect 9539 23140 9680 23168
rect 9539 23137 9551 23140
rect 9493 23131 9551 23137
rect 9674 23128 9680 23140
rect 9732 23128 9738 23180
rect 10520 23177 10548 23276
rect 13078 23236 13084 23248
rect 11808 23208 13084 23236
rect 10505 23171 10563 23177
rect 10505 23137 10517 23171
rect 10551 23137 10563 23171
rect 10505 23131 10563 23137
rect 6546 23100 6552 23112
rect 5552 23072 6552 23100
rect 5445 23063 5503 23069
rect 1765 23035 1823 23041
rect 1765 23032 1777 23035
rect 1688 23004 1777 23032
rect 1688 22976 1716 23004
rect 1765 23001 1777 23004
rect 1811 23001 1823 23035
rect 1765 22995 1823 23001
rect 1854 22992 1860 23044
rect 1912 23032 1918 23044
rect 2409 23035 2467 23041
rect 1912 23004 1957 23032
rect 1912 22992 1918 23004
rect 2409 23001 2421 23035
rect 2455 23032 2467 23035
rect 3602 23032 3608 23044
rect 2455 23004 3608 23032
rect 2455 23001 2467 23004
rect 2409 22995 2467 23001
rect 3602 22992 3608 23004
rect 3660 22992 3666 23044
rect 3970 22992 3976 23044
rect 4028 23032 4034 23044
rect 4893 23035 4951 23041
rect 4893 23032 4905 23035
rect 4028 23004 4905 23032
rect 4028 22992 4034 23004
rect 4893 23001 4905 23004
rect 4939 23001 4951 23035
rect 5460 23032 5488 23063
rect 6546 23060 6552 23072
rect 6604 23060 6610 23112
rect 7006 23060 7012 23112
rect 7064 23100 7070 23112
rect 7374 23100 7380 23112
rect 7064 23072 7380 23100
rect 7064 23060 7070 23072
rect 7374 23060 7380 23072
rect 7432 23060 7438 23112
rect 7742 23100 7748 23112
rect 7703 23072 7748 23100
rect 7742 23060 7748 23072
rect 7800 23060 7806 23112
rect 8386 23100 8392 23112
rect 8347 23072 8392 23100
rect 8386 23060 8392 23072
rect 8444 23060 8450 23112
rect 11057 23103 11115 23109
rect 11057 23069 11069 23103
rect 11103 23100 11115 23103
rect 11330 23100 11336 23112
rect 11103 23072 11336 23100
rect 11103 23069 11115 23072
rect 11057 23063 11115 23069
rect 11330 23060 11336 23072
rect 11388 23060 11394 23112
rect 11808 23109 11836 23208
rect 13078 23196 13084 23208
rect 13136 23196 13142 23248
rect 16482 23236 16488 23248
rect 14384 23208 16488 23236
rect 12529 23171 12587 23177
rect 12529 23137 12541 23171
rect 12575 23168 12587 23171
rect 13354 23168 13360 23180
rect 12575 23140 13360 23168
rect 12575 23137 12587 23140
rect 12529 23131 12587 23137
rect 13354 23128 13360 23140
rect 13412 23128 13418 23180
rect 14384 23177 14412 23208
rect 16482 23196 16488 23208
rect 16540 23196 16546 23248
rect 16758 23236 16764 23248
rect 16719 23208 16764 23236
rect 16758 23196 16764 23208
rect 16816 23196 16822 23248
rect 14369 23171 14427 23177
rect 14369 23137 14381 23171
rect 14415 23137 14427 23171
rect 14734 23168 14740 23180
rect 14695 23140 14740 23168
rect 14369 23131 14427 23137
rect 14734 23128 14740 23140
rect 14792 23128 14798 23180
rect 17236 23168 17264 23276
rect 17402 23264 17408 23316
rect 17460 23304 17466 23316
rect 17773 23307 17831 23313
rect 17773 23304 17785 23307
rect 17460 23276 17785 23304
rect 17460 23264 17466 23276
rect 17773 23273 17785 23276
rect 17819 23273 17831 23307
rect 17773 23267 17831 23273
rect 18417 23307 18475 23313
rect 18417 23273 18429 23307
rect 18463 23304 18475 23307
rect 18966 23304 18972 23316
rect 18463 23276 18972 23304
rect 18463 23273 18475 23276
rect 18417 23267 18475 23273
rect 18966 23264 18972 23276
rect 19024 23264 19030 23316
rect 17310 23196 17316 23248
rect 17368 23236 17374 23248
rect 27341 23239 27399 23245
rect 27341 23236 27353 23239
rect 17368 23208 27353 23236
rect 17368 23196 17374 23208
rect 27341 23205 27353 23208
rect 27387 23205 27399 23239
rect 27341 23199 27399 23205
rect 18874 23168 18880 23180
rect 17236 23140 18880 23168
rect 18874 23128 18880 23140
rect 18932 23128 18938 23180
rect 11793 23103 11851 23109
rect 11793 23069 11805 23103
rect 11839 23069 11851 23103
rect 11793 23063 11851 23069
rect 15010 23060 15016 23112
rect 15068 23100 15074 23112
rect 15473 23103 15531 23109
rect 15473 23100 15485 23103
rect 15068 23072 15485 23100
rect 15068 23060 15074 23072
rect 15473 23069 15485 23072
rect 15519 23069 15531 23103
rect 17586 23100 17592 23112
rect 15473 23063 15531 23069
rect 15580 23072 17592 23100
rect 7190 23032 7196 23044
rect 5460 23004 7196 23032
rect 4893 22995 4951 23001
rect 7190 22992 7196 23004
rect 7248 22992 7254 23044
rect 9582 22992 9588 23044
rect 9640 23032 9646 23044
rect 12621 23035 12679 23041
rect 9640 23004 9685 23032
rect 9640 22992 9646 23004
rect 12621 23001 12633 23035
rect 12667 23001 12679 23035
rect 12621 22995 12679 23001
rect 13541 23035 13599 23041
rect 13541 23001 13553 23035
rect 13587 23001 13599 23035
rect 13541 22995 13599 23001
rect 1670 22924 1676 22976
rect 1728 22924 1734 22976
rect 3329 22967 3387 22973
rect 3329 22933 3341 22967
rect 3375 22964 3387 22967
rect 4062 22964 4068 22976
rect 3375 22936 4068 22964
rect 3375 22933 3387 22936
rect 3329 22927 3387 22933
rect 4062 22924 4068 22936
rect 4120 22924 4126 22976
rect 4249 22967 4307 22973
rect 4249 22933 4261 22967
rect 4295 22964 4307 22967
rect 4614 22964 4620 22976
rect 4295 22936 4620 22964
rect 4295 22933 4307 22936
rect 4249 22927 4307 22933
rect 4614 22924 4620 22936
rect 4672 22924 4678 22976
rect 7101 22967 7159 22973
rect 7101 22933 7113 22967
rect 7147 22964 7159 22967
rect 7466 22964 7472 22976
rect 7147 22936 7472 22964
rect 7147 22933 7159 22936
rect 7101 22927 7159 22933
rect 7466 22924 7472 22936
rect 7524 22924 7530 22976
rect 7558 22924 7564 22976
rect 7616 22964 7622 22976
rect 7837 22967 7895 22973
rect 7837 22964 7849 22967
rect 7616 22936 7849 22964
rect 7616 22924 7622 22936
rect 7837 22933 7849 22936
rect 7883 22933 7895 22967
rect 7837 22927 7895 22933
rect 8481 22967 8539 22973
rect 8481 22933 8493 22967
rect 8527 22964 8539 22967
rect 9398 22964 9404 22976
rect 8527 22936 9404 22964
rect 8527 22933 8539 22936
rect 8481 22927 8539 22933
rect 9398 22924 9404 22936
rect 9456 22924 9462 22976
rect 11146 22964 11152 22976
rect 11107 22936 11152 22964
rect 11146 22924 11152 22936
rect 11204 22924 11210 22976
rect 11885 22967 11943 22973
rect 11885 22933 11897 22967
rect 11931 22964 11943 22967
rect 12636 22964 12664 22995
rect 11931 22936 12664 22964
rect 11931 22933 11943 22936
rect 11885 22927 11943 22933
rect 12710 22924 12716 22976
rect 12768 22964 12774 22976
rect 13556 22964 13584 22995
rect 14458 22992 14464 23044
rect 14516 23032 14522 23044
rect 15580 23032 15608 23072
rect 17586 23060 17592 23072
rect 17644 23060 17650 23112
rect 18322 23100 18328 23112
rect 18283 23072 18328 23100
rect 18322 23060 18328 23072
rect 18380 23060 18386 23112
rect 24765 23103 24823 23109
rect 24765 23069 24777 23103
rect 24811 23100 24823 23103
rect 24811 23072 25268 23100
rect 24811 23069 24823 23072
rect 24765 23063 24823 23069
rect 16574 23032 16580 23044
rect 14516 23004 14561 23032
rect 14660 23004 15608 23032
rect 16535 23004 16580 23032
rect 14516 22992 14522 23004
rect 14660 22964 14688 23004
rect 16574 22992 16580 23004
rect 16632 22992 16638 23044
rect 17678 23032 17684 23044
rect 17639 23004 17684 23032
rect 17678 22992 17684 23004
rect 17736 22992 17742 23044
rect 18138 22992 18144 23044
rect 18196 23032 18202 23044
rect 19426 23032 19432 23044
rect 18196 23004 19432 23032
rect 18196 22992 18202 23004
rect 19426 22992 19432 23004
rect 19484 22992 19490 23044
rect 12768 22936 14688 22964
rect 12768 22924 12774 22936
rect 15194 22924 15200 22976
rect 15252 22964 15258 22976
rect 15565 22967 15623 22973
rect 15565 22964 15577 22967
rect 15252 22936 15577 22964
rect 15252 22924 15258 22936
rect 15565 22933 15577 22936
rect 15611 22933 15623 22967
rect 15565 22927 15623 22933
rect 18874 22924 18880 22976
rect 18932 22964 18938 22976
rect 22370 22964 22376 22976
rect 18932 22936 22376 22964
rect 18932 22924 18938 22936
rect 22370 22924 22376 22936
rect 22428 22924 22434 22976
rect 22646 22924 22652 22976
rect 22704 22964 22710 22976
rect 25240 22973 25268 23072
rect 25406 23060 25412 23112
rect 25464 23100 25470 23112
rect 27249 23103 27307 23109
rect 25464 23072 25557 23100
rect 25464 23060 25470 23072
rect 27249 23069 27261 23103
rect 27295 23100 27307 23103
rect 37826 23100 37832 23112
rect 27295 23072 37832 23100
rect 27295 23069 27307 23072
rect 27249 23063 27307 23069
rect 37826 23060 37832 23072
rect 37884 23060 37890 23112
rect 25424 23032 25452 23060
rect 27982 23032 27988 23044
rect 25424 23004 27988 23032
rect 27982 22992 27988 23004
rect 28040 22992 28046 23044
rect 24581 22967 24639 22973
rect 24581 22964 24593 22967
rect 22704 22936 24593 22964
rect 22704 22924 22710 22936
rect 24581 22933 24593 22936
rect 24627 22933 24639 22967
rect 24581 22927 24639 22933
rect 25225 22967 25283 22973
rect 25225 22933 25237 22967
rect 25271 22933 25283 22967
rect 25225 22927 25283 22933
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 1854 22720 1860 22772
rect 1912 22760 1918 22772
rect 6730 22760 6736 22772
rect 1912 22732 6736 22760
rect 1912 22720 1918 22732
rect 6730 22720 6736 22732
rect 6788 22720 6794 22772
rect 6825 22763 6883 22769
rect 6825 22729 6837 22763
rect 6871 22760 6883 22763
rect 6871 22732 7604 22760
rect 6871 22729 6883 22732
rect 6825 22723 6883 22729
rect 1765 22695 1823 22701
rect 1765 22661 1777 22695
rect 1811 22692 1823 22695
rect 2682 22692 2688 22704
rect 1811 22664 2688 22692
rect 1811 22661 1823 22664
rect 1765 22655 1823 22661
rect 2682 22652 2688 22664
rect 2740 22652 2746 22704
rect 2866 22692 2872 22704
rect 2827 22664 2872 22692
rect 2866 22652 2872 22664
rect 2924 22652 2930 22704
rect 2958 22652 2964 22704
rect 3016 22692 3022 22704
rect 3513 22695 3571 22701
rect 3016 22664 3061 22692
rect 3016 22652 3022 22664
rect 3513 22661 3525 22695
rect 3559 22692 3571 22695
rect 6454 22692 6460 22704
rect 3559 22664 6460 22692
rect 3559 22661 3571 22664
rect 3513 22655 3571 22661
rect 6454 22652 6460 22664
rect 6512 22652 6518 22704
rect 7466 22692 7472 22704
rect 7427 22664 7472 22692
rect 7466 22652 7472 22664
rect 7524 22652 7530 22704
rect 7576 22701 7604 22732
rect 12066 22720 12072 22772
rect 12124 22760 12130 22772
rect 12124 22732 12940 22760
rect 12124 22720 12130 22732
rect 7561 22695 7619 22701
rect 7561 22661 7573 22695
rect 7607 22661 7619 22695
rect 7561 22655 7619 22661
rect 8478 22652 8484 22704
rect 8536 22692 8542 22704
rect 9033 22695 9091 22701
rect 9033 22692 9045 22695
rect 8536 22664 9045 22692
rect 8536 22652 8542 22664
rect 9033 22661 9045 22664
rect 9079 22661 9091 22695
rect 9033 22655 9091 22661
rect 9674 22652 9680 22704
rect 9732 22692 9738 22704
rect 10137 22695 10195 22701
rect 10137 22692 10149 22695
rect 9732 22664 10149 22692
rect 9732 22652 9738 22664
rect 10137 22661 10149 22664
rect 10183 22661 10195 22695
rect 10137 22655 10195 22661
rect 10229 22695 10287 22701
rect 10229 22661 10241 22695
rect 10275 22692 10287 22695
rect 11054 22692 11060 22704
rect 10275 22664 11060 22692
rect 10275 22661 10287 22664
rect 10229 22655 10287 22661
rect 11054 22652 11060 22664
rect 11112 22652 11118 22704
rect 11790 22652 11796 22704
rect 11848 22692 11854 22704
rect 12912 22701 12940 22732
rect 14642 22720 14648 22772
rect 14700 22760 14706 22772
rect 14700 22732 22094 22760
rect 14700 22720 14706 22732
rect 12345 22695 12403 22701
rect 12345 22692 12357 22695
rect 11848 22664 12357 22692
rect 11848 22652 11854 22664
rect 12345 22661 12357 22664
rect 12391 22661 12403 22695
rect 12345 22655 12403 22661
rect 12897 22695 12955 22701
rect 12897 22661 12909 22695
rect 12943 22661 12955 22695
rect 12897 22655 12955 22661
rect 17957 22695 18015 22701
rect 17957 22661 17969 22695
rect 18003 22692 18015 22695
rect 18693 22695 18751 22701
rect 18693 22692 18705 22695
rect 18003 22664 18705 22692
rect 18003 22661 18015 22664
rect 17957 22655 18015 22661
rect 18693 22661 18705 22664
rect 18739 22661 18751 22695
rect 18693 22655 18751 22661
rect 21177 22695 21235 22701
rect 21177 22661 21189 22695
rect 21223 22692 21235 22695
rect 21450 22692 21456 22704
rect 21223 22664 21456 22692
rect 21223 22661 21235 22664
rect 21177 22655 21235 22661
rect 21450 22652 21456 22664
rect 21508 22652 21514 22704
rect 22066 22692 22094 22732
rect 37826 22720 37832 22772
rect 37884 22760 37890 22772
rect 38010 22760 38016 22772
rect 37884 22732 38016 22760
rect 37884 22720 37890 22732
rect 38010 22720 38016 22732
rect 38068 22720 38074 22772
rect 22189 22695 22247 22701
rect 22189 22692 22201 22695
rect 22066 22664 22201 22692
rect 22189 22661 22201 22664
rect 22235 22661 22247 22695
rect 22189 22655 22247 22661
rect 4525 22627 4583 22633
rect 4525 22593 4537 22627
rect 4571 22593 4583 22627
rect 4525 22587 4583 22593
rect 1673 22559 1731 22565
rect 1673 22525 1685 22559
rect 1719 22556 1731 22559
rect 3602 22556 3608 22568
rect 1719 22528 3608 22556
rect 1719 22525 1731 22528
rect 1673 22519 1731 22525
rect 3602 22516 3608 22528
rect 3660 22516 3666 22568
rect 2222 22488 2228 22500
rect 2183 22460 2228 22488
rect 2222 22448 2228 22460
rect 2280 22448 2286 22500
rect 4540 22488 4568 22587
rect 5074 22584 5080 22636
rect 5132 22624 5138 22636
rect 5169 22627 5227 22633
rect 5169 22624 5181 22627
rect 5132 22596 5181 22624
rect 5132 22584 5138 22596
rect 5169 22593 5181 22596
rect 5215 22593 5227 22627
rect 5169 22587 5227 22593
rect 5813 22627 5871 22633
rect 5813 22593 5825 22627
rect 5859 22593 5871 22627
rect 6730 22624 6736 22636
rect 6691 22596 6736 22624
rect 5813 22587 5871 22593
rect 5828 22556 5856 22587
rect 6730 22584 6736 22596
rect 6788 22584 6794 22636
rect 13262 22584 13268 22636
rect 13320 22624 13326 22636
rect 13725 22627 13783 22633
rect 13725 22624 13737 22627
rect 13320 22596 13737 22624
rect 13320 22584 13326 22596
rect 13725 22593 13737 22596
rect 13771 22593 13783 22627
rect 13725 22587 13783 22593
rect 16022 22584 16028 22636
rect 16080 22624 16086 22636
rect 17865 22627 17923 22633
rect 17865 22624 17877 22627
rect 16080 22596 17877 22624
rect 16080 22584 16086 22596
rect 17865 22593 17877 22596
rect 17911 22593 17923 22627
rect 17865 22587 17923 22593
rect 23661 22627 23719 22633
rect 23661 22593 23673 22627
rect 23707 22593 23719 22627
rect 23661 22587 23719 22593
rect 7742 22556 7748 22568
rect 5828 22528 7748 22556
rect 7742 22516 7748 22528
rect 7800 22516 7806 22568
rect 8481 22559 8539 22565
rect 8481 22525 8493 22559
rect 8527 22556 8539 22559
rect 8846 22556 8852 22568
rect 8527 22528 8852 22556
rect 8527 22525 8539 22528
rect 8481 22519 8539 22525
rect 8846 22516 8852 22528
rect 8904 22516 8910 22568
rect 10318 22516 10324 22568
rect 10376 22556 10382 22568
rect 10413 22559 10471 22565
rect 10413 22556 10425 22559
rect 10376 22528 10425 22556
rect 10376 22516 10382 22528
rect 10413 22525 10425 22528
rect 10459 22525 10471 22559
rect 10413 22519 10471 22525
rect 6270 22488 6276 22500
rect 4540 22460 6276 22488
rect 6270 22448 6276 22460
rect 6328 22448 6334 22500
rect 6454 22448 6460 22500
rect 6512 22488 6518 22500
rect 9582 22488 9588 22500
rect 6512 22460 9588 22488
rect 6512 22448 6518 22460
rect 9582 22448 9588 22460
rect 9640 22448 9646 22500
rect 10428 22488 10456 22519
rect 12066 22516 12072 22568
rect 12124 22556 12130 22568
rect 12250 22556 12256 22568
rect 12124 22528 12256 22556
rect 12124 22516 12130 22528
rect 12250 22516 12256 22528
rect 12308 22516 12314 22568
rect 12406 22528 17264 22556
rect 12406 22488 12434 22528
rect 17236 22488 17264 22528
rect 17310 22516 17316 22568
rect 17368 22556 17374 22568
rect 18601 22559 18659 22565
rect 18601 22556 18613 22559
rect 17368 22528 18613 22556
rect 17368 22516 17374 22528
rect 18601 22525 18613 22528
rect 18647 22525 18659 22559
rect 18874 22556 18880 22568
rect 18835 22528 18880 22556
rect 18601 22519 18659 22525
rect 18874 22516 18880 22528
rect 18932 22556 18938 22568
rect 19150 22556 19156 22568
rect 18932 22528 19156 22556
rect 18932 22516 18938 22528
rect 19150 22516 19156 22528
rect 19208 22516 19214 22568
rect 22097 22559 22155 22565
rect 22097 22525 22109 22559
rect 22143 22556 22155 22559
rect 22186 22556 22192 22568
rect 22143 22528 22192 22556
rect 22143 22525 22155 22528
rect 22097 22519 22155 22525
rect 22186 22516 22192 22528
rect 22244 22516 22250 22568
rect 22370 22556 22376 22568
rect 22331 22528 22376 22556
rect 22370 22516 22376 22528
rect 22428 22516 22434 22568
rect 23290 22516 23296 22568
rect 23348 22556 23354 22568
rect 23676 22556 23704 22587
rect 23842 22584 23848 22636
rect 23900 22624 23906 22636
rect 24581 22627 24639 22633
rect 24581 22624 24593 22627
rect 23900 22596 24593 22624
rect 23900 22584 23906 22596
rect 24581 22593 24593 22596
rect 24627 22593 24639 22627
rect 24581 22587 24639 22593
rect 37826 22584 37832 22636
rect 37884 22624 37890 22636
rect 38013 22627 38071 22633
rect 38013 22624 38025 22627
rect 37884 22596 38025 22624
rect 37884 22584 37890 22596
rect 38013 22593 38025 22596
rect 38059 22593 38071 22627
rect 38013 22587 38071 22593
rect 37918 22556 37924 22568
rect 23348 22528 37924 22556
rect 23348 22516 23354 22528
rect 37918 22516 37924 22528
rect 37976 22516 37982 22568
rect 18506 22488 18512 22500
rect 10428 22460 12434 22488
rect 13648 22460 13952 22488
rect 17236 22460 18512 22488
rect 4617 22423 4675 22429
rect 4617 22389 4629 22423
rect 4663 22420 4675 22423
rect 5166 22420 5172 22432
rect 4663 22392 5172 22420
rect 4663 22389 4675 22392
rect 4617 22383 4675 22389
rect 5166 22380 5172 22392
rect 5224 22380 5230 22432
rect 5261 22423 5319 22429
rect 5261 22389 5273 22423
rect 5307 22420 5319 22423
rect 5810 22420 5816 22432
rect 5307 22392 5816 22420
rect 5307 22389 5319 22392
rect 5261 22383 5319 22389
rect 5810 22380 5816 22392
rect 5868 22380 5874 22432
rect 5905 22423 5963 22429
rect 5905 22389 5917 22423
rect 5951 22420 5963 22423
rect 6638 22420 6644 22432
rect 5951 22392 6644 22420
rect 5951 22389 5963 22392
rect 5905 22383 5963 22389
rect 6638 22380 6644 22392
rect 6696 22380 6702 22432
rect 9125 22423 9183 22429
rect 9125 22389 9137 22423
rect 9171 22420 9183 22423
rect 13648 22420 13676 22460
rect 13814 22420 13820 22432
rect 9171 22392 13676 22420
rect 13775 22392 13820 22420
rect 9171 22389 9183 22392
rect 9125 22383 9183 22389
rect 13814 22380 13820 22392
rect 13872 22380 13878 22432
rect 13924 22420 13952 22460
rect 18506 22448 18512 22460
rect 18564 22448 18570 22500
rect 21358 22488 21364 22500
rect 21319 22460 21364 22488
rect 21358 22448 21364 22460
rect 21416 22448 21422 22500
rect 34790 22488 34796 22500
rect 22066 22460 34796 22488
rect 22066 22420 22094 22460
rect 34790 22448 34796 22460
rect 34848 22448 34854 22500
rect 38194 22488 38200 22500
rect 38155 22460 38200 22488
rect 38194 22448 38200 22460
rect 38252 22448 38258 22500
rect 13924 22392 22094 22420
rect 22186 22380 22192 22432
rect 22244 22420 22250 22432
rect 23198 22420 23204 22432
rect 22244 22392 23204 22420
rect 22244 22380 22250 22392
rect 23198 22380 23204 22392
rect 23256 22380 23262 22432
rect 23750 22420 23756 22432
rect 23711 22392 23756 22420
rect 23750 22380 23756 22392
rect 23808 22380 23814 22432
rect 24673 22423 24731 22429
rect 24673 22389 24685 22423
rect 24719 22420 24731 22423
rect 24762 22420 24768 22432
rect 24719 22392 24768 22420
rect 24719 22389 24731 22392
rect 24673 22383 24731 22389
rect 24762 22380 24768 22392
rect 24820 22380 24826 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 3602 22176 3608 22228
rect 3660 22216 3666 22228
rect 16114 22216 16120 22228
rect 3660 22188 16120 22216
rect 3660 22176 3666 22188
rect 16114 22176 16120 22188
rect 16172 22176 16178 22228
rect 17494 22176 17500 22228
rect 17552 22216 17558 22228
rect 17862 22216 17868 22228
rect 17552 22188 17868 22216
rect 17552 22176 17558 22188
rect 17862 22176 17868 22188
rect 17920 22176 17926 22228
rect 7466 22108 7472 22160
rect 7524 22148 7530 22160
rect 8386 22148 8392 22160
rect 7524 22120 8392 22148
rect 7524 22108 7530 22120
rect 8386 22108 8392 22120
rect 8444 22108 8450 22160
rect 11054 22148 11060 22160
rect 9508 22120 11060 22148
rect 1857 22083 1915 22089
rect 1857 22049 1869 22083
rect 1903 22080 1915 22083
rect 2038 22080 2044 22092
rect 1903 22052 2044 22080
rect 1903 22049 1915 22052
rect 1857 22043 1915 22049
rect 2038 22040 2044 22052
rect 2096 22040 2102 22092
rect 2406 22080 2412 22092
rect 2367 22052 2412 22080
rect 2406 22040 2412 22052
rect 2464 22040 2470 22092
rect 4614 22080 4620 22092
rect 4172 22052 4620 22080
rect 4172 22024 4200 22052
rect 4614 22040 4620 22052
rect 4672 22040 4678 22092
rect 4982 22080 4988 22092
rect 4943 22052 4988 22080
rect 4982 22040 4988 22052
rect 5040 22040 5046 22092
rect 5810 22040 5816 22092
rect 5868 22080 5874 22092
rect 6454 22080 6460 22092
rect 5868 22052 6460 22080
rect 5868 22040 5874 22052
rect 6454 22040 6460 22052
rect 6512 22080 6518 22092
rect 6733 22083 6791 22089
rect 6733 22080 6745 22083
rect 6512 22052 6745 22080
rect 6512 22040 6518 22052
rect 6733 22049 6745 22052
rect 6779 22049 6791 22083
rect 6733 22043 6791 22049
rect 7377 22083 7435 22089
rect 7377 22049 7389 22083
rect 7423 22080 7435 22083
rect 7742 22080 7748 22092
rect 7423 22052 7748 22080
rect 7423 22049 7435 22052
rect 7377 22043 7435 22049
rect 7742 22040 7748 22052
rect 7800 22080 7806 22092
rect 9508 22080 9536 22120
rect 11054 22108 11060 22120
rect 11112 22108 11118 22160
rect 12066 22108 12072 22160
rect 12124 22148 12130 22160
rect 12124 22120 12204 22148
rect 12124 22108 12130 22120
rect 7800 22052 9536 22080
rect 7800 22040 7806 22052
rect 9582 22040 9588 22092
rect 9640 22080 9646 22092
rect 9677 22083 9735 22089
rect 9677 22080 9689 22083
rect 9640 22052 9689 22080
rect 9640 22040 9646 22052
rect 9677 22049 9689 22052
rect 9723 22049 9735 22083
rect 9677 22043 9735 22049
rect 1765 22015 1823 22021
rect 1765 21981 1777 22015
rect 1811 22012 1823 22015
rect 1811 21984 2268 22012
rect 1811 21981 1823 21984
rect 1765 21975 1823 21981
rect 2240 21876 2268 21984
rect 4154 21972 4160 22024
rect 4212 21972 4218 22024
rect 4249 22015 4307 22021
rect 4249 21981 4261 22015
rect 4295 22012 4307 22015
rect 4798 22012 4804 22024
rect 4295 21984 4804 22012
rect 4295 21981 4307 21984
rect 4249 21975 4307 21981
rect 4798 21972 4804 21984
rect 4856 21972 4862 22024
rect 8386 22012 8392 22024
rect 8347 21984 8392 22012
rect 8386 21972 8392 21984
rect 8444 21972 8450 22024
rect 12066 22012 12072 22024
rect 11624 21984 12072 22012
rect 2498 21904 2504 21956
rect 2556 21944 2562 21956
rect 3053 21947 3111 21953
rect 2556 21916 2601 21944
rect 2556 21904 2562 21916
rect 3053 21913 3065 21947
rect 3099 21944 3111 21947
rect 3602 21944 3608 21956
rect 3099 21916 3608 21944
rect 3099 21913 3111 21916
rect 3053 21907 3111 21913
rect 3602 21904 3608 21916
rect 3660 21904 3666 21956
rect 5077 21947 5135 21953
rect 5077 21913 5089 21947
rect 5123 21913 5135 21947
rect 5077 21907 5135 21913
rect 5629 21947 5687 21953
rect 5629 21913 5641 21947
rect 5675 21944 5687 21947
rect 5810 21944 5816 21956
rect 5675 21916 5816 21944
rect 5675 21913 5687 21916
rect 5629 21907 5687 21913
rect 4246 21876 4252 21888
rect 2240 21848 4252 21876
rect 4246 21836 4252 21848
rect 4304 21836 4310 21888
rect 4338 21836 4344 21888
rect 4396 21876 4402 21888
rect 5092 21876 5120 21907
rect 5810 21904 5816 21916
rect 5868 21904 5874 21956
rect 6825 21947 6883 21953
rect 6825 21913 6837 21947
rect 6871 21913 6883 21947
rect 9398 21944 9404 21956
rect 9359 21916 9404 21944
rect 6825 21907 6883 21913
rect 5718 21876 5724 21888
rect 4396 21848 4441 21876
rect 5092 21848 5724 21876
rect 4396 21836 4402 21848
rect 5718 21836 5724 21848
rect 5776 21836 5782 21888
rect 6840 21876 6868 21907
rect 9398 21904 9404 21916
rect 9456 21904 9462 21956
rect 9490 21904 9496 21956
rect 9548 21944 9554 21956
rect 10689 21947 10747 21953
rect 9548 21916 9593 21944
rect 9548 21904 9554 21916
rect 10689 21913 10701 21947
rect 10735 21913 10747 21947
rect 10689 21907 10747 21913
rect 10781 21947 10839 21953
rect 10781 21913 10793 21947
rect 10827 21944 10839 21947
rect 11146 21944 11152 21956
rect 10827 21916 11152 21944
rect 10827 21913 10839 21916
rect 10781 21907 10839 21913
rect 7926 21876 7932 21888
rect 6840 21848 7932 21876
rect 7926 21836 7932 21848
rect 7984 21836 7990 21888
rect 8481 21879 8539 21885
rect 8481 21845 8493 21879
rect 8527 21876 8539 21879
rect 9950 21876 9956 21888
rect 8527 21848 9956 21876
rect 8527 21845 8539 21848
rect 8481 21839 8539 21845
rect 9950 21836 9956 21848
rect 10008 21836 10014 21888
rect 10704 21876 10732 21907
rect 11146 21904 11152 21916
rect 11204 21904 11210 21956
rect 11330 21904 11336 21956
rect 11388 21944 11394 21956
rect 11624 21944 11652 21984
rect 12066 21972 12072 21984
rect 12124 21972 12130 22024
rect 11388 21916 11652 21944
rect 11701 21947 11759 21953
rect 11388 21904 11394 21916
rect 11701 21913 11713 21947
rect 11747 21944 11759 21947
rect 11882 21944 11888 21956
rect 11747 21916 11888 21944
rect 11747 21913 11759 21916
rect 11701 21907 11759 21913
rect 11882 21904 11888 21916
rect 11940 21904 11946 21956
rect 12176 21944 12204 22120
rect 17954 22108 17960 22160
rect 18012 22148 18018 22160
rect 22922 22148 22928 22160
rect 18012 22120 22928 22148
rect 18012 22108 18018 22120
rect 22922 22108 22928 22120
rect 22980 22108 22986 22160
rect 14642 22080 14648 22092
rect 14603 22052 14648 22080
rect 14642 22040 14648 22052
rect 14700 22040 14706 22092
rect 13188 21984 13676 22012
rect 12345 21947 12403 21953
rect 12345 21944 12357 21947
rect 12176 21916 12357 21944
rect 12345 21913 12357 21916
rect 12391 21913 12403 21947
rect 12345 21907 12403 21913
rect 12434 21904 12440 21956
rect 12492 21944 12498 21956
rect 12492 21916 12537 21944
rect 12492 21904 12498 21916
rect 12710 21904 12716 21956
rect 12768 21944 12774 21956
rect 13188 21944 13216 21984
rect 12768 21916 13216 21944
rect 13357 21947 13415 21953
rect 12768 21904 12774 21916
rect 13357 21913 13369 21947
rect 13403 21944 13415 21947
rect 13538 21944 13544 21956
rect 13403 21916 13544 21944
rect 13403 21913 13415 21916
rect 13357 21907 13415 21913
rect 13372 21876 13400 21907
rect 13538 21904 13544 21916
rect 13596 21904 13602 21956
rect 10704 21848 13400 21876
rect 13648 21876 13676 21984
rect 14090 21972 14096 22024
rect 14148 22012 14154 22024
rect 14553 22015 14611 22021
rect 14553 22012 14565 22015
rect 14148 21984 14565 22012
rect 14148 21972 14154 21984
rect 14553 21981 14565 21984
rect 14599 21981 14611 22015
rect 15197 22015 15255 22021
rect 15197 22012 15209 22015
rect 14553 21975 14611 21981
rect 14660 21984 15209 22012
rect 13722 21904 13728 21956
rect 13780 21944 13786 21956
rect 14660 21944 14688 21984
rect 15197 21981 15209 21984
rect 15243 21981 15255 22015
rect 15197 21975 15255 21981
rect 22097 22015 22155 22021
rect 22097 21981 22109 22015
rect 22143 22012 22155 22015
rect 23014 22012 23020 22024
rect 22143 21984 23020 22012
rect 22143 21981 22155 21984
rect 22097 21975 22155 21981
rect 23014 21972 23020 21984
rect 23072 21972 23078 22024
rect 23201 22015 23259 22021
rect 23201 21981 23213 22015
rect 23247 22012 23259 22015
rect 23290 22012 23296 22024
rect 23247 21984 23296 22012
rect 23247 21981 23259 21984
rect 23201 21975 23259 21981
rect 23290 21972 23296 21984
rect 23348 21972 23354 22024
rect 38010 22012 38016 22024
rect 37971 21984 38016 22012
rect 38010 21972 38016 21984
rect 38068 21972 38074 22024
rect 18138 21944 18144 21956
rect 13780 21916 14688 21944
rect 14752 21916 18144 21944
rect 13780 21904 13786 21916
rect 14752 21876 14780 21916
rect 18138 21904 18144 21916
rect 18196 21904 18202 21956
rect 15286 21876 15292 21888
rect 13648 21848 14780 21876
rect 15247 21848 15292 21876
rect 15286 21836 15292 21848
rect 15344 21836 15350 21888
rect 21913 21879 21971 21885
rect 21913 21845 21925 21879
rect 21959 21876 21971 21879
rect 22186 21876 22192 21888
rect 21959 21848 22192 21876
rect 21959 21845 21971 21848
rect 21913 21839 21971 21845
rect 22186 21836 22192 21848
rect 22244 21836 22250 21888
rect 23290 21876 23296 21888
rect 23251 21848 23296 21876
rect 23290 21836 23296 21848
rect 23348 21836 23354 21888
rect 37829 21879 37887 21885
rect 37829 21845 37841 21879
rect 37875 21876 37887 21879
rect 37918 21876 37924 21888
rect 37875 21848 37924 21876
rect 37875 21845 37887 21848
rect 37829 21839 37887 21845
rect 37918 21836 37924 21848
rect 37976 21836 37982 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 2498 21632 2504 21684
rect 2556 21672 2562 21684
rect 5905 21675 5963 21681
rect 2556 21644 4660 21672
rect 2556 21632 2562 21644
rect 1857 21607 1915 21613
rect 1857 21573 1869 21607
rect 1903 21604 1915 21607
rect 1946 21604 1952 21616
rect 1903 21576 1952 21604
rect 1903 21573 1915 21576
rect 1857 21567 1915 21573
rect 1946 21564 1952 21576
rect 2004 21564 2010 21616
rect 2038 21564 2044 21616
rect 2096 21604 2102 21616
rect 3329 21607 3387 21613
rect 3329 21604 3341 21607
rect 2096 21576 3341 21604
rect 2096 21564 2102 21576
rect 3329 21573 3341 21576
rect 3375 21573 3387 21607
rect 3329 21567 3387 21573
rect 3421 21607 3479 21613
rect 3421 21573 3433 21607
rect 3467 21604 3479 21607
rect 4154 21604 4160 21616
rect 3467 21576 4160 21604
rect 3467 21573 3479 21576
rect 3421 21567 3479 21573
rect 4154 21564 4160 21576
rect 4212 21564 4218 21616
rect 4632 21613 4660 21644
rect 5905 21641 5917 21675
rect 5951 21672 5963 21675
rect 11885 21675 11943 21681
rect 5951 21644 8800 21672
rect 5951 21641 5963 21644
rect 5905 21635 5963 21641
rect 4617 21607 4675 21613
rect 4617 21573 4629 21607
rect 4663 21573 4675 21607
rect 6730 21604 6736 21616
rect 6691 21576 6736 21604
rect 4617 21567 4675 21573
rect 6730 21564 6736 21576
rect 6788 21564 6794 21616
rect 8772 21613 8800 21644
rect 11885 21641 11897 21675
rect 11931 21672 11943 21675
rect 12434 21672 12440 21684
rect 11931 21644 12440 21672
rect 11931 21641 11943 21644
rect 11885 21635 11943 21641
rect 12434 21632 12440 21644
rect 12492 21632 12498 21684
rect 13170 21632 13176 21684
rect 13228 21672 13234 21684
rect 13446 21672 13452 21684
rect 13228 21644 13452 21672
rect 13228 21632 13234 21644
rect 13446 21632 13452 21644
rect 13504 21632 13510 21684
rect 13538 21632 13544 21684
rect 13596 21672 13602 21684
rect 16298 21672 16304 21684
rect 13596 21644 16304 21672
rect 13596 21632 13602 21644
rect 16298 21632 16304 21644
rect 16356 21632 16362 21684
rect 23198 21632 23204 21684
rect 23256 21672 23262 21684
rect 28813 21675 28871 21681
rect 28813 21672 28825 21675
rect 23256 21644 28825 21672
rect 23256 21632 23262 21644
rect 28813 21641 28825 21644
rect 28859 21641 28871 21675
rect 28813 21635 28871 21641
rect 8750 21607 8808 21613
rect 8750 21573 8762 21607
rect 8796 21573 8808 21607
rect 8750 21567 8808 21573
rect 8938 21564 8944 21616
rect 8996 21604 9002 21616
rect 9674 21604 9680 21616
rect 8996 21576 9680 21604
rect 8996 21564 9002 21576
rect 9674 21564 9680 21576
rect 9732 21564 9738 21616
rect 9950 21564 9956 21616
rect 10008 21604 10014 21616
rect 11057 21607 11115 21613
rect 10008 21576 10053 21604
rect 10008 21564 10014 21576
rect 11057 21573 11069 21607
rect 11103 21604 11115 21607
rect 14645 21607 14703 21613
rect 14645 21604 14657 21607
rect 11103 21576 14657 21604
rect 11103 21573 11115 21576
rect 11057 21567 11115 21573
rect 14645 21573 14657 21576
rect 14691 21573 14703 21607
rect 14645 21567 14703 21573
rect 15010 21564 15016 21616
rect 15068 21604 15074 21616
rect 15197 21607 15255 21613
rect 15197 21604 15209 21607
rect 15068 21576 15209 21604
rect 15068 21564 15074 21576
rect 15197 21573 15209 21576
rect 15243 21573 15255 21607
rect 15197 21567 15255 21573
rect 15654 21564 15660 21616
rect 15712 21604 15718 21616
rect 15930 21604 15936 21616
rect 15712 21576 15936 21604
rect 15712 21564 15718 21576
rect 15930 21564 15936 21576
rect 15988 21564 15994 21616
rect 17494 21604 17500 21616
rect 17455 21576 17500 21604
rect 17494 21564 17500 21576
rect 17552 21564 17558 21616
rect 17586 21564 17592 21616
rect 17644 21604 17650 21616
rect 17644 21576 17689 21604
rect 17644 21564 17650 21576
rect 21542 21564 21548 21616
rect 21600 21604 21606 21616
rect 22189 21607 22247 21613
rect 22189 21604 22201 21607
rect 21600 21576 22201 21604
rect 21600 21564 21606 21576
rect 22189 21573 22201 21576
rect 22235 21573 22247 21607
rect 23106 21604 23112 21616
rect 23067 21576 23112 21604
rect 22189 21567 22247 21573
rect 23106 21564 23112 21576
rect 23164 21564 23170 21616
rect 37366 21604 37372 21616
rect 28736 21576 37372 21604
rect 5813 21539 5871 21545
rect 5813 21505 5825 21539
rect 5859 21536 5871 21539
rect 6362 21536 6368 21548
rect 5859 21508 6368 21536
rect 5859 21505 5871 21508
rect 5813 21499 5871 21505
rect 6362 21496 6368 21508
rect 6420 21496 6426 21548
rect 7576 21508 8524 21536
rect 1765 21471 1823 21477
rect 1765 21437 1777 21471
rect 1811 21437 1823 21471
rect 1765 21431 1823 21437
rect 1780 21400 1808 21431
rect 2222 21428 2228 21480
rect 2280 21468 2286 21480
rect 2406 21468 2412 21480
rect 2280 21440 2412 21468
rect 2280 21428 2286 21440
rect 2406 21428 2412 21440
rect 2464 21428 2470 21480
rect 3602 21468 3608 21480
rect 3563 21440 3608 21468
rect 3602 21428 3608 21440
rect 3660 21428 3666 21480
rect 4525 21471 4583 21477
rect 4525 21468 4537 21471
rect 3804 21440 4537 21468
rect 1780 21372 2774 21400
rect 2746 21332 2774 21372
rect 2866 21360 2872 21412
rect 2924 21400 2930 21412
rect 3804 21400 3832 21440
rect 4525 21437 4537 21440
rect 4571 21437 4583 21471
rect 4525 21431 4583 21437
rect 4798 21428 4804 21480
rect 4856 21468 4862 21480
rect 4856 21440 6408 21468
rect 4856 21428 4862 21440
rect 2924 21372 3832 21400
rect 2924 21360 2930 21372
rect 4246 21360 4252 21412
rect 4304 21400 4310 21412
rect 5074 21400 5080 21412
rect 4304 21372 5080 21400
rect 4304 21360 4310 21372
rect 5074 21360 5080 21372
rect 5132 21360 5138 21412
rect 6380 21400 6408 21440
rect 6454 21428 6460 21480
rect 6512 21468 6518 21480
rect 6641 21471 6699 21477
rect 6641 21468 6653 21471
rect 6512 21440 6653 21468
rect 6512 21428 6518 21440
rect 6641 21437 6653 21440
rect 6687 21437 6699 21471
rect 6641 21431 6699 21437
rect 6822 21428 6828 21480
rect 6880 21468 6886 21480
rect 7576 21468 7604 21508
rect 6880 21440 7604 21468
rect 7653 21471 7711 21477
rect 6880 21428 6886 21440
rect 7653 21437 7665 21471
rect 7699 21468 7711 21471
rect 8110 21468 8116 21480
rect 7699 21440 8116 21468
rect 7699 21437 7711 21440
rect 7653 21431 7711 21437
rect 8110 21428 8116 21440
rect 8168 21428 8174 21480
rect 8202 21400 8208 21412
rect 6380 21372 8208 21400
rect 8202 21360 8208 21372
rect 8260 21360 8266 21412
rect 8496 21400 8524 21508
rect 10962 21496 10968 21548
rect 11020 21536 11026 21548
rect 11020 21508 11065 21536
rect 11020 21496 11026 21508
rect 11330 21496 11336 21548
rect 11388 21536 11394 21548
rect 11793 21539 11851 21545
rect 11793 21536 11805 21539
rect 11388 21508 11805 21536
rect 11388 21496 11394 21508
rect 11793 21505 11805 21508
rect 11839 21505 11851 21539
rect 11793 21499 11851 21505
rect 12434 21496 12440 21548
rect 12492 21536 12498 21548
rect 12492 21508 12537 21536
rect 12492 21496 12498 21508
rect 13170 21496 13176 21548
rect 13228 21536 13234 21548
rect 13265 21539 13323 21545
rect 13265 21536 13277 21539
rect 13228 21508 13277 21536
rect 13228 21496 13234 21508
rect 13265 21505 13277 21508
rect 13311 21505 13323 21539
rect 13722 21536 13728 21548
rect 13683 21508 13728 21536
rect 13265 21499 13323 21505
rect 13722 21496 13728 21508
rect 13780 21496 13786 21548
rect 15838 21536 15844 21548
rect 15799 21508 15844 21536
rect 15838 21496 15844 21508
rect 15896 21496 15902 21548
rect 23014 21496 23020 21548
rect 23072 21536 23078 21548
rect 25317 21539 25375 21545
rect 25317 21536 25329 21539
rect 23072 21508 25329 21536
rect 23072 21496 23078 21508
rect 25317 21505 25329 21508
rect 25363 21536 25375 21539
rect 27062 21536 27068 21548
rect 25363 21508 27068 21536
rect 25363 21505 25375 21508
rect 25317 21499 25375 21505
rect 27062 21496 27068 21508
rect 27120 21496 27126 21548
rect 27982 21536 27988 21548
rect 27943 21508 27988 21536
rect 27982 21496 27988 21508
rect 28040 21496 28046 21548
rect 28736 21545 28764 21576
rect 37366 21564 37372 21576
rect 37424 21564 37430 21616
rect 28721 21539 28779 21545
rect 28721 21505 28733 21539
rect 28767 21505 28779 21539
rect 28721 21499 28779 21505
rect 31386 21496 31392 21548
rect 31444 21536 31450 21548
rect 32493 21539 32551 21545
rect 32493 21536 32505 21539
rect 31444 21508 32505 21536
rect 31444 21496 31450 21508
rect 32493 21505 32505 21508
rect 32539 21505 32551 21539
rect 38013 21539 38071 21545
rect 38013 21536 38025 21539
rect 32493 21499 32551 21505
rect 35866 21508 38025 21536
rect 8665 21471 8723 21477
rect 8665 21437 8677 21471
rect 8711 21456 8723 21471
rect 8846 21468 8852 21480
rect 8772 21456 8852 21468
rect 8711 21440 8852 21456
rect 8711 21437 8800 21440
rect 8665 21431 8800 21437
rect 8680 21428 8800 21431
rect 8846 21428 8852 21440
rect 8904 21428 8910 21480
rect 9861 21471 9919 21477
rect 9861 21437 9873 21471
rect 9907 21468 9919 21471
rect 13630 21468 13636 21480
rect 9907 21456 10824 21468
rect 10980 21456 13636 21468
rect 9907 21440 13636 21456
rect 9907 21437 9919 21440
rect 9861 21431 9919 21437
rect 10796 21428 11008 21440
rect 13630 21428 13636 21440
rect 13688 21428 13694 21480
rect 8938 21400 8944 21412
rect 8496 21372 8944 21400
rect 8938 21360 8944 21372
rect 8996 21360 9002 21412
rect 9217 21403 9275 21409
rect 9217 21369 9229 21403
rect 9263 21369 9275 21403
rect 9217 21363 9275 21369
rect 4798 21332 4804 21344
rect 2746 21304 4804 21332
rect 4798 21292 4804 21304
rect 4856 21292 4862 21344
rect 5810 21292 5816 21344
rect 5868 21332 5874 21344
rect 8754 21332 8760 21344
rect 5868 21304 8760 21332
rect 5868 21292 5874 21304
rect 8754 21292 8760 21304
rect 8812 21292 8818 21344
rect 9232 21332 9260 21363
rect 9582 21360 9588 21412
rect 9640 21400 9646 21412
rect 10413 21403 10471 21409
rect 10413 21400 10425 21403
rect 9640 21372 10425 21400
rect 9640 21360 9646 21372
rect 10413 21369 10425 21372
rect 10459 21369 10471 21403
rect 10413 21363 10471 21369
rect 12250 21360 12256 21412
rect 12308 21400 12314 21412
rect 13740 21400 13768 21496
rect 14553 21471 14611 21477
rect 14553 21437 14565 21471
rect 14599 21468 14611 21471
rect 17310 21468 17316 21480
rect 14599 21440 17316 21468
rect 14599 21437 14611 21440
rect 14553 21431 14611 21437
rect 17310 21428 17316 21440
rect 17368 21428 17374 21480
rect 17678 21428 17684 21480
rect 17736 21468 17742 21480
rect 17957 21471 18015 21477
rect 17957 21468 17969 21471
rect 17736 21440 17969 21468
rect 17736 21428 17742 21440
rect 17957 21437 17969 21440
rect 18003 21437 18015 21471
rect 17957 21431 18015 21437
rect 18046 21428 18052 21480
rect 18104 21468 18110 21480
rect 18874 21468 18880 21480
rect 18104 21440 18880 21468
rect 18104 21428 18110 21440
rect 18874 21428 18880 21440
rect 18932 21428 18938 21480
rect 22097 21471 22155 21477
rect 22097 21437 22109 21471
rect 22143 21468 22155 21471
rect 23750 21468 23756 21480
rect 22143 21440 23756 21468
rect 22143 21437 22155 21440
rect 22097 21431 22155 21437
rect 23750 21428 23756 21440
rect 23808 21468 23814 21480
rect 24029 21471 24087 21477
rect 24029 21468 24041 21471
rect 23808 21440 24041 21468
rect 23808 21428 23814 21440
rect 24029 21437 24041 21440
rect 24075 21437 24087 21471
rect 24029 21431 24087 21437
rect 24213 21471 24271 21477
rect 24213 21437 24225 21471
rect 24259 21468 24271 21471
rect 25409 21471 25467 21477
rect 25409 21468 25421 21471
rect 24259 21440 25421 21468
rect 24259 21437 24271 21440
rect 24213 21431 24271 21437
rect 25409 21437 25421 21440
rect 25455 21437 25467 21471
rect 25409 21431 25467 21437
rect 12308 21372 13768 21400
rect 12308 21360 12314 21372
rect 15010 21360 15016 21412
rect 15068 21400 15074 21412
rect 20162 21400 20168 21412
rect 15068 21372 20168 21400
rect 15068 21360 15074 21372
rect 20162 21360 20168 21372
rect 20220 21360 20226 21412
rect 32309 21403 32367 21409
rect 32309 21369 32321 21403
rect 32355 21400 32367 21403
rect 35866 21400 35894 21508
rect 38013 21505 38025 21508
rect 38059 21505 38071 21539
rect 38013 21499 38071 21505
rect 32355 21372 35894 21400
rect 32355 21369 32367 21372
rect 32309 21363 32367 21369
rect 11698 21332 11704 21344
rect 9232 21304 11704 21332
rect 11698 21292 11704 21304
rect 11756 21292 11762 21344
rect 12526 21332 12532 21344
rect 12487 21304 12532 21332
rect 12526 21292 12532 21304
rect 12584 21292 12590 21344
rect 13081 21335 13139 21341
rect 13081 21301 13093 21335
rect 13127 21332 13139 21335
rect 13722 21332 13728 21344
rect 13127 21304 13728 21332
rect 13127 21301 13139 21304
rect 13081 21295 13139 21301
rect 13722 21292 13728 21304
rect 13780 21292 13786 21344
rect 13817 21335 13875 21341
rect 13817 21301 13829 21335
rect 13863 21332 13875 21335
rect 13906 21332 13912 21344
rect 13863 21304 13912 21332
rect 13863 21301 13875 21304
rect 13817 21295 13875 21301
rect 13906 21292 13912 21304
rect 13964 21292 13970 21344
rect 13998 21292 14004 21344
rect 14056 21332 14062 21344
rect 15657 21335 15715 21341
rect 15657 21332 15669 21335
rect 14056 21304 15669 21332
rect 14056 21292 14062 21304
rect 15657 21301 15669 21304
rect 15703 21301 15715 21335
rect 15657 21295 15715 21301
rect 16298 21292 16304 21344
rect 16356 21332 16362 21344
rect 18690 21332 18696 21344
rect 16356 21304 18696 21332
rect 16356 21292 16362 21304
rect 18690 21292 18696 21304
rect 18748 21332 18754 21344
rect 23106 21332 23112 21344
rect 18748 21304 23112 21332
rect 18748 21292 18754 21304
rect 23106 21292 23112 21304
rect 23164 21292 23170 21344
rect 24486 21332 24492 21344
rect 24447 21304 24492 21332
rect 24486 21292 24492 21304
rect 24544 21292 24550 21344
rect 27798 21332 27804 21344
rect 27759 21304 27804 21332
rect 27798 21292 27804 21304
rect 27856 21292 27862 21344
rect 38194 21332 38200 21344
rect 38155 21304 38200 21332
rect 38194 21292 38200 21304
rect 38252 21292 38258 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 1762 21128 1768 21140
rect 1723 21100 1768 21128
rect 1762 21088 1768 21100
rect 1820 21088 1826 21140
rect 3878 21128 3884 21140
rect 2240 21100 3884 21128
rect 1581 20927 1639 20933
rect 1581 20893 1593 20927
rect 1627 20924 1639 20927
rect 2240 20924 2268 21100
rect 3878 21088 3884 21100
rect 3936 21088 3942 21140
rect 8754 21088 8760 21140
rect 8812 21128 8818 21140
rect 9306 21128 9312 21140
rect 8812 21100 9312 21128
rect 8812 21088 8818 21100
rect 9306 21088 9312 21100
rect 9364 21088 9370 21140
rect 9401 21131 9459 21137
rect 9401 21097 9413 21131
rect 9447 21128 9459 21131
rect 15838 21128 15844 21140
rect 9447 21100 15844 21128
rect 9447 21097 9459 21100
rect 9401 21091 9459 21097
rect 15838 21088 15844 21100
rect 15896 21088 15902 21140
rect 17313 21131 17371 21137
rect 17313 21097 17325 21131
rect 17359 21128 17371 21131
rect 17586 21128 17592 21140
rect 17359 21100 17592 21128
rect 17359 21097 17371 21100
rect 17313 21091 17371 21097
rect 17586 21088 17592 21100
rect 17644 21088 17650 21140
rect 21450 21128 21456 21140
rect 17972 21100 21456 21128
rect 3602 21020 3608 21072
rect 3660 21060 3666 21072
rect 3660 21032 5580 21060
rect 3660 21020 3666 21032
rect 2409 20995 2467 21001
rect 2409 20961 2421 20995
rect 2455 20992 2467 20995
rect 3050 20992 3056 21004
rect 2455 20964 3056 20992
rect 2455 20961 2467 20964
rect 2409 20955 2467 20961
rect 3050 20952 3056 20964
rect 3108 20952 3114 21004
rect 4246 20952 4252 21004
rect 4304 20992 4310 21004
rect 4706 20992 4712 21004
rect 4304 20964 4712 20992
rect 4304 20952 4310 20964
rect 4706 20952 4712 20964
rect 4764 20952 4770 21004
rect 5258 20992 5264 21004
rect 5219 20964 5264 20992
rect 5258 20952 5264 20964
rect 5316 20952 5322 21004
rect 5552 21001 5580 21032
rect 5718 21020 5724 21072
rect 5776 21060 5782 21072
rect 6822 21060 6828 21072
rect 5776 21032 6828 21060
rect 5776 21020 5782 21032
rect 6822 21020 6828 21032
rect 6880 21020 6886 21072
rect 7745 21063 7803 21069
rect 7745 21029 7757 21063
rect 7791 21060 7803 21063
rect 13538 21060 13544 21072
rect 7791 21032 13544 21060
rect 7791 21029 7803 21032
rect 7745 21023 7803 21029
rect 13538 21020 13544 21032
rect 13596 21020 13602 21072
rect 13630 21020 13636 21072
rect 13688 21060 13694 21072
rect 13688 21032 14596 21060
rect 13688 21020 13694 21032
rect 5537 20995 5595 21001
rect 5537 20961 5549 20995
rect 5583 20961 5595 20995
rect 7190 20992 7196 21004
rect 7151 20964 7196 20992
rect 5537 20955 5595 20961
rect 7190 20952 7196 20964
rect 7248 20952 7254 21004
rect 9398 20952 9404 21004
rect 9456 20992 9462 21004
rect 9674 20992 9680 21004
rect 9456 20964 9680 20992
rect 9456 20952 9462 20964
rect 9674 20952 9680 20964
rect 9732 20952 9738 21004
rect 10152 21001 10272 21004
rect 10138 20995 10272 21001
rect 10138 20961 10150 20995
rect 10184 20992 10272 20995
rect 10778 20992 10784 21004
rect 10184 20976 10784 20992
rect 10184 20961 10196 20976
rect 10244 20964 10784 20976
rect 10138 20955 10196 20961
rect 10778 20952 10784 20964
rect 10836 20952 10842 21004
rect 11149 20995 11207 21001
rect 11149 20961 11161 20995
rect 11195 20992 11207 20995
rect 12158 20992 12164 21004
rect 11195 20964 12164 20992
rect 11195 20961 11207 20964
rect 11149 20955 11207 20961
rect 12158 20952 12164 20964
rect 12216 20952 12222 21004
rect 12618 20992 12624 21004
rect 12579 20964 12624 20992
rect 12618 20952 12624 20964
rect 12676 20952 12682 21004
rect 13814 20952 13820 21004
rect 13872 20992 13878 21004
rect 14461 20995 14519 21001
rect 14461 20992 14473 20995
rect 13872 20964 14473 20992
rect 13872 20952 13878 20964
rect 14461 20961 14473 20964
rect 14507 20961 14519 20995
rect 14568 20992 14596 21032
rect 15470 21020 15476 21072
rect 15528 21060 15534 21072
rect 16574 21060 16580 21072
rect 15528 21032 16580 21060
rect 15528 21020 15534 21032
rect 16574 21020 16580 21032
rect 16632 21020 16638 21072
rect 17972 20992 18000 21100
rect 21450 21088 21456 21100
rect 21508 21088 21514 21140
rect 31386 21128 31392 21140
rect 31347 21100 31392 21128
rect 31386 21088 31392 21100
rect 31444 21088 31450 21140
rect 37369 21131 37427 21137
rect 37369 21097 37381 21131
rect 37415 21128 37427 21131
rect 38470 21128 38476 21140
rect 37415 21100 38476 21128
rect 37415 21097 37427 21100
rect 37369 21091 37427 21097
rect 38470 21088 38476 21100
rect 38528 21088 38534 21140
rect 23198 21060 23204 21072
rect 19444 21032 23204 21060
rect 19444 21001 19472 21032
rect 23198 21020 23204 21032
rect 23256 21020 23262 21072
rect 14568 20964 16436 20992
rect 14461 20955 14519 20961
rect 1627 20896 2268 20924
rect 6457 20927 6515 20933
rect 1627 20893 1639 20896
rect 1581 20887 1639 20893
rect 6457 20893 6469 20927
rect 6503 20924 6515 20927
rect 6822 20924 6828 20936
rect 6503 20896 6828 20924
rect 6503 20893 6515 20896
rect 6457 20887 6515 20893
rect 6822 20884 6828 20896
rect 6880 20884 6886 20936
rect 8389 20927 8447 20933
rect 8389 20893 8401 20927
rect 8435 20924 8447 20927
rect 9122 20924 9128 20936
rect 8435 20896 9128 20924
rect 8435 20893 8447 20896
rect 8389 20887 8447 20893
rect 9122 20884 9128 20896
rect 9180 20884 9186 20936
rect 9593 20923 9651 20929
rect 13722 20924 13728 20936
rect 9593 20889 9605 20923
rect 9639 20920 9651 20923
rect 9639 20889 9674 20920
rect 13683 20896 13728 20924
rect 9593 20883 9674 20889
rect 13722 20884 13728 20896
rect 13780 20884 13786 20936
rect 14274 20924 14280 20936
rect 14235 20896 14280 20924
rect 14274 20884 14280 20896
rect 14332 20884 14338 20936
rect 14642 20884 14648 20936
rect 14700 20924 14706 20936
rect 14918 20924 14924 20936
rect 14700 20896 14924 20924
rect 14700 20884 14706 20896
rect 14918 20884 14924 20896
rect 14976 20884 14982 20936
rect 15381 20927 15439 20933
rect 15381 20893 15393 20927
rect 15427 20924 15439 20927
rect 15470 20924 15476 20936
rect 15427 20896 15476 20924
rect 15427 20893 15439 20896
rect 15381 20887 15439 20893
rect 15470 20884 15476 20896
rect 15528 20884 15534 20936
rect 2501 20859 2559 20865
rect 2501 20825 2513 20859
rect 2547 20856 2559 20859
rect 2590 20856 2596 20868
rect 2547 20828 2596 20856
rect 2547 20825 2559 20828
rect 2501 20819 2559 20825
rect 2590 20816 2596 20828
rect 2648 20816 2654 20868
rect 3053 20859 3111 20865
rect 3053 20856 3065 20859
rect 2746 20828 3065 20856
rect 2406 20748 2412 20800
rect 2464 20788 2470 20800
rect 2746 20788 2774 20828
rect 3053 20825 3065 20828
rect 3099 20825 3111 20859
rect 4065 20859 4123 20865
rect 4065 20856 4077 20859
rect 3053 20819 3111 20825
rect 3988 20828 4077 20856
rect 3988 20800 4016 20828
rect 4065 20825 4077 20828
rect 4111 20825 4123 20859
rect 4065 20819 4123 20825
rect 4157 20859 4215 20865
rect 4157 20825 4169 20859
rect 4203 20856 4215 20859
rect 4246 20856 4252 20868
rect 4203 20828 4252 20856
rect 4203 20825 4215 20828
rect 4157 20819 4215 20825
rect 4246 20816 4252 20828
rect 4304 20816 4310 20868
rect 4709 20859 4767 20865
rect 4709 20825 4721 20859
rect 4755 20856 4767 20859
rect 4798 20856 4804 20868
rect 4755 20828 4804 20856
rect 4755 20825 4767 20828
rect 4709 20819 4767 20825
rect 4798 20816 4804 20828
rect 4856 20816 4862 20868
rect 5350 20856 5356 20868
rect 5311 20828 5356 20856
rect 5350 20816 5356 20828
rect 5408 20816 5414 20868
rect 7285 20859 7343 20865
rect 7285 20825 7297 20859
rect 7331 20856 7343 20859
rect 7558 20856 7564 20868
rect 7331 20828 7564 20856
rect 7331 20825 7343 20828
rect 7285 20819 7343 20825
rect 7558 20816 7564 20828
rect 7616 20816 7622 20868
rect 8481 20859 8539 20865
rect 8481 20825 8493 20859
rect 8527 20856 8539 20859
rect 8938 20856 8944 20868
rect 8527 20828 8944 20856
rect 8527 20825 8539 20828
rect 8481 20819 8539 20825
rect 8938 20816 8944 20828
rect 8996 20816 9002 20868
rect 2464 20760 2774 20788
rect 2464 20748 2470 20760
rect 3970 20748 3976 20800
rect 4028 20748 4034 20800
rect 6086 20748 6092 20800
rect 6144 20788 6150 20800
rect 6362 20788 6368 20800
rect 6144 20760 6368 20788
rect 6144 20748 6150 20760
rect 6362 20748 6368 20760
rect 6420 20748 6426 20800
rect 6549 20791 6607 20797
rect 6549 20757 6561 20791
rect 6595 20788 6607 20791
rect 9214 20788 9220 20800
rect 6595 20760 9220 20788
rect 6595 20757 6607 20760
rect 6549 20751 6607 20757
rect 9214 20748 9220 20760
rect 9272 20748 9278 20800
rect 9398 20748 9404 20800
rect 9456 20788 9462 20800
rect 9646 20788 9674 20883
rect 10134 20816 10140 20868
rect 10192 20856 10198 20868
rect 10229 20859 10287 20865
rect 10229 20856 10241 20859
rect 10192 20828 10241 20856
rect 10192 20816 10198 20828
rect 10229 20825 10241 20828
rect 10275 20825 10287 20859
rect 10229 20819 10287 20825
rect 11701 20859 11759 20865
rect 11701 20825 11713 20859
rect 11747 20825 11759 20859
rect 11701 20819 11759 20825
rect 9456 20760 9674 20788
rect 11716 20788 11744 20819
rect 11790 20816 11796 20868
rect 11848 20856 11854 20868
rect 13354 20856 13360 20868
rect 11848 20828 11893 20856
rect 12406 20828 13360 20856
rect 11848 20816 11854 20828
rect 12406 20788 12434 20828
rect 13354 20816 13360 20828
rect 13412 20816 13418 20868
rect 16408 20856 16436 20964
rect 16592 20964 18000 20992
rect 19429 20995 19487 21001
rect 16592 20936 16620 20964
rect 19429 20961 19441 20995
rect 19475 20961 19487 20995
rect 20714 20992 20720 21004
rect 20675 20964 20720 20992
rect 19429 20955 19487 20961
rect 20714 20952 20720 20964
rect 20772 20952 20778 21004
rect 38378 20992 38384 21004
rect 22664 20964 38384 20992
rect 16574 20884 16580 20936
rect 16632 20924 16638 20936
rect 16632 20896 16725 20924
rect 16632 20884 16638 20896
rect 16942 20884 16948 20936
rect 17000 20924 17006 20936
rect 17221 20927 17279 20933
rect 17221 20924 17233 20927
rect 17000 20896 17233 20924
rect 17000 20884 17006 20896
rect 17221 20893 17233 20896
rect 17267 20893 17279 20927
rect 17221 20887 17279 20893
rect 19334 20884 19340 20936
rect 19392 20924 19398 20936
rect 19613 20927 19671 20933
rect 19613 20924 19625 20927
rect 19392 20896 19625 20924
rect 19392 20884 19398 20896
rect 19613 20893 19625 20896
rect 19659 20893 19671 20927
rect 20898 20924 20904 20936
rect 20859 20896 20904 20924
rect 19613 20887 19671 20893
rect 20898 20884 20904 20896
rect 20956 20884 20962 20936
rect 22189 20927 22247 20933
rect 22189 20924 22201 20927
rect 22066 20896 22201 20924
rect 16408 20828 17908 20856
rect 13538 20788 13544 20800
rect 11716 20760 12434 20788
rect 13499 20760 13544 20788
rect 9456 20748 9462 20760
rect 13538 20748 13544 20760
rect 13596 20748 13602 20800
rect 15378 20748 15384 20800
rect 15436 20788 15442 20800
rect 15473 20791 15531 20797
rect 15473 20788 15485 20791
rect 15436 20760 15485 20788
rect 15436 20748 15442 20760
rect 15473 20757 15485 20760
rect 15519 20757 15531 20791
rect 16666 20788 16672 20800
rect 16627 20760 16672 20788
rect 15473 20751 15531 20757
rect 16666 20748 16672 20760
rect 16724 20748 16730 20800
rect 17880 20788 17908 20828
rect 17954 20816 17960 20868
rect 18012 20856 18018 20868
rect 22066 20856 22094 20896
rect 22189 20893 22201 20896
rect 22235 20893 22247 20927
rect 22370 20924 22376 20936
rect 22331 20896 22376 20924
rect 22189 20887 22247 20893
rect 22370 20884 22376 20896
rect 22428 20884 22434 20936
rect 18012 20828 22094 20856
rect 18012 20816 18018 20828
rect 20073 20791 20131 20797
rect 20073 20788 20085 20791
rect 17880 20760 20085 20788
rect 20073 20757 20085 20760
rect 20119 20788 20131 20791
rect 21361 20791 21419 20797
rect 21361 20788 21373 20791
rect 20119 20760 21373 20788
rect 20119 20757 20131 20760
rect 20073 20751 20131 20757
rect 21361 20757 21373 20760
rect 21407 20757 21419 20791
rect 21361 20751 21419 20757
rect 21450 20748 21456 20800
rect 21508 20788 21514 20800
rect 22664 20788 22692 20964
rect 38378 20952 38384 20964
rect 38436 20952 38442 21004
rect 26053 20927 26111 20933
rect 26053 20893 26065 20927
rect 26099 20893 26111 20927
rect 26053 20887 26111 20893
rect 26068 20856 26096 20887
rect 26234 20884 26240 20936
rect 26292 20924 26298 20936
rect 31297 20927 31355 20933
rect 31297 20924 31309 20927
rect 26292 20896 31309 20924
rect 26292 20884 26298 20896
rect 31297 20893 31309 20896
rect 31343 20893 31355 20927
rect 31297 20887 31355 20893
rect 37366 20884 37372 20936
rect 37424 20924 37430 20936
rect 37553 20927 37611 20933
rect 37553 20924 37565 20927
rect 37424 20896 37565 20924
rect 37424 20884 37430 20896
rect 37553 20893 37565 20896
rect 37599 20893 37611 20927
rect 38010 20924 38016 20936
rect 37971 20896 38016 20924
rect 37553 20887 37611 20893
rect 38010 20884 38016 20896
rect 38068 20884 38074 20936
rect 35342 20856 35348 20868
rect 26068 20828 35348 20856
rect 35342 20816 35348 20828
rect 35400 20816 35406 20868
rect 21508 20760 22692 20788
rect 22833 20791 22891 20797
rect 21508 20748 21514 20760
rect 22833 20757 22845 20791
rect 22879 20788 22891 20791
rect 24486 20788 24492 20800
rect 22879 20760 24492 20788
rect 22879 20757 22891 20760
rect 22833 20751 22891 20757
rect 24486 20748 24492 20760
rect 24544 20748 24550 20800
rect 24670 20748 24676 20800
rect 24728 20788 24734 20800
rect 26145 20791 26203 20797
rect 26145 20788 26157 20791
rect 24728 20760 26157 20788
rect 24728 20748 24734 20760
rect 26145 20757 26157 20760
rect 26191 20757 26203 20791
rect 38194 20788 38200 20800
rect 38155 20760 38200 20788
rect 26145 20751 26203 20757
rect 38194 20748 38200 20760
rect 38252 20748 38258 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 1578 20544 1584 20596
rect 1636 20544 1642 20596
rect 3694 20584 3700 20596
rect 1780 20556 3700 20584
rect 1596 20516 1624 20544
rect 1780 20525 1808 20556
rect 3694 20544 3700 20556
rect 3752 20544 3758 20596
rect 7098 20584 7104 20596
rect 6012 20556 7104 20584
rect 6012 20528 6040 20556
rect 7098 20544 7104 20556
rect 7156 20544 7162 20596
rect 8018 20544 8024 20596
rect 8076 20584 8082 20596
rect 13998 20584 14004 20596
rect 8076 20556 14004 20584
rect 8076 20544 8082 20556
rect 13998 20544 14004 20556
rect 14056 20544 14062 20596
rect 14093 20587 14151 20593
rect 14093 20553 14105 20587
rect 14139 20584 14151 20587
rect 14642 20584 14648 20596
rect 14139 20556 14648 20584
rect 14139 20553 14151 20556
rect 14093 20547 14151 20553
rect 14642 20544 14648 20556
rect 14700 20544 14706 20596
rect 14752 20556 15332 20584
rect 1673 20519 1731 20525
rect 1673 20516 1685 20519
rect 1596 20488 1685 20516
rect 1673 20485 1685 20488
rect 1719 20485 1731 20519
rect 1673 20479 1731 20485
rect 1765 20519 1823 20525
rect 1765 20485 1777 20519
rect 1811 20485 1823 20519
rect 3326 20516 3332 20528
rect 3287 20488 3332 20516
rect 1765 20479 1823 20485
rect 3326 20476 3332 20488
rect 3384 20476 3390 20528
rect 3881 20519 3939 20525
rect 3881 20485 3893 20519
rect 3927 20516 3939 20519
rect 4798 20516 4804 20528
rect 3927 20488 4804 20516
rect 3927 20485 3939 20488
rect 3881 20479 3939 20485
rect 4798 20476 4804 20488
rect 4856 20476 4862 20528
rect 5166 20476 5172 20528
rect 5224 20516 5230 20528
rect 5445 20519 5503 20525
rect 5445 20516 5457 20519
rect 5224 20488 5457 20516
rect 5224 20476 5230 20488
rect 5445 20485 5457 20488
rect 5491 20485 5503 20519
rect 5994 20516 6000 20528
rect 5907 20488 6000 20516
rect 5445 20479 5503 20485
rect 5994 20476 6000 20488
rect 6052 20476 6058 20528
rect 7006 20516 7012 20528
rect 6967 20488 7012 20516
rect 7006 20476 7012 20488
rect 7064 20476 7070 20528
rect 7561 20519 7619 20525
rect 7561 20485 7573 20519
rect 7607 20516 7619 20519
rect 7742 20516 7748 20528
rect 7607 20488 7748 20516
rect 7607 20485 7619 20488
rect 7561 20479 7619 20485
rect 4154 20408 4160 20460
rect 4212 20448 4218 20460
rect 4617 20451 4675 20457
rect 4617 20448 4629 20451
rect 4212 20420 4629 20448
rect 4212 20408 4218 20420
rect 4617 20417 4629 20420
rect 4663 20417 4675 20451
rect 4617 20411 4675 20417
rect 2685 20383 2743 20389
rect 2685 20349 2697 20383
rect 2731 20380 2743 20383
rect 3050 20380 3056 20392
rect 2731 20352 3056 20380
rect 2731 20349 2743 20352
rect 2685 20343 2743 20349
rect 3050 20340 3056 20352
rect 3108 20340 3114 20392
rect 3237 20383 3295 20389
rect 3237 20349 3249 20383
rect 3283 20380 3295 20383
rect 3326 20380 3332 20392
rect 3283 20352 3332 20380
rect 3283 20349 3295 20352
rect 3237 20343 3295 20349
rect 3326 20340 3332 20352
rect 3384 20340 3390 20392
rect 5353 20383 5411 20389
rect 5353 20349 5365 20383
rect 5399 20380 5411 20383
rect 6917 20383 6975 20389
rect 5399 20352 6868 20380
rect 5399 20349 5411 20352
rect 5353 20343 5411 20349
rect 6178 20312 6184 20324
rect 3988 20284 6184 20312
rect 3694 20204 3700 20256
rect 3752 20244 3758 20256
rect 3988 20244 4016 20284
rect 6178 20272 6184 20284
rect 6236 20272 6242 20324
rect 6840 20312 6868 20352
rect 6917 20349 6929 20383
rect 6963 20380 6975 20383
rect 7098 20380 7104 20392
rect 6963 20352 7104 20380
rect 6963 20349 6975 20352
rect 6917 20343 6975 20349
rect 7098 20340 7104 20352
rect 7156 20340 7162 20392
rect 7576 20312 7604 20479
rect 7742 20476 7748 20488
rect 7800 20476 7806 20528
rect 8202 20516 8208 20528
rect 8163 20488 8208 20516
rect 8202 20476 8208 20488
rect 8260 20476 8266 20528
rect 8386 20476 8392 20528
rect 8444 20516 8450 20528
rect 9401 20519 9459 20525
rect 9401 20516 9413 20519
rect 8444 20488 9413 20516
rect 8444 20476 8450 20488
rect 9401 20485 9413 20488
rect 9447 20485 9459 20519
rect 10318 20516 10324 20528
rect 10279 20488 10324 20516
rect 9401 20479 9459 20485
rect 10318 20476 10324 20488
rect 10376 20476 10382 20528
rect 11882 20516 11888 20528
rect 11843 20488 11888 20516
rect 11882 20476 11888 20488
rect 11940 20476 11946 20528
rect 11977 20519 12035 20525
rect 11977 20485 11989 20519
rect 12023 20516 12035 20519
rect 12526 20516 12532 20528
rect 12023 20488 12532 20516
rect 12023 20485 12035 20488
rect 11977 20479 12035 20485
rect 12526 20476 12532 20488
rect 12584 20476 12590 20528
rect 12986 20476 12992 20528
rect 13044 20516 13050 20528
rect 14752 20516 14780 20556
rect 15194 20516 15200 20528
rect 13044 20488 14780 20516
rect 15155 20488 15200 20516
rect 13044 20476 13050 20488
rect 15194 20476 15200 20488
rect 15252 20476 15258 20528
rect 15304 20516 15332 20556
rect 15930 20544 15936 20596
rect 15988 20584 15994 20596
rect 15988 20556 20484 20584
rect 15988 20544 15994 20556
rect 16117 20519 16175 20525
rect 15304 20488 15976 20516
rect 8754 20408 8760 20460
rect 8812 20448 8818 20460
rect 8812 20420 9168 20448
rect 8812 20408 8818 20420
rect 7926 20340 7932 20392
rect 7984 20380 7990 20392
rect 8113 20383 8171 20389
rect 8113 20380 8125 20383
rect 7984 20352 8125 20380
rect 7984 20340 7990 20352
rect 8113 20349 8125 20352
rect 8159 20349 8171 20383
rect 8846 20380 8852 20392
rect 8113 20343 8171 20349
rect 8220 20352 8852 20380
rect 6840 20284 7604 20312
rect 7742 20272 7748 20324
rect 7800 20312 7806 20324
rect 8220 20312 8248 20352
rect 8846 20340 8852 20352
rect 8904 20340 8910 20392
rect 7800 20284 8248 20312
rect 9140 20312 9168 20420
rect 10778 20408 10784 20460
rect 10836 20448 10842 20460
rect 10965 20451 11023 20457
rect 10965 20448 10977 20451
rect 10836 20420 10977 20448
rect 10836 20408 10842 20420
rect 10965 20417 10977 20420
rect 11011 20417 11023 20451
rect 10965 20411 11023 20417
rect 12802 20408 12808 20460
rect 12860 20448 12866 20460
rect 13262 20448 13268 20460
rect 12860 20420 13268 20448
rect 12860 20408 12866 20420
rect 13262 20408 13268 20420
rect 13320 20408 13326 20460
rect 13538 20408 13544 20460
rect 13596 20448 13602 20460
rect 13633 20451 13691 20457
rect 13633 20448 13645 20451
rect 13596 20420 13645 20448
rect 13596 20408 13602 20420
rect 13633 20417 13645 20420
rect 13679 20417 13691 20451
rect 15948 20448 15976 20488
rect 16117 20485 16129 20519
rect 16163 20516 16175 20519
rect 16298 20516 16304 20528
rect 16163 20488 16304 20516
rect 16163 20485 16175 20488
rect 16117 20479 16175 20485
rect 16298 20476 16304 20488
rect 16356 20476 16362 20528
rect 16390 20476 16396 20528
rect 16448 20516 16454 20528
rect 17405 20519 17463 20525
rect 17405 20516 17417 20519
rect 16448 20488 17417 20516
rect 16448 20476 16454 20488
rect 17405 20485 17417 20488
rect 17451 20485 17463 20519
rect 19518 20516 19524 20528
rect 19479 20488 19524 20516
rect 17405 20479 17463 20485
rect 19518 20476 19524 20488
rect 19576 20476 19582 20528
rect 19613 20519 19671 20525
rect 19613 20485 19625 20519
rect 19659 20516 19671 20519
rect 20456 20516 20484 20556
rect 20898 20544 20904 20596
rect 20956 20584 20962 20596
rect 21085 20587 21143 20593
rect 21085 20584 21097 20587
rect 20956 20556 21097 20584
rect 20956 20544 20962 20556
rect 21085 20553 21097 20556
rect 21131 20553 21143 20587
rect 21085 20547 21143 20553
rect 22005 20587 22063 20593
rect 22005 20553 22017 20587
rect 22051 20584 22063 20587
rect 22370 20584 22376 20596
rect 22051 20556 22376 20584
rect 22051 20553 22063 20556
rect 22005 20547 22063 20553
rect 22370 20544 22376 20556
rect 22428 20544 22434 20596
rect 37734 20584 37740 20596
rect 37695 20556 37740 20584
rect 37734 20544 37740 20556
rect 37792 20544 37798 20596
rect 38102 20516 38108 20528
rect 19659 20488 20392 20516
rect 20456 20488 21036 20516
rect 19659 20485 19671 20488
rect 19613 20479 19671 20485
rect 15948 20420 16804 20448
rect 13633 20411 13691 20417
rect 9306 20380 9312 20392
rect 9267 20352 9312 20380
rect 9306 20340 9312 20352
rect 9364 20340 9370 20392
rect 9674 20340 9680 20392
rect 9732 20380 9738 20392
rect 12161 20383 12219 20389
rect 12161 20380 12173 20383
rect 9732 20352 12173 20380
rect 9732 20340 9738 20352
rect 12161 20349 12173 20352
rect 12207 20349 12219 20383
rect 13449 20383 13507 20389
rect 13449 20380 13461 20383
rect 12161 20343 12219 20349
rect 12406 20352 13461 20380
rect 11057 20315 11115 20321
rect 9140 20284 10180 20312
rect 7800 20272 7806 20284
rect 3752 20216 4016 20244
rect 4709 20247 4767 20253
rect 3752 20204 3758 20216
rect 4709 20213 4721 20247
rect 4755 20244 4767 20247
rect 9490 20244 9496 20256
rect 4755 20216 9496 20244
rect 4755 20213 4767 20216
rect 4709 20207 4767 20213
rect 9490 20204 9496 20216
rect 9548 20204 9554 20256
rect 10152 20244 10180 20284
rect 11057 20281 11069 20315
rect 11103 20312 11115 20315
rect 12406 20312 12434 20352
rect 13449 20349 13461 20352
rect 13495 20380 13507 20383
rect 13906 20380 13912 20392
rect 13495 20352 13912 20380
rect 13495 20349 13507 20352
rect 13449 20343 13507 20349
rect 13906 20340 13912 20352
rect 13964 20340 13970 20392
rect 15105 20383 15163 20389
rect 15105 20349 15117 20383
rect 15151 20349 15163 20383
rect 15105 20343 15163 20349
rect 11103 20284 12434 20312
rect 11103 20281 11115 20284
rect 11057 20275 11115 20281
rect 12710 20272 12716 20324
rect 12768 20312 12774 20324
rect 13354 20312 13360 20324
rect 12768 20284 13360 20312
rect 12768 20272 12774 20284
rect 13354 20272 13360 20284
rect 13412 20272 13418 20324
rect 15120 20312 15148 20343
rect 16666 20312 16672 20324
rect 15120 20284 16672 20312
rect 16666 20272 16672 20284
rect 16724 20272 16730 20324
rect 16776 20312 16804 20420
rect 18690 20408 18696 20460
rect 18748 20448 18754 20460
rect 18785 20451 18843 20457
rect 18785 20448 18797 20451
rect 18748 20420 18797 20448
rect 18748 20408 18754 20420
rect 18785 20417 18797 20420
rect 18831 20417 18843 20451
rect 18785 20411 18843 20417
rect 18877 20451 18935 20457
rect 18877 20417 18889 20451
rect 18923 20448 18935 20451
rect 19334 20448 19340 20460
rect 18923 20420 19340 20448
rect 18923 20417 18935 20420
rect 18877 20411 18935 20417
rect 19334 20408 19340 20420
rect 19392 20408 19398 20460
rect 17310 20380 17316 20392
rect 17271 20352 17316 20380
rect 17310 20340 17316 20352
rect 17368 20340 17374 20392
rect 18138 20380 18144 20392
rect 18099 20352 18144 20380
rect 18138 20340 18144 20352
rect 18196 20340 18202 20392
rect 19797 20383 19855 20389
rect 19797 20380 19809 20383
rect 19306 20352 19809 20380
rect 17402 20312 17408 20324
rect 16776 20284 17408 20312
rect 17402 20272 17408 20284
rect 17460 20272 17466 20324
rect 17586 20272 17592 20324
rect 17644 20312 17650 20324
rect 19306 20312 19334 20352
rect 19797 20349 19809 20352
rect 19843 20349 19855 20383
rect 20364 20380 20392 20488
rect 21008 20457 21036 20488
rect 35866 20488 38108 20516
rect 20993 20451 21051 20457
rect 20993 20417 21005 20451
rect 21039 20417 21051 20451
rect 22186 20448 22192 20460
rect 22147 20420 22192 20448
rect 20993 20411 21051 20417
rect 22186 20408 22192 20420
rect 22244 20408 22250 20460
rect 27798 20448 27804 20460
rect 27759 20420 27804 20448
rect 27798 20408 27804 20420
rect 27856 20408 27862 20460
rect 35342 20448 35348 20460
rect 35303 20420 35348 20448
rect 35342 20408 35348 20420
rect 35400 20448 35406 20460
rect 35866 20448 35894 20488
rect 38102 20476 38108 20488
rect 38160 20476 38166 20528
rect 35400 20420 35894 20448
rect 35400 20408 35406 20420
rect 36814 20408 36820 20460
rect 36872 20448 36878 20460
rect 37921 20451 37979 20457
rect 37921 20448 37933 20451
rect 36872 20420 37933 20448
rect 36872 20408 36878 20420
rect 37921 20417 37933 20420
rect 37967 20417 37979 20451
rect 37921 20411 37979 20417
rect 22370 20380 22376 20392
rect 20364 20352 22376 20380
rect 19797 20343 19855 20349
rect 22370 20340 22376 20352
rect 22428 20340 22434 20392
rect 17644 20284 19334 20312
rect 17644 20272 17650 20284
rect 19702 20272 19708 20324
rect 19760 20312 19766 20324
rect 31110 20312 31116 20324
rect 19760 20284 31116 20312
rect 19760 20272 19766 20284
rect 31110 20272 31116 20284
rect 31168 20272 31174 20324
rect 16850 20244 16856 20256
rect 10152 20216 16856 20244
rect 16850 20204 16856 20216
rect 16908 20204 16914 20256
rect 17218 20204 17224 20256
rect 17276 20244 17282 20256
rect 22554 20244 22560 20256
rect 17276 20216 22560 20244
rect 17276 20204 17282 20216
rect 22554 20204 22560 20216
rect 22612 20204 22618 20256
rect 26786 20204 26792 20256
rect 26844 20244 26850 20256
rect 27617 20247 27675 20253
rect 27617 20244 27629 20247
rect 26844 20216 27629 20244
rect 26844 20204 26850 20216
rect 27617 20213 27629 20216
rect 27663 20213 27675 20247
rect 27617 20207 27675 20213
rect 34790 20204 34796 20256
rect 34848 20244 34854 20256
rect 35161 20247 35219 20253
rect 35161 20244 35173 20247
rect 34848 20216 35173 20244
rect 34848 20204 34854 20216
rect 35161 20213 35173 20216
rect 35207 20213 35219 20247
rect 35161 20207 35219 20213
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 2866 20000 2872 20052
rect 2924 20040 2930 20052
rect 3970 20040 3976 20052
rect 2924 20012 3976 20040
rect 2924 20000 2930 20012
rect 3970 20000 3976 20012
rect 4028 20000 4034 20052
rect 4062 20000 4068 20052
rect 4120 20040 4126 20052
rect 4522 20040 4528 20052
rect 4120 20012 4528 20040
rect 4120 20000 4126 20012
rect 4522 20000 4528 20012
rect 4580 20000 4586 20052
rect 7190 20000 7196 20052
rect 7248 20040 7254 20052
rect 7742 20040 7748 20052
rect 7248 20012 7748 20040
rect 7248 20000 7254 20012
rect 7742 20000 7748 20012
rect 7800 20000 7806 20052
rect 8202 20000 8208 20052
rect 8260 20040 8266 20052
rect 9217 20043 9275 20049
rect 9217 20040 9229 20043
rect 8260 20012 9229 20040
rect 8260 20000 8266 20012
rect 9217 20009 9229 20012
rect 9263 20009 9275 20043
rect 9217 20003 9275 20009
rect 11882 20000 11888 20052
rect 11940 20040 11946 20052
rect 17218 20040 17224 20052
rect 11940 20012 17224 20040
rect 11940 20000 11946 20012
rect 17218 20000 17224 20012
rect 17276 20000 17282 20052
rect 17402 20000 17408 20052
rect 17460 20040 17466 20052
rect 18874 20040 18880 20052
rect 17460 20012 18880 20040
rect 17460 20000 17466 20012
rect 18874 20000 18880 20012
rect 18932 20000 18938 20052
rect 37737 20043 37795 20049
rect 37737 20009 37749 20043
rect 37783 20040 37795 20043
rect 38010 20040 38016 20052
rect 37783 20012 38016 20040
rect 37783 20009 37795 20012
rect 37737 20003 37795 20009
rect 38010 20000 38016 20012
rect 38068 20000 38074 20052
rect 8754 19932 8760 19984
rect 8812 19972 8818 19984
rect 12986 19972 12992 19984
rect 8812 19944 12992 19972
rect 8812 19932 8818 19944
rect 12986 19932 12992 19944
rect 13044 19932 13050 19984
rect 20438 19972 20444 19984
rect 13096 19944 20444 19972
rect 1765 19907 1823 19913
rect 1765 19873 1777 19907
rect 1811 19904 1823 19907
rect 2130 19904 2136 19916
rect 1811 19876 2136 19904
rect 1811 19873 1823 19876
rect 1765 19867 1823 19873
rect 2130 19864 2136 19876
rect 2188 19864 2194 19916
rect 2777 19907 2835 19913
rect 2777 19873 2789 19907
rect 2823 19904 2835 19907
rect 2823 19876 3556 19904
rect 2823 19873 2835 19876
rect 2777 19867 2835 19873
rect 3237 19839 3295 19845
rect 3237 19805 3249 19839
rect 3283 19805 3295 19839
rect 3528 19836 3556 19876
rect 3602 19864 3608 19916
rect 3660 19904 3666 19916
rect 4065 19907 4123 19913
rect 4065 19904 4077 19907
rect 3660 19876 4077 19904
rect 3660 19864 3666 19876
rect 4065 19873 4077 19876
rect 4111 19873 4123 19907
rect 4065 19867 4123 19873
rect 4154 19864 4160 19916
rect 4212 19904 4218 19916
rect 4212 19876 5304 19904
rect 4212 19864 4218 19876
rect 5276 19836 5304 19876
rect 6730 19864 6736 19916
rect 6788 19904 6794 19916
rect 6788 19876 6833 19904
rect 6788 19864 6794 19876
rect 7558 19864 7564 19916
rect 7616 19904 7622 19916
rect 7929 19907 7987 19913
rect 7929 19904 7941 19907
rect 7616 19876 7941 19904
rect 7616 19864 7622 19876
rect 7929 19873 7941 19876
rect 7975 19873 7987 19907
rect 9858 19904 9864 19916
rect 9819 19876 9864 19904
rect 7929 19867 7987 19873
rect 9858 19864 9864 19876
rect 9916 19864 9922 19916
rect 10873 19907 10931 19913
rect 10873 19873 10885 19907
rect 10919 19904 10931 19907
rect 13096 19904 13124 19944
rect 20438 19932 20444 19944
rect 20496 19932 20502 19984
rect 20622 19932 20628 19984
rect 20680 19972 20686 19984
rect 20680 19944 21312 19972
rect 20680 19932 20686 19944
rect 13262 19904 13268 19916
rect 10919 19876 13124 19904
rect 13223 19876 13268 19904
rect 10919 19873 10931 19876
rect 10873 19867 10931 19873
rect 13262 19864 13268 19876
rect 13320 19864 13326 19916
rect 13998 19864 14004 19916
rect 14056 19904 14062 19916
rect 18690 19904 18696 19916
rect 14056 19876 18696 19904
rect 14056 19864 14062 19876
rect 5718 19836 5724 19848
rect 3528 19808 3924 19836
rect 5276 19808 5724 19836
rect 3237 19799 3295 19805
rect 1854 19768 1860 19780
rect 1815 19740 1860 19768
rect 1854 19728 1860 19740
rect 1912 19728 1918 19780
rect 3252 19768 3280 19799
rect 3602 19768 3608 19780
rect 3252 19740 3608 19768
rect 3602 19728 3608 19740
rect 3660 19728 3666 19780
rect 3896 19768 3924 19808
rect 5718 19796 5724 19808
rect 5776 19796 5782 19848
rect 5997 19839 6055 19845
rect 5997 19805 6009 19839
rect 6043 19836 6055 19839
rect 6178 19836 6184 19848
rect 6043 19808 6184 19836
rect 6043 19805 6055 19808
rect 5997 19799 6055 19805
rect 6178 19796 6184 19808
rect 6236 19796 6242 19848
rect 9122 19836 9128 19848
rect 9083 19808 9128 19836
rect 9122 19796 9128 19808
rect 9180 19796 9186 19848
rect 15473 19839 15531 19845
rect 15473 19805 15485 19839
rect 15519 19836 15531 19839
rect 16206 19836 16212 19848
rect 15519 19808 16212 19836
rect 15519 19805 15531 19808
rect 15473 19799 15531 19805
rect 16206 19796 16212 19808
rect 16264 19796 16270 19848
rect 18156 19845 18184 19876
rect 18690 19864 18696 19876
rect 18748 19864 18754 19916
rect 19521 19907 19579 19913
rect 19521 19873 19533 19907
rect 19567 19904 19579 19907
rect 20806 19904 20812 19916
rect 19567 19876 20812 19904
rect 19567 19873 19579 19876
rect 19521 19867 19579 19873
rect 20806 19864 20812 19876
rect 20864 19864 20870 19916
rect 21284 19913 21312 19944
rect 21269 19907 21327 19913
rect 21269 19873 21281 19907
rect 21315 19873 21327 19907
rect 22462 19904 22468 19916
rect 22423 19876 22468 19904
rect 21269 19867 21327 19873
rect 22462 19864 22468 19876
rect 22520 19864 22526 19916
rect 22646 19904 22652 19916
rect 22607 19876 22652 19904
rect 22646 19864 22652 19876
rect 22704 19864 22710 19916
rect 24946 19904 24952 19916
rect 24907 19876 24952 19904
rect 24946 19864 24952 19876
rect 25004 19864 25010 19916
rect 26786 19904 26792 19916
rect 26747 19876 26792 19904
rect 26786 19864 26792 19876
rect 26844 19864 26850 19916
rect 16301 19839 16359 19845
rect 16301 19805 16313 19839
rect 16347 19836 16359 19839
rect 16761 19839 16819 19845
rect 16761 19836 16773 19839
rect 16347 19808 16528 19836
rect 16347 19805 16359 19808
rect 16301 19799 16359 19805
rect 16500 19780 16528 19808
rect 16592 19808 16773 19836
rect 16592 19780 16620 19808
rect 16761 19805 16773 19808
rect 16807 19805 16819 19839
rect 16761 19799 16819 19805
rect 18141 19839 18199 19845
rect 18141 19805 18153 19839
rect 18187 19805 18199 19839
rect 18141 19799 18199 19805
rect 20162 19796 20168 19848
rect 20220 19836 20226 19848
rect 25961 19839 26019 19845
rect 20220 19808 20265 19836
rect 20220 19796 20226 19808
rect 25961 19805 25973 19839
rect 26007 19836 26019 19839
rect 26605 19839 26663 19845
rect 26605 19836 26617 19839
rect 26007 19808 26617 19836
rect 26007 19805 26019 19808
rect 25961 19799 26019 19805
rect 26605 19805 26617 19808
rect 26651 19805 26663 19839
rect 26605 19799 26663 19805
rect 34514 19796 34520 19848
rect 34572 19836 34578 19848
rect 36909 19839 36967 19845
rect 36909 19836 36921 19839
rect 34572 19808 36921 19836
rect 34572 19796 34578 19808
rect 36909 19805 36921 19808
rect 36955 19805 36967 19839
rect 36909 19799 36967 19805
rect 37001 19839 37059 19845
rect 37001 19805 37013 19839
rect 37047 19836 37059 19839
rect 37921 19839 37979 19845
rect 37921 19836 37933 19839
rect 37047 19808 37933 19836
rect 37047 19805 37059 19808
rect 37001 19799 37059 19805
rect 37921 19805 37933 19808
rect 37967 19805 37979 19839
rect 37921 19799 37979 19805
rect 4062 19768 4068 19780
rect 3896 19740 4068 19768
rect 4062 19728 4068 19740
rect 4120 19728 4126 19780
rect 4157 19771 4215 19777
rect 4157 19737 4169 19771
rect 4203 19768 4215 19771
rect 4890 19768 4896 19780
rect 4203 19740 4896 19768
rect 4203 19737 4215 19740
rect 4157 19731 4215 19737
rect 4890 19728 4896 19740
rect 4948 19728 4954 19780
rect 5074 19768 5080 19780
rect 5035 19740 5080 19768
rect 5074 19728 5080 19740
rect 5132 19728 5138 19780
rect 5350 19728 5356 19780
rect 5408 19768 5414 19780
rect 6454 19768 6460 19780
rect 5408 19740 6460 19768
rect 5408 19728 5414 19740
rect 6454 19728 6460 19740
rect 6512 19728 6518 19780
rect 6834 19771 6892 19777
rect 6834 19737 6846 19771
rect 6880 19768 6892 19771
rect 7377 19771 7435 19777
rect 6880 19740 6960 19768
rect 6880 19737 6892 19740
rect 6834 19731 6892 19737
rect 3329 19703 3387 19709
rect 3329 19669 3341 19703
rect 3375 19700 3387 19703
rect 5258 19700 5264 19712
rect 3375 19672 5264 19700
rect 3375 19669 3387 19672
rect 3329 19663 3387 19669
rect 5258 19660 5264 19672
rect 5316 19660 5322 19712
rect 6089 19703 6147 19709
rect 6089 19669 6101 19703
rect 6135 19700 6147 19703
rect 6932 19700 6960 19740
rect 7377 19737 7389 19771
rect 7423 19768 7435 19771
rect 7742 19768 7748 19780
rect 7423 19740 7748 19768
rect 7423 19737 7435 19740
rect 7377 19731 7435 19737
rect 7742 19728 7748 19740
rect 7800 19728 7806 19780
rect 8018 19768 8024 19780
rect 7979 19740 8024 19768
rect 8018 19728 8024 19740
rect 8076 19728 8082 19780
rect 8573 19771 8631 19777
rect 8573 19737 8585 19771
rect 8619 19768 8631 19771
rect 9674 19768 9680 19780
rect 8619 19740 9680 19768
rect 8619 19737 8631 19740
rect 8573 19731 8631 19737
rect 9674 19728 9680 19740
rect 9732 19728 9738 19780
rect 9953 19771 10011 19777
rect 9953 19768 9965 19771
rect 9784 19740 9965 19768
rect 6135 19672 6960 19700
rect 6135 19669 6147 19672
rect 6089 19663 6147 19669
rect 9214 19660 9220 19712
rect 9272 19700 9278 19712
rect 9784 19700 9812 19740
rect 9953 19737 9965 19740
rect 9999 19737 10011 19771
rect 9953 19731 10011 19737
rect 10962 19728 10968 19780
rect 11020 19768 11026 19780
rect 11793 19771 11851 19777
rect 11793 19768 11805 19771
rect 11020 19740 11805 19768
rect 11020 19728 11026 19740
rect 11793 19737 11805 19740
rect 11839 19737 11851 19771
rect 11793 19731 11851 19737
rect 11885 19771 11943 19777
rect 11885 19737 11897 19771
rect 11931 19737 11943 19771
rect 11885 19731 11943 19737
rect 9272 19672 9812 19700
rect 9272 19660 9278 19672
rect 9858 19660 9864 19712
rect 9916 19700 9922 19712
rect 10870 19700 10876 19712
rect 9916 19672 10876 19700
rect 9916 19660 9922 19672
rect 10870 19660 10876 19672
rect 10928 19660 10934 19712
rect 11900 19700 11928 19731
rect 12250 19728 12256 19780
rect 12308 19768 12314 19780
rect 12437 19771 12495 19777
rect 12437 19768 12449 19771
rect 12308 19740 12449 19768
rect 12308 19728 12314 19740
rect 12437 19737 12449 19740
rect 12483 19737 12495 19771
rect 12437 19731 12495 19737
rect 12526 19728 12532 19780
rect 12584 19768 12590 19780
rect 12989 19771 13047 19777
rect 12989 19768 13001 19771
rect 12584 19740 13001 19768
rect 12584 19728 12590 19740
rect 12989 19737 13001 19740
rect 13035 19737 13047 19771
rect 12989 19731 13047 19737
rect 13081 19771 13139 19777
rect 13081 19737 13093 19771
rect 13127 19768 13139 19771
rect 13354 19768 13360 19780
rect 13127 19740 13360 19768
rect 13127 19737 13139 19740
rect 13081 19731 13139 19737
rect 13354 19728 13360 19740
rect 13412 19728 13418 19780
rect 14366 19768 14372 19780
rect 14327 19740 14372 19768
rect 14366 19728 14372 19740
rect 14424 19728 14430 19780
rect 14461 19771 14519 19777
rect 14461 19737 14473 19771
rect 14507 19737 14519 19771
rect 15010 19768 15016 19780
rect 14971 19740 15016 19768
rect 14461 19731 14519 19737
rect 13814 19700 13820 19712
rect 11900 19672 13820 19700
rect 13814 19660 13820 19672
rect 13872 19660 13878 19712
rect 14476 19700 14504 19731
rect 15010 19728 15016 19740
rect 15068 19728 15074 19780
rect 15102 19728 15108 19780
rect 15160 19768 15166 19780
rect 15160 19740 16160 19768
rect 15160 19728 15166 19740
rect 15286 19700 15292 19712
rect 14476 19672 15292 19700
rect 15286 19660 15292 19672
rect 15344 19660 15350 19712
rect 15562 19700 15568 19712
rect 15523 19672 15568 19700
rect 15562 19660 15568 19672
rect 15620 19660 15626 19712
rect 16132 19709 16160 19740
rect 16482 19728 16488 19780
rect 16540 19728 16546 19780
rect 16574 19728 16580 19780
rect 16632 19728 16638 19780
rect 19613 19771 19671 19777
rect 19613 19737 19625 19771
rect 19659 19768 19671 19771
rect 19978 19768 19984 19780
rect 19659 19740 19984 19768
rect 19659 19737 19671 19740
rect 19613 19731 19671 19737
rect 19978 19728 19984 19740
rect 20036 19728 20042 19780
rect 20993 19771 21051 19777
rect 20993 19737 21005 19771
rect 21039 19737 21051 19771
rect 20993 19731 21051 19737
rect 16117 19703 16175 19709
rect 16117 19669 16129 19703
rect 16163 19669 16175 19703
rect 16117 19663 16175 19669
rect 16758 19660 16764 19712
rect 16816 19700 16822 19712
rect 16853 19703 16911 19709
rect 16853 19700 16865 19703
rect 16816 19672 16865 19700
rect 16816 19660 16822 19672
rect 16853 19669 16865 19672
rect 16899 19669 16911 19703
rect 16853 19663 16911 19669
rect 17034 19660 17040 19712
rect 17092 19700 17098 19712
rect 18233 19703 18291 19709
rect 18233 19700 18245 19703
rect 17092 19672 18245 19700
rect 17092 19660 17098 19672
rect 18233 19669 18245 19672
rect 18279 19669 18291 19703
rect 21008 19700 21036 19731
rect 21082 19728 21088 19780
rect 21140 19768 21146 19780
rect 21140 19740 21185 19768
rect 21140 19728 21146 19740
rect 24394 19728 24400 19780
rect 24452 19768 24458 19780
rect 24670 19768 24676 19780
rect 24452 19740 24676 19768
rect 24452 19728 24458 19740
rect 24670 19728 24676 19740
rect 24728 19728 24734 19780
rect 24762 19728 24768 19780
rect 24820 19768 24826 19780
rect 24820 19740 24865 19768
rect 24820 19728 24826 19740
rect 22554 19700 22560 19712
rect 21008 19672 22560 19700
rect 18233 19663 18291 19669
rect 22554 19660 22560 19672
rect 22612 19660 22618 19712
rect 23109 19703 23167 19709
rect 23109 19669 23121 19703
rect 23155 19700 23167 19703
rect 23934 19700 23940 19712
rect 23155 19672 23940 19700
rect 23155 19669 23167 19672
rect 23109 19663 23167 19669
rect 23934 19660 23940 19672
rect 23992 19700 23998 19712
rect 24578 19700 24584 19712
rect 23992 19672 24584 19700
rect 23992 19660 23998 19672
rect 24578 19660 24584 19672
rect 24636 19660 24642 19712
rect 27246 19700 27252 19712
rect 27207 19672 27252 19700
rect 27246 19660 27252 19672
rect 27304 19660 27310 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 3050 19456 3056 19508
rect 3108 19496 3114 19508
rect 4709 19499 4767 19505
rect 3108 19468 3832 19496
rect 3108 19456 3114 19468
rect 1673 19431 1731 19437
rect 1673 19397 1685 19431
rect 1719 19428 1731 19431
rect 2774 19428 2780 19440
rect 1719 19400 2780 19428
rect 1719 19397 1731 19400
rect 1673 19391 1731 19397
rect 2774 19388 2780 19400
rect 2832 19388 2838 19440
rect 2869 19431 2927 19437
rect 2869 19397 2881 19431
rect 2915 19428 2927 19431
rect 3142 19428 3148 19440
rect 2915 19400 3148 19428
rect 2915 19397 2927 19400
rect 2869 19391 2927 19397
rect 3142 19388 3148 19400
rect 3200 19388 3206 19440
rect 3804 19437 3832 19468
rect 4709 19465 4721 19499
rect 4755 19496 4767 19499
rect 7006 19496 7012 19508
rect 4755 19468 7012 19496
rect 4755 19465 4767 19468
rect 4709 19459 4767 19465
rect 7006 19456 7012 19468
rect 7064 19456 7070 19508
rect 10410 19496 10416 19508
rect 7116 19468 10416 19496
rect 3789 19431 3847 19437
rect 3789 19397 3801 19431
rect 3835 19428 3847 19431
rect 5166 19428 5172 19440
rect 3835 19400 5172 19428
rect 3835 19397 3847 19400
rect 3789 19391 3847 19397
rect 5166 19388 5172 19400
rect 5224 19388 5230 19440
rect 5442 19428 5448 19440
rect 5403 19400 5448 19428
rect 5442 19388 5448 19400
rect 5500 19388 5506 19440
rect 5994 19428 6000 19440
rect 5955 19400 6000 19428
rect 5994 19388 6000 19400
rect 6052 19388 6058 19440
rect 6454 19388 6460 19440
rect 6512 19428 6518 19440
rect 6641 19431 6699 19437
rect 6641 19428 6653 19431
rect 6512 19400 6653 19428
rect 6512 19388 6518 19400
rect 6641 19397 6653 19400
rect 6687 19397 6699 19431
rect 6641 19391 6699 19397
rect 4617 19363 4675 19369
rect 4617 19329 4629 19363
rect 4663 19360 4675 19363
rect 4890 19360 4896 19372
rect 4663 19332 4896 19360
rect 4663 19329 4675 19332
rect 4617 19323 4675 19329
rect 4890 19320 4896 19332
rect 4948 19320 4954 19372
rect 6549 19363 6607 19369
rect 6549 19329 6561 19363
rect 6595 19360 6607 19363
rect 7116 19360 7144 19468
rect 10410 19456 10416 19468
rect 10468 19496 10474 19508
rect 13354 19496 13360 19508
rect 10468 19468 11008 19496
rect 10468 19456 10474 19468
rect 7374 19428 7380 19440
rect 7335 19400 7380 19428
rect 7374 19388 7380 19400
rect 7432 19388 7438 19440
rect 9030 19428 9036 19440
rect 8991 19400 9036 19428
rect 9030 19388 9036 19400
rect 9088 19388 9094 19440
rect 9490 19388 9496 19440
rect 9548 19388 9554 19440
rect 10980 19428 11008 19468
rect 11808 19468 13360 19496
rect 11808 19437 11836 19468
rect 13354 19456 13360 19468
rect 13412 19456 13418 19508
rect 14274 19496 14280 19508
rect 13464 19468 14280 19496
rect 11793 19431 11851 19437
rect 10980 19400 11652 19428
rect 10980 19369 11008 19400
rect 6595 19332 7144 19360
rect 10965 19363 11023 19369
rect 6595 19329 6607 19332
rect 6549 19323 6607 19329
rect 10965 19329 10977 19363
rect 11011 19329 11023 19363
rect 10965 19323 11023 19329
rect 11054 19320 11060 19372
rect 11112 19360 11118 19372
rect 11112 19332 11157 19360
rect 11112 19320 11118 19332
rect 2777 19295 2835 19301
rect 2777 19261 2789 19295
rect 2823 19292 2835 19295
rect 2958 19292 2964 19304
rect 2823 19264 2964 19292
rect 2823 19261 2835 19264
rect 2777 19255 2835 19261
rect 2958 19252 2964 19264
rect 3016 19252 3022 19304
rect 3878 19252 3884 19304
rect 3936 19292 3942 19304
rect 5074 19292 5080 19304
rect 3936 19264 5080 19292
rect 3936 19252 3942 19264
rect 5074 19252 5080 19264
rect 5132 19252 5138 19304
rect 5350 19292 5356 19304
rect 5311 19264 5356 19292
rect 5350 19252 5356 19264
rect 5408 19252 5414 19304
rect 5718 19252 5724 19304
rect 5776 19292 5782 19304
rect 6822 19292 6828 19304
rect 5776 19264 6828 19292
rect 5776 19252 5782 19264
rect 6822 19252 6828 19264
rect 6880 19292 6886 19304
rect 7285 19295 7343 19301
rect 7285 19292 7297 19295
rect 6880 19264 7297 19292
rect 6880 19252 6886 19264
rect 7285 19261 7297 19264
rect 7331 19261 7343 19295
rect 7285 19255 7343 19261
rect 7466 19252 7472 19304
rect 7524 19292 7530 19304
rect 7561 19295 7619 19301
rect 7561 19292 7573 19295
rect 7524 19264 7573 19292
rect 7524 19252 7530 19264
rect 7561 19261 7573 19264
rect 7607 19261 7619 19295
rect 8754 19292 8760 19304
rect 8715 19264 8760 19292
rect 7561 19255 7619 19261
rect 8754 19252 8760 19264
rect 8812 19252 8818 19304
rect 8864 19264 10088 19292
rect 1857 19227 1915 19233
rect 1857 19193 1869 19227
rect 1903 19224 1915 19227
rect 2222 19224 2228 19236
rect 1903 19196 2228 19224
rect 1903 19193 1915 19196
rect 1857 19187 1915 19193
rect 2222 19184 2228 19196
rect 2280 19184 2286 19236
rect 3970 19184 3976 19236
rect 4028 19224 4034 19236
rect 8864 19224 8892 19264
rect 4028 19196 8892 19224
rect 10060 19224 10088 19264
rect 10318 19252 10324 19304
rect 10376 19292 10382 19304
rect 10686 19292 10692 19304
rect 10376 19264 10692 19292
rect 10376 19252 10382 19264
rect 10686 19252 10692 19264
rect 10744 19252 10750 19304
rect 11624 19292 11652 19400
rect 11793 19397 11805 19431
rect 11839 19397 11851 19431
rect 11793 19391 11851 19397
rect 11885 19431 11943 19437
rect 11885 19397 11897 19431
rect 11931 19428 11943 19431
rect 11974 19428 11980 19440
rect 11931 19400 11980 19428
rect 11931 19397 11943 19400
rect 11885 19391 11943 19397
rect 11974 19388 11980 19400
rect 12032 19388 12038 19440
rect 12066 19388 12072 19440
rect 12124 19428 12130 19440
rect 13464 19428 13492 19468
rect 14274 19456 14280 19468
rect 14332 19456 14338 19508
rect 17402 19496 17408 19508
rect 15396 19468 17408 19496
rect 14001 19431 14059 19437
rect 14001 19428 14013 19431
rect 12124 19400 13492 19428
rect 13556 19400 14013 19428
rect 12124 19388 12130 19400
rect 13078 19320 13084 19372
rect 13136 19360 13142 19372
rect 13173 19363 13231 19369
rect 13173 19360 13185 19363
rect 13136 19332 13185 19360
rect 13136 19320 13142 19332
rect 13173 19329 13185 19332
rect 13219 19360 13231 19363
rect 13446 19360 13452 19372
rect 13219 19332 13452 19360
rect 13219 19329 13231 19332
rect 13173 19323 13231 19329
rect 13446 19320 13452 19332
rect 13504 19320 13510 19372
rect 12066 19292 12072 19304
rect 11624 19264 12072 19292
rect 12066 19252 12072 19264
rect 12124 19252 12130 19304
rect 12161 19295 12219 19301
rect 12161 19261 12173 19295
rect 12207 19292 12219 19295
rect 12802 19292 12808 19304
rect 12207 19264 12808 19292
rect 12207 19261 12219 19264
rect 12161 19255 12219 19261
rect 12176 19224 12204 19255
rect 12802 19252 12808 19264
rect 12860 19252 12866 19304
rect 13265 19295 13323 19301
rect 13265 19261 13277 19295
rect 13311 19292 13323 19295
rect 13556 19292 13584 19400
rect 14001 19397 14013 19400
rect 14047 19397 14059 19431
rect 15396 19428 15424 19468
rect 17402 19456 17408 19468
rect 17460 19456 17466 19508
rect 20346 19496 20352 19508
rect 18340 19468 20352 19496
rect 15562 19428 15568 19440
rect 14001 19391 14059 19397
rect 15304 19400 15424 19428
rect 15523 19400 15568 19428
rect 13906 19292 13912 19304
rect 13311 19264 13584 19292
rect 13867 19264 13912 19292
rect 13311 19261 13323 19264
rect 13265 19255 13323 19261
rect 13906 19252 13912 19264
rect 13964 19252 13970 19304
rect 14366 19292 14372 19304
rect 14327 19264 14372 19292
rect 14366 19252 14372 19264
rect 14424 19252 14430 19304
rect 15194 19292 15200 19304
rect 14752 19264 15200 19292
rect 10060 19196 12204 19224
rect 4028 19184 4034 19196
rect 12342 19184 12348 19236
rect 12400 19224 12406 19236
rect 14752 19224 14780 19264
rect 15194 19252 15200 19264
rect 15252 19252 15258 19304
rect 15304 19292 15332 19400
rect 15562 19388 15568 19400
rect 15620 19388 15626 19440
rect 17034 19428 17040 19440
rect 16995 19400 17040 19428
rect 17034 19388 17040 19400
rect 17092 19388 17098 19440
rect 18340 19437 18368 19468
rect 20346 19456 20352 19468
rect 20404 19456 20410 19508
rect 20438 19456 20444 19508
rect 20496 19496 20502 19508
rect 23106 19496 23112 19508
rect 20496 19468 23112 19496
rect 20496 19456 20502 19468
rect 23106 19456 23112 19468
rect 23164 19456 23170 19508
rect 26053 19499 26111 19505
rect 26053 19465 26065 19499
rect 26099 19465 26111 19499
rect 36814 19496 36820 19508
rect 36775 19468 36820 19496
rect 26053 19459 26111 19465
rect 18325 19431 18383 19437
rect 18325 19397 18337 19431
rect 18371 19397 18383 19431
rect 18325 19391 18383 19397
rect 18417 19431 18475 19437
rect 18417 19397 18429 19431
rect 18463 19428 18475 19431
rect 19889 19431 19947 19437
rect 19889 19428 19901 19431
rect 18463 19400 19901 19428
rect 18463 19397 18475 19400
rect 18417 19391 18475 19397
rect 19889 19397 19901 19400
rect 19935 19397 19947 19431
rect 19889 19391 19947 19397
rect 16666 19320 16672 19372
rect 16724 19360 16730 19372
rect 19797 19363 19855 19369
rect 16724 19332 16804 19360
rect 16724 19320 16730 19332
rect 15473 19295 15531 19301
rect 15473 19292 15485 19295
rect 15304 19264 15485 19292
rect 15473 19261 15485 19264
rect 15519 19261 15531 19295
rect 15473 19255 15531 19261
rect 15749 19295 15807 19301
rect 15749 19261 15761 19295
rect 15795 19261 15807 19295
rect 16776 19292 16804 19332
rect 19797 19329 19809 19363
rect 19843 19360 19855 19363
rect 20438 19360 20444 19372
rect 19843 19332 20444 19360
rect 19843 19329 19855 19332
rect 19797 19323 19855 19329
rect 20438 19320 20444 19332
rect 20496 19320 20502 19372
rect 24118 19360 24124 19372
rect 24079 19332 24124 19360
rect 24118 19320 24124 19332
rect 24176 19360 24182 19372
rect 25593 19363 25651 19369
rect 24176 19332 25544 19360
rect 24176 19320 24182 19332
rect 16945 19295 17003 19301
rect 16945 19292 16957 19295
rect 16776 19264 16957 19292
rect 15749 19255 15807 19261
rect 16945 19261 16957 19264
rect 16991 19261 17003 19295
rect 17310 19292 17316 19304
rect 17271 19264 17316 19292
rect 16945 19255 17003 19261
rect 12400 19196 14780 19224
rect 12400 19184 12406 19196
rect 14826 19184 14832 19236
rect 14884 19224 14890 19236
rect 15764 19224 15792 19255
rect 17310 19252 17316 19264
rect 17368 19252 17374 19304
rect 19245 19295 19303 19301
rect 19245 19261 19257 19295
rect 19291 19292 19303 19295
rect 20346 19292 20352 19304
rect 19291 19264 20352 19292
rect 19291 19261 19303 19264
rect 19245 19255 19303 19261
rect 20346 19252 20352 19264
rect 20404 19292 20410 19304
rect 20622 19292 20628 19304
rect 20404 19264 20628 19292
rect 20404 19252 20410 19264
rect 20622 19252 20628 19264
rect 20680 19252 20686 19304
rect 24670 19252 24676 19304
rect 24728 19292 24734 19304
rect 24765 19295 24823 19301
rect 24765 19292 24777 19295
rect 24728 19264 24777 19292
rect 24728 19252 24734 19264
rect 24765 19261 24777 19264
rect 24811 19261 24823 19295
rect 25516 19292 25544 19332
rect 25593 19329 25605 19363
rect 25639 19360 25651 19363
rect 26068 19360 26096 19459
rect 36814 19456 36820 19468
rect 36872 19456 36878 19508
rect 37826 19496 37832 19508
rect 37787 19468 37832 19496
rect 37826 19456 37832 19468
rect 37884 19456 37890 19508
rect 26237 19363 26295 19369
rect 26237 19360 26249 19363
rect 25639 19332 26096 19360
rect 26160 19332 26249 19360
rect 25639 19329 25651 19332
rect 25593 19323 25651 19329
rect 26160 19292 26188 19332
rect 26237 19329 26249 19332
rect 26283 19329 26295 19363
rect 26237 19323 26295 19329
rect 27706 19320 27712 19372
rect 27764 19360 27770 19372
rect 36725 19363 36783 19369
rect 36725 19360 36737 19363
rect 27764 19332 36737 19360
rect 27764 19320 27770 19332
rect 36725 19329 36737 19332
rect 36771 19329 36783 19363
rect 38010 19360 38016 19372
rect 37971 19332 38016 19360
rect 36725 19323 36783 19329
rect 38010 19320 38016 19332
rect 38068 19320 38074 19372
rect 25516 19264 26188 19292
rect 24765 19255 24823 19261
rect 14884 19196 15792 19224
rect 14884 19184 14890 19196
rect 16850 19184 16856 19236
rect 16908 19224 16914 19236
rect 17328 19224 17356 19252
rect 16908 19196 17356 19224
rect 16908 19184 16914 19196
rect 23198 19184 23204 19236
rect 23256 19224 23262 19236
rect 26234 19224 26240 19236
rect 23256 19196 26240 19224
rect 23256 19184 23262 19196
rect 26234 19184 26240 19196
rect 26292 19184 26298 19236
rect 4062 19116 4068 19168
rect 4120 19156 4126 19168
rect 6546 19156 6552 19168
rect 4120 19128 6552 19156
rect 4120 19116 4126 19128
rect 6546 19116 6552 19128
rect 6604 19116 6610 19168
rect 6638 19116 6644 19168
rect 6696 19156 6702 19168
rect 10226 19156 10232 19168
rect 6696 19128 10232 19156
rect 6696 19116 6702 19128
rect 10226 19116 10232 19128
rect 10284 19116 10290 19168
rect 10502 19156 10508 19168
rect 10463 19128 10508 19156
rect 10502 19116 10508 19128
rect 10560 19116 10566 19168
rect 10962 19116 10968 19168
rect 11020 19156 11026 19168
rect 17218 19156 17224 19168
rect 11020 19128 17224 19156
rect 11020 19116 11026 19128
rect 17218 19116 17224 19128
rect 17276 19116 17282 19168
rect 17954 19116 17960 19168
rect 18012 19156 18018 19168
rect 18414 19156 18420 19168
rect 18012 19128 18420 19156
rect 18012 19116 18018 19128
rect 18414 19116 18420 19128
rect 18472 19156 18478 19168
rect 19242 19156 19248 19168
rect 18472 19128 19248 19156
rect 18472 19116 18478 19128
rect 19242 19116 19248 19128
rect 19300 19116 19306 19168
rect 23474 19116 23480 19168
rect 23532 19156 23538 19168
rect 24213 19159 24271 19165
rect 24213 19156 24225 19159
rect 23532 19128 24225 19156
rect 23532 19116 23538 19128
rect 24213 19125 24225 19128
rect 24259 19125 24271 19159
rect 24213 19119 24271 19125
rect 24854 19116 24860 19168
rect 24912 19156 24918 19168
rect 25409 19159 25467 19165
rect 25409 19156 25421 19159
rect 24912 19128 25421 19156
rect 24912 19116 24918 19128
rect 25409 19125 25421 19128
rect 25455 19125 25467 19159
rect 25409 19119 25467 19125
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 4341 18955 4399 18961
rect 4341 18921 4353 18955
rect 4387 18952 4399 18955
rect 5350 18952 5356 18964
rect 4387 18924 5356 18952
rect 4387 18921 4399 18924
rect 4341 18915 4399 18921
rect 5350 18912 5356 18924
rect 5408 18912 5414 18964
rect 5442 18912 5448 18964
rect 5500 18952 5506 18964
rect 7282 18952 7288 18964
rect 5500 18924 7288 18952
rect 5500 18912 5506 18924
rect 7282 18912 7288 18924
rect 7340 18952 7346 18964
rect 7742 18952 7748 18964
rect 7340 18924 7748 18952
rect 7340 18912 7346 18924
rect 7742 18912 7748 18924
rect 7800 18912 7806 18964
rect 10042 18952 10048 18964
rect 9232 18924 10048 18952
rect 2958 18844 2964 18896
rect 3016 18884 3022 18896
rect 3016 18856 6132 18884
rect 3016 18844 3022 18856
rect 2225 18819 2283 18825
rect 2225 18785 2237 18819
rect 2271 18816 2283 18819
rect 3234 18816 3240 18828
rect 2271 18788 3240 18816
rect 2271 18785 2283 18788
rect 2225 18779 2283 18785
rect 3234 18776 3240 18788
rect 3292 18776 3298 18828
rect 4985 18819 5043 18825
rect 4985 18785 4997 18819
rect 5031 18816 5043 18819
rect 5166 18816 5172 18828
rect 5031 18788 5172 18816
rect 5031 18785 5043 18788
rect 4985 18779 5043 18785
rect 5166 18776 5172 18788
rect 5224 18776 5230 18828
rect 5629 18819 5687 18825
rect 5629 18785 5641 18819
rect 5675 18816 5687 18819
rect 5994 18816 6000 18828
rect 5675 18788 6000 18816
rect 5675 18785 5687 18788
rect 5629 18779 5687 18785
rect 5994 18776 6000 18788
rect 6052 18776 6058 18828
rect 6104 18816 6132 18856
rect 6546 18844 6552 18896
rect 6604 18884 6610 18896
rect 7190 18884 7196 18896
rect 6604 18856 7196 18884
rect 6604 18844 6610 18856
rect 7190 18844 7196 18856
rect 7248 18844 7254 18896
rect 7466 18844 7472 18896
rect 7524 18884 7530 18896
rect 9232 18884 9260 18924
rect 10042 18912 10048 18924
rect 10100 18912 10106 18964
rect 10134 18912 10140 18964
rect 10192 18952 10198 18964
rect 10873 18955 10931 18961
rect 10873 18952 10885 18955
rect 10192 18924 10885 18952
rect 10192 18912 10198 18924
rect 10873 18921 10885 18924
rect 10919 18952 10931 18955
rect 11422 18952 11428 18964
rect 10919 18924 11428 18952
rect 10919 18921 10931 18924
rect 10873 18915 10931 18921
rect 11422 18912 11428 18924
rect 11480 18912 11486 18964
rect 11882 18912 11888 18964
rect 11940 18952 11946 18964
rect 12250 18952 12256 18964
rect 11940 18924 12256 18952
rect 11940 18912 11946 18924
rect 12250 18912 12256 18924
rect 12308 18952 12314 18964
rect 17678 18952 17684 18964
rect 12308 18924 17684 18952
rect 12308 18912 12314 18924
rect 17678 18912 17684 18924
rect 17736 18912 17742 18964
rect 21542 18952 21548 18964
rect 21503 18924 21548 18952
rect 21542 18912 21548 18924
rect 21600 18912 21606 18964
rect 26234 18952 26240 18964
rect 22940 18924 26240 18952
rect 13170 18884 13176 18896
rect 7524 18856 9260 18884
rect 10428 18856 13176 18884
rect 7524 18844 7530 18856
rect 6104 18788 6592 18816
rect 4246 18748 4252 18760
rect 4159 18720 4252 18748
rect 4246 18708 4252 18720
rect 4304 18708 4310 18760
rect 6089 18751 6147 18757
rect 6089 18717 6101 18751
rect 6135 18748 6147 18751
rect 6362 18748 6368 18760
rect 6135 18720 6368 18748
rect 6135 18717 6147 18720
rect 6089 18711 6147 18717
rect 6362 18708 6368 18720
rect 6420 18708 6426 18760
rect 2314 18640 2320 18692
rect 2372 18680 2378 18692
rect 2869 18683 2927 18689
rect 2372 18652 2417 18680
rect 2372 18640 2378 18652
rect 2869 18649 2881 18683
rect 2915 18680 2927 18683
rect 4154 18680 4160 18692
rect 2915 18652 4160 18680
rect 2915 18649 2927 18652
rect 2869 18643 2927 18649
rect 4154 18640 4160 18652
rect 4212 18640 4218 18692
rect 1486 18572 1492 18624
rect 1544 18612 1550 18624
rect 4264 18612 4292 18708
rect 5074 18640 5080 18692
rect 5132 18680 5138 18692
rect 6564 18680 6592 18788
rect 8570 18776 8576 18828
rect 8628 18816 8634 18828
rect 9401 18819 9459 18825
rect 9401 18816 9413 18819
rect 8628 18788 9413 18816
rect 8628 18776 8634 18788
rect 9401 18785 9413 18788
rect 9447 18816 9459 18819
rect 10428 18816 10456 18856
rect 13170 18844 13176 18856
rect 13228 18844 13234 18896
rect 14734 18844 14740 18896
rect 14792 18884 14798 18896
rect 22940 18884 22968 18924
rect 26234 18912 26240 18924
rect 26292 18912 26298 18964
rect 37461 18955 37519 18961
rect 28966 18924 35894 18952
rect 14792 18856 22968 18884
rect 14792 18844 14798 18856
rect 23934 18844 23940 18896
rect 23992 18884 23998 18896
rect 28966 18884 28994 18924
rect 23992 18856 28994 18884
rect 35866 18884 35894 18924
rect 37461 18921 37473 18955
rect 37507 18952 37519 18955
rect 38562 18952 38568 18964
rect 37507 18924 38568 18952
rect 37507 18921 37519 18924
rect 37461 18915 37519 18921
rect 38562 18912 38568 18924
rect 38620 18912 38626 18964
rect 38194 18884 38200 18896
rect 35866 18856 38200 18884
rect 23992 18844 23998 18856
rect 38194 18844 38200 18856
rect 38252 18844 38258 18896
rect 11514 18816 11520 18828
rect 9447 18788 10456 18816
rect 11475 18788 11520 18816
rect 9447 18785 9459 18788
rect 9401 18779 9459 18785
rect 11514 18776 11520 18788
rect 11572 18776 11578 18828
rect 12250 18776 12256 18828
rect 12308 18816 12314 18828
rect 12526 18816 12532 18828
rect 12308 18788 12532 18816
rect 12308 18776 12314 18788
rect 12526 18776 12532 18788
rect 12584 18776 12590 18828
rect 12713 18819 12771 18825
rect 12713 18785 12725 18819
rect 12759 18816 12771 18819
rect 12986 18816 12992 18828
rect 12759 18788 12992 18816
rect 12759 18785 12771 18788
rect 12713 18779 12771 18785
rect 12986 18776 12992 18788
rect 13044 18776 13050 18828
rect 13078 18776 13084 18828
rect 13136 18816 13142 18828
rect 13538 18816 13544 18828
rect 13136 18788 13544 18816
rect 13136 18776 13142 18788
rect 13538 18776 13544 18788
rect 13596 18776 13602 18828
rect 15838 18776 15844 18828
rect 15896 18816 15902 18828
rect 21542 18816 21548 18828
rect 15896 18788 21548 18816
rect 15896 18776 15902 18788
rect 21542 18776 21548 18788
rect 21600 18776 21606 18828
rect 24670 18816 24676 18828
rect 24631 18788 24676 18816
rect 24670 18776 24676 18788
rect 24728 18776 24734 18828
rect 8389 18751 8447 18757
rect 8389 18717 8401 18751
rect 8435 18717 8447 18751
rect 8389 18711 8447 18717
rect 6825 18683 6883 18689
rect 6825 18680 6837 18683
rect 5132 18652 5177 18680
rect 6564 18652 6837 18680
rect 5132 18640 5138 18652
rect 6825 18649 6837 18652
rect 6871 18649 6883 18683
rect 6825 18643 6883 18649
rect 6917 18683 6975 18689
rect 6917 18649 6929 18683
rect 6963 18680 6975 18683
rect 7006 18680 7012 18692
rect 6963 18652 7012 18680
rect 6963 18649 6975 18652
rect 6917 18643 6975 18649
rect 7006 18640 7012 18652
rect 7064 18640 7070 18692
rect 7282 18640 7288 18692
rect 7340 18680 7346 18692
rect 7466 18680 7472 18692
rect 7340 18652 7472 18680
rect 7340 18640 7346 18652
rect 7466 18640 7472 18652
rect 7524 18640 7530 18692
rect 7837 18683 7895 18689
rect 7837 18649 7849 18683
rect 7883 18680 7895 18683
rect 8018 18680 8024 18692
rect 7883 18652 8024 18680
rect 7883 18649 7895 18652
rect 7837 18643 7895 18649
rect 8018 18640 8024 18652
rect 8076 18640 8082 18692
rect 8404 18680 8432 18711
rect 8846 18708 8852 18760
rect 8904 18748 8910 18760
rect 9125 18751 9183 18757
rect 9125 18748 9137 18751
rect 8904 18720 9137 18748
rect 8904 18708 8910 18720
rect 9125 18717 9137 18720
rect 9171 18717 9183 18751
rect 9125 18711 9183 18717
rect 12161 18751 12219 18757
rect 12161 18717 12173 18751
rect 12207 18748 12219 18751
rect 12342 18748 12348 18760
rect 12207 18720 12348 18748
rect 12207 18717 12219 18720
rect 12161 18711 12219 18717
rect 12342 18708 12348 18720
rect 12400 18708 12406 18760
rect 13906 18708 13912 18760
rect 13964 18748 13970 18760
rect 14369 18751 14427 18757
rect 14369 18748 14381 18751
rect 13964 18720 14381 18748
rect 13964 18708 13970 18720
rect 14369 18717 14381 18720
rect 14415 18717 14427 18751
rect 14369 18711 14427 18717
rect 16025 18751 16083 18757
rect 16025 18717 16037 18751
rect 16071 18748 16083 18751
rect 16206 18748 16212 18760
rect 16071 18720 16212 18748
rect 16071 18717 16083 18720
rect 16025 18711 16083 18717
rect 16206 18708 16212 18720
rect 16264 18708 16270 18760
rect 16666 18708 16672 18760
rect 16724 18748 16730 18760
rect 16942 18748 16948 18760
rect 16724 18720 16948 18748
rect 16724 18708 16730 18720
rect 16942 18708 16948 18720
rect 17000 18708 17006 18760
rect 17954 18748 17960 18760
rect 17052 18720 17960 18748
rect 9398 18680 9404 18692
rect 8404 18652 9404 18680
rect 9398 18640 9404 18652
rect 9456 18640 9462 18692
rect 9858 18640 9864 18692
rect 9916 18640 9922 18692
rect 11609 18683 11667 18689
rect 11609 18680 11621 18683
rect 11440 18652 11621 18680
rect 11440 18624 11468 18652
rect 11609 18649 11621 18652
rect 11655 18649 11667 18683
rect 12802 18680 12808 18692
rect 12763 18652 12808 18680
rect 11609 18643 11667 18649
rect 12802 18640 12808 18652
rect 12860 18640 12866 18692
rect 13630 18640 13636 18692
rect 13688 18680 13694 18692
rect 15378 18680 15384 18692
rect 13688 18652 14596 18680
rect 15339 18652 15384 18680
rect 13688 18640 13694 18652
rect 1544 18584 4292 18612
rect 6181 18615 6239 18621
rect 1544 18572 1550 18584
rect 6181 18581 6193 18615
rect 6227 18612 6239 18615
rect 8294 18612 8300 18624
rect 6227 18584 8300 18612
rect 6227 18581 6239 18584
rect 6181 18575 6239 18581
rect 8294 18572 8300 18584
rect 8352 18572 8358 18624
rect 8481 18615 8539 18621
rect 8481 18581 8493 18615
rect 8527 18612 8539 18615
rect 10042 18612 10048 18624
rect 8527 18584 10048 18612
rect 8527 18581 8539 18584
rect 8481 18575 8539 18581
rect 10042 18572 10048 18584
rect 10100 18572 10106 18624
rect 10318 18572 10324 18624
rect 10376 18612 10382 18624
rect 10870 18612 10876 18624
rect 10376 18584 10876 18612
rect 10376 18572 10382 18584
rect 10870 18572 10876 18584
rect 10928 18572 10934 18624
rect 11422 18572 11428 18624
rect 11480 18572 11486 18624
rect 11514 18572 11520 18624
rect 11572 18612 11578 18624
rect 12250 18612 12256 18624
rect 11572 18584 12256 18612
rect 11572 18572 11578 18584
rect 12250 18572 12256 18584
rect 12308 18572 12314 18624
rect 14458 18612 14464 18624
rect 14419 18584 14464 18612
rect 14458 18572 14464 18584
rect 14516 18572 14522 18624
rect 14568 18612 14596 18652
rect 15378 18640 15384 18652
rect 15436 18640 15442 18692
rect 15470 18640 15476 18692
rect 15528 18680 15534 18692
rect 17052 18680 17080 18720
rect 17954 18708 17960 18720
rect 18012 18708 18018 18760
rect 18138 18708 18144 18760
rect 18196 18748 18202 18760
rect 18233 18751 18291 18757
rect 18233 18748 18245 18751
rect 18196 18720 18245 18748
rect 18196 18708 18202 18720
rect 18233 18717 18245 18720
rect 18279 18748 18291 18751
rect 18414 18748 18420 18760
rect 18279 18720 18420 18748
rect 18279 18717 18291 18720
rect 18233 18711 18291 18717
rect 18414 18708 18420 18720
rect 18472 18708 18478 18760
rect 20254 18708 20260 18760
rect 20312 18748 20318 18760
rect 21453 18751 21511 18757
rect 21453 18748 21465 18751
rect 20312 18720 21465 18748
rect 20312 18708 20318 18720
rect 21453 18717 21465 18720
rect 21499 18717 21511 18751
rect 21453 18711 21511 18717
rect 26234 18708 26240 18760
rect 26292 18748 26298 18760
rect 26789 18751 26847 18757
rect 26789 18748 26801 18751
rect 26292 18720 26801 18748
rect 26292 18708 26298 18720
rect 26789 18717 26801 18720
rect 26835 18748 26847 18751
rect 27982 18748 27988 18760
rect 26835 18720 27988 18748
rect 26835 18717 26847 18720
rect 26789 18711 26847 18717
rect 27982 18708 27988 18720
rect 28040 18708 28046 18760
rect 37458 18708 37464 18760
rect 37516 18748 37522 18760
rect 37645 18751 37703 18757
rect 37645 18748 37657 18751
rect 37516 18720 37657 18748
rect 37516 18708 37522 18720
rect 37645 18717 37657 18720
rect 37691 18717 37703 18751
rect 38286 18748 38292 18760
rect 38247 18720 38292 18748
rect 37645 18711 37703 18717
rect 38286 18708 38292 18720
rect 38344 18708 38350 18760
rect 15528 18652 15573 18680
rect 15672 18652 17080 18680
rect 15528 18640 15534 18652
rect 15672 18612 15700 18652
rect 17218 18640 17224 18692
rect 17276 18680 17282 18692
rect 23385 18683 23443 18689
rect 23385 18680 23397 18683
rect 17276 18652 23397 18680
rect 17276 18640 17282 18652
rect 23385 18649 23397 18652
rect 23431 18649 23443 18683
rect 23385 18643 23443 18649
rect 23474 18640 23480 18692
rect 23532 18680 23538 18692
rect 24029 18683 24087 18689
rect 23532 18652 23577 18680
rect 23532 18640 23538 18652
rect 24029 18649 24041 18683
rect 24075 18649 24087 18683
rect 24029 18643 24087 18649
rect 24765 18683 24823 18689
rect 24765 18649 24777 18683
rect 24811 18680 24823 18683
rect 24854 18680 24860 18692
rect 24811 18652 24860 18680
rect 24811 18649 24823 18652
rect 24765 18643 24823 18649
rect 17034 18612 17040 18624
rect 14568 18584 15700 18612
rect 16995 18584 17040 18612
rect 17034 18572 17040 18584
rect 17092 18572 17098 18624
rect 17402 18572 17408 18624
rect 17460 18612 17466 18624
rect 18325 18615 18383 18621
rect 18325 18612 18337 18615
rect 17460 18584 18337 18612
rect 17460 18572 17466 18584
rect 18325 18581 18337 18584
rect 18371 18581 18383 18615
rect 18325 18575 18383 18581
rect 18414 18572 18420 18624
rect 18472 18612 18478 18624
rect 23934 18612 23940 18624
rect 18472 18584 23940 18612
rect 18472 18572 18478 18584
rect 23934 18572 23940 18584
rect 23992 18572 23998 18624
rect 24044 18612 24072 18643
rect 24854 18640 24860 18652
rect 24912 18640 24918 18692
rect 25317 18683 25375 18689
rect 25317 18649 25329 18683
rect 25363 18680 25375 18683
rect 34514 18680 34520 18692
rect 25363 18652 34520 18680
rect 25363 18649 25375 18652
rect 25317 18643 25375 18649
rect 25332 18612 25360 18643
rect 34514 18640 34520 18652
rect 34572 18640 34578 18692
rect 24044 18584 25360 18612
rect 26881 18615 26939 18621
rect 26881 18581 26893 18615
rect 26927 18612 26939 18615
rect 27338 18612 27344 18624
rect 26927 18584 27344 18612
rect 26927 18581 26939 18584
rect 26881 18575 26939 18581
rect 27338 18572 27344 18584
rect 27396 18572 27402 18624
rect 38102 18612 38108 18624
rect 38063 18584 38108 18612
rect 38102 18572 38108 18584
rect 38160 18572 38166 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 1670 18368 1676 18420
rect 1728 18408 1734 18420
rect 2041 18411 2099 18417
rect 2041 18408 2053 18411
rect 1728 18380 2053 18408
rect 1728 18368 1734 18380
rect 2041 18377 2053 18380
rect 2087 18377 2099 18411
rect 4706 18408 4712 18420
rect 2041 18371 2099 18377
rect 2792 18380 4712 18408
rect 2792 18349 2820 18380
rect 4706 18368 4712 18380
rect 4764 18368 4770 18420
rect 5258 18368 5264 18420
rect 5316 18408 5322 18420
rect 5316 18380 6868 18408
rect 5316 18368 5322 18380
rect 2777 18343 2835 18349
rect 2777 18309 2789 18343
rect 2823 18309 2835 18343
rect 2777 18303 2835 18309
rect 3329 18343 3387 18349
rect 3329 18309 3341 18343
rect 3375 18340 3387 18343
rect 3970 18340 3976 18352
rect 3375 18312 3976 18340
rect 3375 18309 3387 18312
rect 3329 18303 3387 18309
rect 3970 18300 3976 18312
rect 4028 18300 4034 18352
rect 4065 18343 4123 18349
rect 4065 18309 4077 18343
rect 4111 18340 4123 18343
rect 5166 18340 5172 18352
rect 4111 18312 5172 18340
rect 4111 18309 4123 18312
rect 4065 18303 4123 18309
rect 5166 18300 5172 18312
rect 5224 18300 5230 18352
rect 6733 18343 6791 18349
rect 6733 18340 6745 18343
rect 5828 18312 6745 18340
rect 1854 18272 1860 18284
rect 1815 18244 1860 18272
rect 1854 18232 1860 18244
rect 1912 18232 1918 18284
rect 5074 18272 5080 18284
rect 5035 18244 5080 18272
rect 5074 18232 5080 18244
rect 5132 18232 5138 18284
rect 2685 18207 2743 18213
rect 2685 18173 2697 18207
rect 2731 18204 2743 18207
rect 3326 18204 3332 18216
rect 2731 18176 3332 18204
rect 2731 18173 2743 18176
rect 2685 18167 2743 18173
rect 3326 18164 3332 18176
rect 3384 18164 3390 18216
rect 3973 18207 4031 18213
rect 3973 18173 3985 18207
rect 4019 18204 4031 18207
rect 4062 18204 4068 18216
rect 4019 18176 4068 18204
rect 4019 18173 4031 18176
rect 3973 18167 4031 18173
rect 2958 18096 2964 18148
rect 3016 18136 3022 18148
rect 3988 18136 4016 18167
rect 4062 18164 4068 18176
rect 4120 18164 4126 18216
rect 4617 18207 4675 18213
rect 4617 18173 4629 18207
rect 4663 18204 4675 18207
rect 5718 18204 5724 18216
rect 4663 18176 5724 18204
rect 4663 18173 4675 18176
rect 4617 18167 4675 18173
rect 5718 18164 5724 18176
rect 5776 18164 5782 18216
rect 5828 18136 5856 18312
rect 6733 18309 6745 18312
rect 6779 18309 6791 18343
rect 6840 18340 6868 18380
rect 6914 18368 6920 18420
rect 6972 18408 6978 18420
rect 8754 18408 8760 18420
rect 6972 18380 8760 18408
rect 6972 18368 6978 18380
rect 8754 18368 8760 18380
rect 8812 18368 8818 18420
rect 15470 18368 15476 18420
rect 15528 18408 15534 18420
rect 16945 18411 17003 18417
rect 16945 18408 16957 18411
rect 15528 18380 16957 18408
rect 15528 18368 15534 18380
rect 16945 18377 16957 18380
rect 16991 18377 17003 18411
rect 16945 18371 17003 18377
rect 19978 18368 19984 18420
rect 20036 18408 20042 18420
rect 20533 18411 20591 18417
rect 20533 18408 20545 18411
rect 20036 18380 20545 18408
rect 20036 18368 20042 18380
rect 20533 18377 20545 18380
rect 20579 18377 20591 18411
rect 36354 18408 36360 18420
rect 20533 18371 20591 18377
rect 22066 18380 36360 18408
rect 10606 18343 10664 18349
rect 6840 18312 8602 18340
rect 6733 18303 6791 18309
rect 10606 18309 10618 18343
rect 10652 18340 10664 18343
rect 10870 18340 10876 18352
rect 10652 18312 10876 18340
rect 10652 18309 10664 18312
rect 10606 18303 10664 18309
rect 10870 18300 10876 18312
rect 10928 18300 10934 18352
rect 11882 18340 11888 18352
rect 11843 18312 11888 18340
rect 11882 18300 11888 18312
rect 11940 18300 11946 18352
rect 11977 18343 12035 18349
rect 11977 18309 11989 18343
rect 12023 18340 12035 18343
rect 12986 18340 12992 18352
rect 12023 18312 12992 18340
rect 12023 18309 12035 18312
rect 11977 18303 12035 18309
rect 12986 18300 12992 18312
rect 13044 18300 13050 18352
rect 13538 18340 13544 18352
rect 13499 18312 13544 18340
rect 13538 18300 13544 18312
rect 13596 18300 13602 18352
rect 13630 18300 13636 18352
rect 13688 18340 13694 18352
rect 13688 18312 15700 18340
rect 13688 18300 13694 18312
rect 10318 18232 10324 18284
rect 10376 18232 10382 18284
rect 15013 18275 15071 18281
rect 15013 18241 15025 18275
rect 15059 18241 15071 18275
rect 15194 18272 15200 18284
rect 15155 18244 15200 18272
rect 15013 18235 15071 18241
rect 5905 18207 5963 18213
rect 5905 18173 5917 18207
rect 5951 18173 5963 18207
rect 6638 18204 6644 18216
rect 6599 18176 6644 18204
rect 5905 18167 5963 18173
rect 3016 18108 4016 18136
rect 4080 18108 5856 18136
rect 5920 18136 5948 18167
rect 6638 18164 6644 18176
rect 6696 18164 6702 18216
rect 7837 18207 7895 18213
rect 7837 18204 7849 18207
rect 6748 18176 7849 18204
rect 6546 18136 6552 18148
rect 5920 18108 6552 18136
rect 3016 18096 3022 18108
rect 1762 18028 1768 18080
rect 1820 18068 1826 18080
rect 4080 18068 4108 18108
rect 6546 18096 6552 18108
rect 6604 18136 6610 18148
rect 6748 18136 6776 18176
rect 7837 18173 7849 18176
rect 7883 18173 7895 18207
rect 8113 18207 8171 18213
rect 8113 18204 8125 18207
rect 7837 18167 7895 18173
rect 7944 18176 8125 18204
rect 6604 18108 6776 18136
rect 7193 18139 7251 18145
rect 6604 18096 6610 18108
rect 7193 18105 7205 18139
rect 7239 18105 7251 18139
rect 7193 18099 7251 18105
rect 1820 18040 4108 18068
rect 1820 18028 1826 18040
rect 4154 18028 4160 18080
rect 4212 18068 4218 18080
rect 4798 18068 4804 18080
rect 4212 18040 4804 18068
rect 4212 18028 4218 18040
rect 4798 18028 4804 18040
rect 4856 18068 4862 18080
rect 7208 18068 7236 18099
rect 7742 18096 7748 18148
rect 7800 18136 7806 18148
rect 7944 18136 7972 18176
rect 8113 18173 8125 18176
rect 8159 18173 8171 18207
rect 8113 18167 8171 18173
rect 8662 18164 8668 18216
rect 8720 18204 8726 18216
rect 10042 18204 10048 18216
rect 8720 18176 10048 18204
rect 8720 18164 8726 18176
rect 10042 18164 10048 18176
rect 10100 18164 10106 18216
rect 10336 18204 10364 18232
rect 10505 18207 10563 18213
rect 10505 18204 10517 18207
rect 10336 18176 10517 18204
rect 10505 18173 10517 18176
rect 10551 18173 10563 18207
rect 10505 18167 10563 18173
rect 12897 18207 12955 18213
rect 12897 18173 12909 18207
rect 12943 18204 12955 18207
rect 13078 18204 13084 18216
rect 12943 18176 13084 18204
rect 12943 18173 12955 18176
rect 12897 18167 12955 18173
rect 13078 18164 13084 18176
rect 13136 18164 13142 18216
rect 13449 18207 13507 18213
rect 13449 18173 13461 18207
rect 13495 18173 13507 18207
rect 14366 18204 14372 18216
rect 14327 18176 14372 18204
rect 13449 18167 13507 18173
rect 7800 18108 7972 18136
rect 7800 18096 7806 18108
rect 9674 18096 9680 18148
rect 9732 18136 9738 18148
rect 10962 18136 10968 18148
rect 9732 18108 10968 18136
rect 9732 18096 9738 18108
rect 10962 18096 10968 18108
rect 11020 18136 11026 18148
rect 11057 18139 11115 18145
rect 11057 18136 11069 18139
rect 11020 18108 11069 18136
rect 11020 18096 11026 18108
rect 11057 18105 11069 18108
rect 11103 18105 11115 18139
rect 11057 18099 11115 18105
rect 11422 18096 11428 18148
rect 11480 18136 11486 18148
rect 11606 18136 11612 18148
rect 11480 18108 11612 18136
rect 11480 18096 11486 18108
rect 11606 18096 11612 18108
rect 11664 18096 11670 18148
rect 13354 18096 13360 18148
rect 13412 18136 13418 18148
rect 13464 18136 13492 18167
rect 14366 18164 14372 18176
rect 14424 18204 14430 18216
rect 14826 18204 14832 18216
rect 14424 18176 14832 18204
rect 14424 18164 14430 18176
rect 14826 18164 14832 18176
rect 14884 18164 14890 18216
rect 15028 18204 15056 18235
rect 15194 18232 15200 18244
rect 15252 18232 15258 18284
rect 15672 18281 15700 18312
rect 16206 18300 16212 18352
rect 16264 18340 16270 18352
rect 17034 18340 17040 18352
rect 16264 18312 17040 18340
rect 16264 18300 16270 18312
rect 17034 18300 17040 18312
rect 17092 18300 17098 18352
rect 22066 18340 22094 18380
rect 36354 18368 36360 18380
rect 36412 18368 36418 18420
rect 38010 18368 38016 18420
rect 38068 18408 38074 18420
rect 38105 18411 38163 18417
rect 38105 18408 38117 18411
rect 38068 18380 38117 18408
rect 38068 18368 38074 18380
rect 38105 18377 38117 18380
rect 38151 18377 38163 18411
rect 38105 18371 38163 18377
rect 17512 18312 22094 18340
rect 22189 18343 22247 18349
rect 15657 18275 15715 18281
rect 15657 18241 15669 18275
rect 15703 18272 15715 18275
rect 16482 18272 16488 18284
rect 15703 18244 16488 18272
rect 15703 18241 15715 18244
rect 15657 18235 15715 18241
rect 16482 18232 16488 18244
rect 16540 18232 16546 18284
rect 16574 18232 16580 18284
rect 16632 18272 16638 18284
rect 17512 18281 17540 18312
rect 22189 18309 22201 18343
rect 22235 18340 22247 18343
rect 22278 18340 22284 18352
rect 22235 18312 22284 18340
rect 22235 18309 22247 18312
rect 22189 18303 22247 18309
rect 22278 18300 22284 18312
rect 22336 18300 22342 18352
rect 23109 18343 23167 18349
rect 23109 18309 23121 18343
rect 23155 18340 23167 18343
rect 23198 18340 23204 18352
rect 23155 18312 23204 18340
rect 23155 18309 23167 18312
rect 23109 18303 23167 18309
rect 16853 18275 16911 18281
rect 16853 18272 16865 18275
rect 16632 18244 16865 18272
rect 16632 18232 16638 18244
rect 16853 18241 16865 18244
rect 16899 18241 16911 18275
rect 16853 18235 16911 18241
rect 17497 18275 17555 18281
rect 17497 18241 17509 18275
rect 17543 18241 17555 18275
rect 17497 18235 17555 18241
rect 17512 18204 17540 18235
rect 20070 18232 20076 18284
rect 20128 18272 20134 18284
rect 20441 18275 20499 18281
rect 20441 18272 20453 18275
rect 20128 18244 20453 18272
rect 20128 18232 20134 18244
rect 20441 18241 20453 18244
rect 20487 18241 20499 18275
rect 20441 18235 20499 18241
rect 15028 18176 17540 18204
rect 22094 18164 22100 18216
rect 22152 18204 22158 18216
rect 22152 18176 22197 18204
rect 22152 18164 22158 18176
rect 17589 18139 17647 18145
rect 17589 18136 17601 18139
rect 13412 18108 17601 18136
rect 13412 18096 13418 18108
rect 17589 18105 17601 18108
rect 17635 18105 17647 18139
rect 17589 18099 17647 18105
rect 21450 18096 21456 18148
rect 21508 18136 21514 18148
rect 23124 18136 23152 18303
rect 23198 18300 23204 18312
rect 23256 18300 23262 18352
rect 23845 18343 23903 18349
rect 23845 18309 23857 18343
rect 23891 18340 23903 18343
rect 24949 18343 25007 18349
rect 24949 18340 24961 18343
rect 23891 18312 24961 18340
rect 23891 18309 23903 18312
rect 23845 18303 23903 18309
rect 24949 18309 24961 18312
rect 24995 18309 25007 18343
rect 24949 18303 25007 18309
rect 27246 18300 27252 18352
rect 27304 18340 27310 18352
rect 27801 18343 27859 18349
rect 27801 18340 27813 18343
rect 27304 18312 27813 18340
rect 27304 18300 27310 18312
rect 27801 18309 27813 18312
rect 27847 18309 27859 18343
rect 27801 18303 27859 18309
rect 24857 18275 24915 18281
rect 24857 18241 24869 18275
rect 24903 18272 24915 18275
rect 25130 18272 25136 18284
rect 24903 18244 25136 18272
rect 24903 18241 24915 18244
rect 24857 18235 24915 18241
rect 25130 18232 25136 18244
rect 25188 18232 25194 18284
rect 27338 18272 27344 18284
rect 27299 18244 27344 18272
rect 27338 18232 27344 18244
rect 27396 18232 27402 18284
rect 31481 18275 31539 18281
rect 31481 18241 31493 18275
rect 31527 18272 31539 18275
rect 38102 18272 38108 18284
rect 31527 18244 38108 18272
rect 31527 18241 31539 18244
rect 31481 18235 31539 18241
rect 38102 18232 38108 18244
rect 38160 18232 38166 18284
rect 38286 18272 38292 18284
rect 38247 18244 38292 18272
rect 38286 18232 38292 18244
rect 38344 18232 38350 18284
rect 23750 18204 23756 18216
rect 23711 18176 23756 18204
rect 23750 18164 23756 18176
rect 23808 18164 23814 18216
rect 24397 18207 24455 18213
rect 24397 18173 24409 18207
rect 24443 18204 24455 18207
rect 24946 18204 24952 18216
rect 24443 18176 24952 18204
rect 24443 18173 24455 18176
rect 24397 18167 24455 18173
rect 21508 18108 23152 18136
rect 21508 18096 21514 18108
rect 4856 18040 7236 18068
rect 4856 18028 4862 18040
rect 7466 18028 7472 18080
rect 7524 18068 7530 18080
rect 9585 18071 9643 18077
rect 9585 18068 9597 18071
rect 7524 18040 9597 18068
rect 7524 18028 7530 18040
rect 9585 18037 9597 18040
rect 9631 18068 9643 18071
rect 12158 18068 12164 18080
rect 9631 18040 12164 18068
rect 9631 18037 9643 18040
rect 9585 18031 9643 18037
rect 12158 18028 12164 18040
rect 12216 18028 12222 18080
rect 13538 18028 13544 18080
rect 13596 18068 13602 18080
rect 15749 18071 15807 18077
rect 15749 18068 15761 18071
rect 13596 18040 15761 18068
rect 13596 18028 13602 18040
rect 15749 18037 15761 18040
rect 15795 18037 15807 18071
rect 15749 18031 15807 18037
rect 17678 18028 17684 18080
rect 17736 18068 17742 18080
rect 24412 18068 24440 18167
rect 24946 18164 24952 18176
rect 25004 18164 25010 18216
rect 27154 18204 27160 18216
rect 27115 18176 27160 18204
rect 27154 18164 27160 18176
rect 27212 18164 27218 18216
rect 17736 18040 24440 18068
rect 17736 18028 17742 18040
rect 26234 18028 26240 18080
rect 26292 18068 26298 18080
rect 31573 18071 31631 18077
rect 31573 18068 31585 18071
rect 26292 18040 31585 18068
rect 26292 18028 26298 18040
rect 31573 18037 31585 18040
rect 31619 18037 31631 18071
rect 31573 18031 31631 18037
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 3329 17867 3387 17873
rect 3329 17833 3341 17867
rect 3375 17864 3387 17867
rect 4614 17864 4620 17876
rect 3375 17836 4620 17864
rect 3375 17833 3387 17836
rect 3329 17827 3387 17833
rect 4614 17824 4620 17836
rect 4672 17824 4678 17876
rect 4982 17824 4988 17876
rect 5040 17864 5046 17876
rect 5721 17867 5779 17873
rect 5721 17864 5733 17867
rect 5040 17836 5733 17864
rect 5040 17824 5046 17836
rect 5721 17833 5733 17836
rect 5767 17833 5779 17867
rect 11422 17864 11428 17876
rect 5721 17827 5779 17833
rect 6196 17836 11428 17864
rect 6196 17728 6224 17836
rect 11422 17824 11428 17836
rect 11480 17824 11486 17876
rect 12526 17864 12532 17876
rect 11532 17836 12532 17864
rect 8573 17799 8631 17805
rect 8573 17765 8585 17799
rect 8619 17796 8631 17799
rect 8754 17796 8760 17808
rect 8619 17768 8760 17796
rect 8619 17765 8631 17768
rect 8573 17759 8631 17765
rect 8754 17756 8760 17768
rect 8812 17756 8818 17808
rect 10870 17756 10876 17808
rect 10928 17796 10934 17808
rect 11532 17796 11560 17836
rect 12526 17824 12532 17836
rect 12584 17824 12590 17876
rect 12618 17824 12624 17876
rect 12676 17864 12682 17876
rect 18049 17867 18107 17873
rect 18049 17864 18061 17867
rect 12676 17836 18061 17864
rect 12676 17824 12682 17836
rect 18049 17833 18061 17836
rect 18095 17833 18107 17867
rect 20990 17864 20996 17876
rect 18049 17827 18107 17833
rect 19720 17836 20996 17864
rect 14090 17796 14096 17808
rect 10928 17768 11560 17796
rect 13096 17768 14096 17796
rect 10928 17756 10934 17768
rect 2976 17700 6224 17728
rect 6273 17731 6331 17737
rect 1578 17660 1584 17672
rect 1539 17632 1584 17660
rect 1578 17620 1584 17632
rect 1636 17620 1642 17672
rect 2976 17646 3004 17700
rect 6273 17697 6285 17731
rect 6319 17728 6331 17731
rect 7098 17728 7104 17740
rect 6319 17700 7104 17728
rect 6319 17697 6331 17700
rect 6273 17691 6331 17697
rect 7098 17688 7104 17700
rect 7156 17728 7162 17740
rect 12158 17728 12164 17740
rect 7156 17700 12164 17728
rect 7156 17688 7162 17700
rect 12158 17688 12164 17700
rect 12216 17688 12222 17740
rect 12526 17688 12532 17740
rect 12584 17728 12590 17740
rect 13096 17728 13124 17768
rect 14090 17756 14096 17768
rect 14148 17756 14154 17808
rect 15565 17799 15623 17805
rect 15565 17765 15577 17799
rect 15611 17796 15623 17799
rect 16114 17796 16120 17808
rect 15611 17768 16120 17796
rect 15611 17765 15623 17768
rect 15565 17759 15623 17765
rect 16114 17756 16120 17768
rect 16172 17756 16178 17808
rect 16761 17799 16819 17805
rect 16761 17765 16773 17799
rect 16807 17796 16819 17799
rect 19720 17796 19748 17836
rect 20990 17824 20996 17836
rect 21048 17824 21054 17876
rect 21174 17824 21180 17876
rect 21232 17864 21238 17876
rect 24118 17864 24124 17876
rect 21232 17836 24124 17864
rect 21232 17824 21238 17836
rect 24118 17824 24124 17836
rect 24176 17824 24182 17876
rect 22097 17799 22155 17805
rect 16807 17768 19748 17796
rect 19812 17768 22048 17796
rect 16807 17765 16819 17768
rect 16761 17759 16819 17765
rect 12584 17700 13124 17728
rect 13541 17731 13599 17737
rect 12584 17688 12590 17700
rect 13541 17697 13553 17731
rect 13587 17728 13599 17731
rect 13814 17728 13820 17740
rect 13587 17700 13820 17728
rect 13587 17697 13599 17700
rect 13541 17691 13599 17697
rect 13814 17688 13820 17700
rect 13872 17688 13878 17740
rect 14550 17688 14556 17740
rect 14608 17728 14614 17740
rect 19812 17728 19840 17768
rect 14608 17700 19840 17728
rect 19889 17731 19947 17737
rect 14608 17688 14614 17700
rect 19889 17697 19901 17731
rect 19935 17728 19947 17731
rect 20806 17728 20812 17740
rect 19935 17700 20812 17728
rect 19935 17697 19947 17700
rect 19889 17691 19947 17697
rect 20806 17688 20812 17700
rect 20864 17688 20870 17740
rect 22020 17672 22048 17768
rect 22097 17765 22109 17799
rect 22143 17796 22155 17799
rect 22370 17796 22376 17808
rect 22143 17768 22376 17796
rect 22143 17765 22155 17768
rect 22097 17759 22155 17765
rect 22370 17756 22376 17768
rect 22428 17756 22434 17808
rect 30745 17731 30803 17737
rect 30745 17728 30757 17731
rect 22112 17700 30757 17728
rect 3973 17663 4031 17669
rect 3973 17629 3985 17663
rect 4019 17629 4031 17663
rect 3973 17623 4031 17629
rect 6181 17663 6239 17669
rect 6181 17629 6193 17663
rect 6227 17629 6239 17663
rect 6822 17660 6828 17672
rect 6783 17632 6828 17660
rect 6181 17623 6239 17629
rect 1854 17592 1860 17604
rect 1815 17564 1860 17592
rect 1854 17552 1860 17564
rect 1912 17552 1918 17604
rect 3988 17592 4016 17623
rect 4246 17592 4252 17604
rect 3988 17564 4108 17592
rect 4207 17564 4252 17592
rect 4080 17536 4108 17564
rect 4246 17552 4252 17564
rect 4304 17552 4310 17604
rect 4706 17552 4712 17604
rect 4764 17552 4770 17604
rect 5994 17552 6000 17604
rect 6052 17592 6058 17604
rect 6196 17592 6224 17623
rect 6822 17620 6828 17632
rect 6880 17620 6886 17672
rect 8846 17620 8852 17672
rect 8904 17660 8910 17672
rect 9493 17663 9551 17669
rect 9493 17660 9505 17663
rect 8904 17632 9505 17660
rect 8904 17620 8910 17632
rect 9493 17629 9505 17632
rect 9539 17629 9551 17663
rect 9493 17623 9551 17629
rect 10870 17620 10876 17672
rect 10928 17620 10934 17672
rect 11146 17620 11152 17672
rect 11204 17620 11210 17672
rect 11790 17660 11796 17672
rect 11751 17632 11796 17660
rect 11790 17620 11796 17632
rect 11848 17620 11854 17672
rect 14274 17620 14280 17672
rect 14332 17660 14338 17672
rect 17310 17660 17316 17672
rect 14332 17632 14377 17660
rect 17271 17632 17316 17660
rect 14332 17620 14338 17632
rect 17310 17620 17316 17632
rect 17368 17620 17374 17672
rect 17494 17620 17500 17672
rect 17552 17660 17558 17672
rect 17957 17663 18015 17669
rect 17957 17660 17969 17663
rect 17552 17632 17969 17660
rect 17552 17620 17558 17632
rect 17957 17629 17969 17632
rect 18003 17629 18015 17663
rect 22002 17660 22008 17672
rect 21915 17632 22008 17660
rect 17957 17623 18015 17629
rect 22002 17620 22008 17632
rect 22060 17620 22066 17672
rect 6730 17592 6736 17604
rect 6052 17564 6736 17592
rect 6052 17552 6058 17564
rect 6730 17552 6736 17564
rect 6788 17552 6794 17604
rect 7101 17595 7159 17601
rect 7101 17561 7113 17595
rect 7147 17561 7159 17595
rect 7101 17555 7159 17561
rect 4062 17484 4068 17536
rect 4120 17484 4126 17536
rect 7116 17524 7144 17555
rect 7558 17552 7564 17604
rect 7616 17552 7622 17604
rect 9769 17595 9827 17601
rect 8404 17564 9720 17592
rect 8404 17524 8432 17564
rect 7116 17496 8432 17524
rect 9692 17524 9720 17564
rect 9769 17561 9781 17595
rect 9815 17592 9827 17595
rect 10042 17592 10048 17604
rect 9815 17564 10048 17592
rect 9815 17561 9827 17564
rect 9769 17555 9827 17561
rect 10042 17552 10048 17564
rect 10100 17552 10106 17604
rect 11164 17592 11192 17620
rect 12069 17595 12127 17601
rect 12069 17592 12081 17595
rect 11164 17564 12081 17592
rect 12069 17561 12081 17564
rect 12115 17592 12127 17595
rect 12342 17592 12348 17604
rect 12115 17564 12348 17592
rect 12115 17561 12127 17564
rect 12069 17555 12127 17561
rect 12342 17552 12348 17564
rect 12400 17552 12406 17604
rect 13354 17592 13360 17604
rect 13294 17564 13360 17592
rect 13354 17552 13360 17564
rect 13412 17552 13418 17604
rect 15010 17592 15016 17604
rect 14971 17564 15016 17592
rect 15010 17552 15016 17564
rect 15068 17552 15074 17604
rect 15105 17595 15163 17601
rect 15105 17561 15117 17595
rect 15151 17592 15163 17595
rect 16206 17592 16212 17604
rect 15151 17564 15240 17592
rect 16167 17564 16212 17592
rect 15151 17561 15163 17564
rect 15105 17555 15163 17561
rect 10686 17524 10692 17536
rect 9692 17496 10692 17524
rect 10686 17484 10692 17496
rect 10744 17484 10750 17536
rect 11146 17484 11152 17536
rect 11204 17524 11210 17536
rect 11241 17527 11299 17533
rect 11241 17524 11253 17527
rect 11204 17496 11253 17524
rect 11204 17484 11210 17496
rect 11241 17493 11253 17496
rect 11287 17524 11299 17527
rect 13078 17524 13084 17536
rect 11287 17496 13084 17524
rect 11287 17493 11299 17496
rect 11241 17487 11299 17493
rect 13078 17484 13084 17496
rect 13136 17484 13142 17536
rect 13630 17484 13636 17536
rect 13688 17524 13694 17536
rect 14369 17527 14427 17533
rect 14369 17524 14381 17527
rect 13688 17496 14381 17524
rect 13688 17484 13694 17496
rect 14369 17493 14381 17496
rect 14415 17493 14427 17527
rect 15212 17524 15240 17564
rect 16206 17552 16212 17564
rect 16264 17552 16270 17604
rect 16298 17552 16304 17604
rect 16356 17592 16362 17604
rect 16356 17564 16401 17592
rect 16356 17552 16362 17564
rect 17126 17552 17132 17604
rect 17184 17592 17190 17604
rect 17184 17564 17540 17592
rect 17184 17552 17190 17564
rect 17405 17527 17463 17533
rect 17405 17524 17417 17527
rect 15212 17496 17417 17524
rect 14369 17487 14427 17493
rect 17405 17493 17417 17496
rect 17451 17493 17463 17527
rect 17512 17524 17540 17564
rect 17678 17552 17684 17604
rect 17736 17592 17742 17604
rect 19886 17592 19892 17604
rect 17736 17564 19892 17592
rect 17736 17552 17742 17564
rect 19886 17552 19892 17564
rect 19944 17552 19950 17604
rect 19978 17552 19984 17604
rect 20036 17592 20042 17604
rect 20036 17564 20081 17592
rect 20036 17552 20042 17564
rect 20162 17552 20168 17604
rect 20220 17592 20226 17604
rect 20533 17595 20591 17601
rect 20533 17592 20545 17595
rect 20220 17564 20545 17592
rect 20220 17552 20226 17564
rect 20533 17561 20545 17564
rect 20579 17592 20591 17595
rect 20622 17592 20628 17604
rect 20579 17564 20628 17592
rect 20579 17561 20591 17564
rect 20533 17555 20591 17561
rect 20622 17552 20628 17564
rect 20680 17552 20686 17604
rect 22112 17592 22140 17700
rect 30745 17697 30757 17700
rect 30791 17697 30803 17731
rect 30745 17691 30803 17697
rect 22922 17660 22928 17672
rect 22883 17632 22928 17660
rect 22922 17620 22928 17632
rect 22980 17620 22986 17672
rect 28077 17663 28135 17669
rect 28077 17629 28089 17663
rect 28123 17660 28135 17663
rect 28258 17660 28264 17672
rect 28123 17632 28264 17660
rect 28123 17629 28135 17632
rect 28077 17623 28135 17629
rect 28258 17620 28264 17632
rect 28316 17620 28322 17672
rect 28368 17632 35894 17660
rect 22066 17564 22140 17592
rect 23109 17595 23167 17601
rect 22066 17524 22094 17564
rect 23109 17561 23121 17595
rect 23155 17592 23167 17595
rect 28368 17592 28396 17632
rect 30558 17592 30564 17604
rect 23155 17564 28396 17592
rect 30519 17564 30564 17592
rect 23155 17561 23167 17564
rect 23109 17555 23167 17561
rect 30558 17552 30564 17564
rect 30616 17552 30622 17604
rect 17512 17496 22094 17524
rect 17405 17487 17463 17493
rect 27338 17484 27344 17536
rect 27396 17524 27402 17536
rect 27893 17527 27951 17533
rect 27893 17524 27905 17527
rect 27396 17496 27905 17524
rect 27396 17484 27402 17496
rect 27893 17493 27905 17496
rect 27939 17493 27951 17527
rect 35866 17524 35894 17632
rect 37826 17524 37832 17536
rect 35866 17496 37832 17524
rect 27893 17487 27951 17493
rect 37826 17484 37832 17496
rect 37884 17484 37890 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 1946 17280 1952 17332
rect 2004 17320 2010 17332
rect 3694 17320 3700 17332
rect 2004 17292 3556 17320
rect 3655 17292 3700 17320
rect 2004 17280 2010 17292
rect 2866 17212 2872 17264
rect 2924 17212 2930 17264
rect 3528 17252 3556 17292
rect 3694 17280 3700 17292
rect 3752 17280 3758 17332
rect 5997 17323 6055 17329
rect 5997 17320 6009 17323
rect 3804 17292 6009 17320
rect 3804 17252 3832 17292
rect 5997 17289 6009 17292
rect 6043 17320 6055 17323
rect 8478 17320 8484 17332
rect 6043 17292 8484 17320
rect 6043 17289 6055 17292
rect 5997 17283 6055 17289
rect 8478 17280 8484 17292
rect 8536 17280 8542 17332
rect 8662 17280 8668 17332
rect 8720 17320 8726 17332
rect 10042 17320 10048 17332
rect 8720 17292 10048 17320
rect 8720 17280 8726 17292
rect 10042 17280 10048 17292
rect 10100 17280 10106 17332
rect 12158 17280 12164 17332
rect 12216 17320 12222 17332
rect 16206 17320 16212 17332
rect 12216 17292 16212 17320
rect 12216 17280 12222 17292
rect 16206 17280 16212 17292
rect 16264 17280 16270 17332
rect 16482 17280 16488 17332
rect 16540 17320 16546 17332
rect 16666 17320 16672 17332
rect 16540 17292 16672 17320
rect 16540 17280 16546 17292
rect 16666 17280 16672 17292
rect 16724 17280 16730 17332
rect 18417 17323 18475 17329
rect 18417 17289 18429 17323
rect 18463 17320 18475 17323
rect 19978 17320 19984 17332
rect 18463 17292 19984 17320
rect 18463 17289 18475 17292
rect 18417 17283 18475 17289
rect 19978 17280 19984 17292
rect 20036 17280 20042 17332
rect 25041 17323 25099 17329
rect 25041 17289 25053 17323
rect 25087 17320 25099 17323
rect 27154 17320 27160 17332
rect 25087 17292 27160 17320
rect 25087 17289 25099 17292
rect 25041 17283 25099 17289
rect 3528 17224 3832 17252
rect 4525 17255 4583 17261
rect 4525 17221 4537 17255
rect 4571 17252 4583 17255
rect 4614 17252 4620 17264
rect 4571 17224 4620 17252
rect 4571 17221 4583 17224
rect 4525 17215 4583 17221
rect 4614 17212 4620 17224
rect 4672 17212 4678 17264
rect 5534 17212 5540 17264
rect 5592 17212 5598 17264
rect 7834 17212 7840 17264
rect 7892 17212 7898 17264
rect 11054 17252 11060 17264
rect 10350 17224 11060 17252
rect 11054 17212 11060 17224
rect 11112 17212 11118 17264
rect 11146 17212 11152 17264
rect 11204 17252 11210 17264
rect 12250 17252 12256 17264
rect 11204 17224 12256 17252
rect 11204 17212 11210 17224
rect 12250 17212 12256 17224
rect 12308 17212 12314 17264
rect 13814 17212 13820 17264
rect 13872 17252 13878 17264
rect 14550 17252 14556 17264
rect 13872 17224 14556 17252
rect 13872 17212 13878 17224
rect 14550 17212 14556 17224
rect 14608 17212 14614 17264
rect 16850 17252 16856 17264
rect 15778 17224 16856 17252
rect 16850 17212 16856 17224
rect 16908 17212 16914 17264
rect 17770 17252 17776 17264
rect 17420 17224 17776 17252
rect 6546 17184 6552 17196
rect 6507 17156 6552 17184
rect 6546 17144 6552 17156
rect 6604 17144 6610 17196
rect 10594 17144 10600 17196
rect 10652 17184 10658 17196
rect 11790 17184 11796 17196
rect 10652 17156 11796 17184
rect 10652 17144 10658 17156
rect 11790 17144 11796 17156
rect 11848 17184 11854 17196
rect 11977 17187 12035 17193
rect 11977 17184 11989 17187
rect 11848 17156 11989 17184
rect 11848 17144 11854 17156
rect 11977 17153 11989 17156
rect 12023 17153 12035 17187
rect 17037 17187 17095 17193
rect 11977 17147 12035 17153
rect 1578 17076 1584 17128
rect 1636 17116 1642 17128
rect 1949 17119 2007 17125
rect 1949 17116 1961 17119
rect 1636 17088 1961 17116
rect 1636 17076 1642 17088
rect 1949 17085 1961 17088
rect 1995 17085 2007 17119
rect 1949 17079 2007 17085
rect 2225 17119 2283 17125
rect 2225 17085 2237 17119
rect 2271 17116 2283 17119
rect 2271 17088 3924 17116
rect 2271 17085 2283 17088
rect 2225 17079 2283 17085
rect 3896 16980 3924 17088
rect 4062 17076 4068 17128
rect 4120 17116 4126 17128
rect 4249 17119 4307 17125
rect 4249 17116 4261 17119
rect 4120 17088 4261 17116
rect 4120 17076 4126 17088
rect 4249 17085 4261 17088
rect 4295 17085 4307 17119
rect 6825 17119 6883 17125
rect 6825 17116 6837 17119
rect 4249 17079 4307 17085
rect 4356 17088 6837 17116
rect 3970 17008 3976 17060
rect 4028 17048 4034 17060
rect 4356 17048 4384 17088
rect 6825 17085 6837 17088
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 6914 17076 6920 17128
rect 6972 17116 6978 17128
rect 8846 17116 8852 17128
rect 6972 17088 8852 17116
rect 6972 17076 6978 17088
rect 8846 17076 8852 17088
rect 8904 17076 8910 17128
rect 9125 17119 9183 17125
rect 9125 17085 9137 17119
rect 9171 17116 9183 17119
rect 10134 17116 10140 17128
rect 9171 17088 10140 17116
rect 9171 17085 9183 17088
rect 9125 17079 9183 17085
rect 10134 17076 10140 17088
rect 10192 17076 10198 17128
rect 10873 17119 10931 17125
rect 10873 17116 10885 17119
rect 10244 17088 10885 17116
rect 10244 17060 10272 17088
rect 10873 17085 10885 17088
rect 10919 17085 10931 17119
rect 12253 17119 12311 17125
rect 12253 17116 12265 17119
rect 10873 17079 10931 17085
rect 10980 17088 12265 17116
rect 4028 17020 4384 17048
rect 4028 17008 4034 17020
rect 10226 17008 10232 17060
rect 10284 17008 10290 17060
rect 10686 17008 10692 17060
rect 10744 17048 10750 17060
rect 10980 17048 11008 17088
rect 12253 17085 12265 17088
rect 12299 17085 12311 17119
rect 12253 17079 12311 17085
rect 10744 17020 11008 17048
rect 13372 17048 13400 17170
rect 17037 17153 17049 17187
rect 17083 17184 17095 17187
rect 17420 17184 17448 17224
rect 17770 17212 17776 17224
rect 17828 17252 17834 17264
rect 19153 17255 19211 17261
rect 17828 17224 18920 17252
rect 17828 17212 17834 17224
rect 17083 17156 17448 17184
rect 17083 17153 17095 17156
rect 17037 17147 17095 17153
rect 17494 17144 17500 17196
rect 17552 17184 17558 17196
rect 17681 17187 17739 17193
rect 17681 17184 17693 17187
rect 17552 17156 17693 17184
rect 17552 17144 17558 17156
rect 17681 17153 17693 17156
rect 17727 17153 17739 17187
rect 17681 17147 17739 17153
rect 18325 17187 18383 17193
rect 18325 17153 18337 17187
rect 18371 17153 18383 17187
rect 18325 17147 18383 17153
rect 13722 17116 13728 17128
rect 13683 17088 13728 17116
rect 13722 17076 13728 17088
rect 13780 17076 13786 17128
rect 14277 17119 14335 17125
rect 14277 17085 14289 17119
rect 14323 17116 14335 17119
rect 14550 17116 14556 17128
rect 14323 17088 14556 17116
rect 14323 17085 14335 17088
rect 14277 17079 14335 17085
rect 14550 17076 14556 17088
rect 14608 17076 14614 17128
rect 17129 17119 17187 17125
rect 17129 17116 17141 17119
rect 15672 17088 17141 17116
rect 15672 17060 15700 17088
rect 17129 17085 17141 17088
rect 17175 17085 17187 17119
rect 17129 17079 17187 17085
rect 17310 17076 17316 17128
rect 17368 17116 17374 17128
rect 17773 17119 17831 17125
rect 17773 17116 17785 17119
rect 17368 17088 17785 17116
rect 17368 17076 17374 17088
rect 17773 17085 17785 17088
rect 17819 17085 17831 17119
rect 17773 17079 17831 17085
rect 13372 17020 14412 17048
rect 10744 17008 10750 17020
rect 6270 16980 6276 16992
rect 3896 16952 6276 16980
rect 6270 16940 6276 16952
rect 6328 16940 6334 16992
rect 6914 16940 6920 16992
rect 6972 16980 6978 16992
rect 7466 16980 7472 16992
rect 6972 16952 7472 16980
rect 6972 16940 6978 16952
rect 7466 16940 7472 16952
rect 7524 16940 7530 16992
rect 8297 16983 8355 16989
rect 8297 16949 8309 16983
rect 8343 16980 8355 16983
rect 8478 16980 8484 16992
rect 8343 16952 8484 16980
rect 8343 16949 8355 16952
rect 8297 16943 8355 16949
rect 8478 16940 8484 16952
rect 8536 16980 8542 16992
rect 14274 16980 14280 16992
rect 8536 16952 14280 16980
rect 8536 16940 8542 16952
rect 14274 16940 14280 16952
rect 14332 16940 14338 16992
rect 14384 16980 14412 17020
rect 15654 17008 15660 17060
rect 15712 17008 15718 17060
rect 16942 17048 16948 17060
rect 15948 17020 16948 17048
rect 15948 16980 15976 17020
rect 16942 17008 16948 17020
rect 17000 17008 17006 17060
rect 14384 16952 15976 16980
rect 16025 16983 16083 16989
rect 16025 16949 16037 16983
rect 16071 16980 16083 16983
rect 16114 16980 16120 16992
rect 16071 16952 16120 16980
rect 16071 16949 16083 16952
rect 16025 16943 16083 16949
rect 16114 16940 16120 16952
rect 16172 16940 16178 16992
rect 16482 16940 16488 16992
rect 16540 16980 16546 16992
rect 18340 16980 18368 17147
rect 18892 17048 18920 17224
rect 19153 17221 19165 17255
rect 19199 17252 19211 17255
rect 19426 17252 19432 17264
rect 19199 17224 19432 17252
rect 19199 17221 19211 17224
rect 19153 17215 19211 17221
rect 19426 17212 19432 17224
rect 19484 17212 19490 17264
rect 20530 17212 20536 17264
rect 20588 17252 20594 17264
rect 22189 17255 22247 17261
rect 22189 17252 22201 17255
rect 20588 17224 22201 17252
rect 20588 17212 20594 17224
rect 22189 17221 22201 17224
rect 22235 17221 22247 17255
rect 22189 17215 22247 17221
rect 22922 17212 22928 17264
rect 22980 17212 22986 17264
rect 19702 17144 19708 17196
rect 19760 17184 19766 17196
rect 20165 17187 20223 17193
rect 20165 17184 20177 17187
rect 19760 17156 20177 17184
rect 19760 17144 19766 17156
rect 20165 17153 20177 17156
rect 20211 17153 20223 17187
rect 22940 17184 22968 17212
rect 24949 17187 25007 17193
rect 24949 17184 24961 17187
rect 22940 17156 24961 17184
rect 20165 17147 20223 17153
rect 24949 17153 24961 17156
rect 24995 17153 25007 17187
rect 24949 17147 25007 17153
rect 19061 17119 19119 17125
rect 19061 17085 19073 17119
rect 19107 17116 19119 17119
rect 22097 17119 22155 17125
rect 19107 17088 20576 17116
rect 19107 17085 19119 17088
rect 19061 17079 19119 17085
rect 19518 17048 19524 17060
rect 18892 17020 19524 17048
rect 19518 17008 19524 17020
rect 19576 17008 19582 17060
rect 19613 17051 19671 17057
rect 19613 17017 19625 17051
rect 19659 17048 19671 17051
rect 20162 17048 20168 17060
rect 19659 17020 20168 17048
rect 19659 17017 19671 17020
rect 19613 17011 19671 17017
rect 16540 16952 18368 16980
rect 16540 16940 16546 16952
rect 19334 16940 19340 16992
rect 19392 16980 19398 16992
rect 19628 16980 19656 17011
rect 20162 17008 20168 17020
rect 20220 17008 20226 17060
rect 19392 16952 19656 16980
rect 19392 16940 19398 16952
rect 19702 16940 19708 16992
rect 19760 16980 19766 16992
rect 20257 16983 20315 16989
rect 20257 16980 20269 16983
rect 19760 16952 20269 16980
rect 19760 16940 19766 16952
rect 20257 16949 20269 16952
rect 20303 16949 20315 16983
rect 20548 16980 20576 17088
rect 22097 17085 22109 17119
rect 22143 17085 22155 17119
rect 22370 17116 22376 17128
rect 22331 17088 22376 17116
rect 22097 17079 22155 17085
rect 22112 17048 22140 17079
rect 22370 17076 22376 17088
rect 22428 17076 22434 17128
rect 25056 17048 25084 17283
rect 27154 17280 27160 17292
rect 27212 17280 27218 17332
rect 28258 17320 28264 17332
rect 28219 17292 28264 17320
rect 28258 17280 28264 17292
rect 28316 17280 28322 17332
rect 27338 17184 27344 17196
rect 27299 17156 27344 17184
rect 27338 17144 27344 17156
rect 27396 17144 27402 17196
rect 28442 17184 28448 17196
rect 28403 17156 28448 17184
rect 28442 17144 28448 17156
rect 28500 17144 28506 17196
rect 27157 17119 27215 17125
rect 27157 17085 27169 17119
rect 27203 17116 27215 17119
rect 27246 17116 27252 17128
rect 27203 17088 27252 17116
rect 27203 17085 27215 17088
rect 27157 17079 27215 17085
rect 27246 17076 27252 17088
rect 27304 17076 27310 17128
rect 22112 17020 25084 17048
rect 24394 16980 24400 16992
rect 20548 16952 24400 16980
rect 20257 16943 20315 16949
rect 24394 16940 24400 16952
rect 24452 16940 24458 16992
rect 27614 16980 27620 16992
rect 27575 16952 27620 16980
rect 27614 16940 27620 16952
rect 27672 16940 27678 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 3234 16736 3240 16788
rect 3292 16776 3298 16788
rect 3970 16776 3976 16788
rect 3292 16748 3976 16776
rect 3292 16736 3298 16748
rect 3970 16736 3976 16748
rect 4028 16736 4034 16788
rect 4880 16779 4938 16785
rect 4880 16745 4892 16779
rect 4926 16776 4938 16779
rect 4982 16776 4988 16788
rect 4926 16748 4988 16776
rect 4926 16745 4938 16748
rect 4880 16739 4938 16745
rect 4982 16736 4988 16748
rect 5040 16736 5046 16788
rect 7742 16736 7748 16788
rect 7800 16776 7806 16788
rect 8662 16776 8668 16788
rect 7800 16748 8668 16776
rect 7800 16736 7806 16748
rect 8662 16736 8668 16748
rect 8720 16736 8726 16788
rect 8772 16748 12572 16776
rect 1857 16643 1915 16649
rect 1857 16609 1869 16643
rect 1903 16640 1915 16643
rect 3418 16640 3424 16652
rect 1903 16612 3424 16640
rect 1903 16609 1915 16612
rect 1857 16603 1915 16609
rect 3418 16600 3424 16612
rect 3476 16600 3482 16652
rect 4246 16600 4252 16652
rect 4304 16640 4310 16652
rect 4617 16643 4675 16649
rect 4617 16640 4629 16643
rect 4304 16612 4629 16640
rect 4304 16600 4310 16612
rect 4617 16609 4629 16612
rect 4663 16640 4675 16643
rect 6546 16640 6552 16652
rect 4663 16612 6552 16640
rect 4663 16609 4675 16612
rect 4617 16603 4675 16609
rect 6546 16600 6552 16612
rect 6604 16600 6610 16652
rect 7101 16643 7159 16649
rect 7101 16609 7113 16643
rect 7147 16640 7159 16643
rect 8772 16640 8800 16748
rect 9214 16668 9220 16720
rect 9272 16708 9278 16720
rect 9398 16708 9404 16720
rect 9272 16680 9404 16708
rect 9272 16668 9278 16680
rect 9398 16668 9404 16680
rect 9456 16708 9462 16720
rect 10686 16708 10692 16720
rect 9456 16680 10692 16708
rect 9456 16668 9462 16680
rect 10686 16668 10692 16680
rect 10744 16668 10750 16720
rect 12066 16668 12072 16720
rect 12124 16708 12130 16720
rect 12544 16708 12572 16748
rect 13170 16736 13176 16788
rect 13228 16776 13234 16788
rect 13722 16776 13728 16788
rect 13228 16748 13728 16776
rect 13228 16736 13234 16748
rect 13722 16736 13728 16748
rect 13780 16736 13786 16788
rect 15010 16736 15016 16788
rect 15068 16776 15074 16788
rect 15654 16776 15660 16788
rect 15068 16748 15660 16776
rect 15068 16736 15074 16748
rect 15654 16736 15660 16748
rect 15712 16736 15718 16788
rect 16298 16736 16304 16788
rect 16356 16776 16362 16788
rect 18693 16779 18751 16785
rect 18693 16776 18705 16779
rect 16356 16748 18705 16776
rect 16356 16736 16362 16748
rect 18693 16745 18705 16748
rect 18739 16745 18751 16779
rect 22370 16776 22376 16788
rect 18693 16739 18751 16745
rect 18800 16748 22376 16776
rect 14090 16708 14096 16720
rect 12124 16680 12388 16708
rect 12544 16680 14096 16708
rect 12124 16668 12130 16680
rect 7147 16612 8800 16640
rect 7147 16609 7159 16612
rect 7101 16603 7159 16609
rect 8846 16600 8852 16652
rect 8904 16640 8910 16652
rect 9861 16643 9919 16649
rect 9861 16640 9873 16643
rect 8904 16612 9873 16640
rect 8904 16600 8910 16612
rect 9861 16609 9873 16612
rect 9907 16609 9919 16643
rect 9861 16603 9919 16609
rect 10965 16643 11023 16649
rect 10965 16609 10977 16643
rect 11011 16640 11023 16643
rect 11330 16640 11336 16652
rect 11011 16612 11336 16640
rect 11011 16609 11023 16612
rect 10965 16603 11023 16609
rect 11330 16600 11336 16612
rect 11388 16640 11394 16652
rect 12360 16640 12388 16680
rect 14090 16668 14096 16680
rect 14148 16668 14154 16720
rect 17862 16668 17868 16720
rect 17920 16708 17926 16720
rect 18800 16708 18828 16748
rect 22370 16736 22376 16748
rect 22428 16736 22434 16788
rect 17920 16680 18828 16708
rect 17920 16668 17926 16680
rect 18966 16668 18972 16720
rect 19024 16708 19030 16720
rect 19024 16680 20208 16708
rect 19024 16668 19030 16680
rect 20180 16652 20208 16680
rect 14550 16640 14556 16652
rect 11388 16612 12296 16640
rect 12360 16612 13584 16640
rect 11388 16600 11394 16612
rect 1578 16572 1584 16584
rect 1539 16544 1584 16572
rect 1578 16532 1584 16544
rect 1636 16532 1642 16584
rect 3973 16575 4031 16581
rect 3973 16541 3985 16575
rect 4019 16572 4031 16575
rect 4522 16572 4528 16584
rect 4019 16544 4528 16572
rect 4019 16541 4031 16544
rect 3973 16535 4031 16541
rect 4522 16532 4528 16544
rect 4580 16532 4586 16584
rect 6822 16572 6828 16584
rect 6783 16544 6828 16572
rect 6822 16532 6828 16544
rect 6880 16532 6886 16584
rect 9306 16532 9312 16584
rect 9364 16572 9370 16584
rect 9364 16544 10549 16572
rect 9364 16532 9370 16544
rect 3786 16504 3792 16516
rect 3082 16476 3792 16504
rect 3786 16464 3792 16476
rect 3844 16464 3850 16516
rect 4614 16504 4620 16516
rect 3988 16476 4620 16504
rect 3329 16439 3387 16445
rect 3329 16405 3341 16439
rect 3375 16436 3387 16439
rect 3988 16436 4016 16476
rect 4614 16464 4620 16476
rect 4672 16464 4678 16516
rect 5626 16464 5632 16516
rect 5684 16464 5690 16516
rect 6196 16476 7512 16504
rect 3375 16408 4016 16436
rect 3375 16405 3387 16408
rect 3329 16399 3387 16405
rect 4062 16396 4068 16448
rect 4120 16436 4126 16448
rect 4120 16408 4165 16436
rect 4120 16396 4126 16408
rect 5074 16396 5080 16448
rect 5132 16436 5138 16448
rect 6196 16436 6224 16476
rect 6362 16436 6368 16448
rect 5132 16408 6224 16436
rect 6323 16408 6368 16436
rect 5132 16396 5138 16408
rect 6362 16396 6368 16408
rect 6420 16396 6426 16448
rect 7484 16436 7512 16476
rect 7650 16464 7656 16516
rect 7708 16464 7714 16516
rect 9125 16507 9183 16513
rect 9125 16504 9137 16507
rect 8396 16476 9137 16504
rect 8396 16436 8424 16476
rect 9125 16473 9137 16476
rect 9171 16504 9183 16507
rect 9674 16504 9680 16516
rect 9171 16476 9680 16504
rect 9171 16473 9183 16476
rect 9125 16467 9183 16473
rect 9674 16464 9680 16476
rect 9732 16464 9738 16516
rect 10521 16504 10549 16544
rect 10594 16532 10600 16584
rect 10652 16572 10658 16584
rect 10689 16575 10747 16581
rect 10689 16572 10701 16575
rect 10652 16544 10701 16572
rect 10652 16532 10658 16544
rect 10689 16541 10701 16544
rect 10735 16541 10747 16575
rect 12268 16572 12296 16612
rect 12434 16572 12440 16584
rect 12268 16544 12440 16572
rect 10689 16535 10747 16541
rect 12434 16532 12440 16544
rect 12492 16532 12498 16584
rect 13556 16581 13584 16612
rect 14292 16612 14556 16640
rect 14292 16584 14320 16612
rect 14550 16600 14556 16612
rect 14608 16600 14614 16652
rect 15746 16600 15752 16652
rect 15804 16640 15810 16652
rect 15930 16640 15936 16652
rect 15804 16612 15936 16640
rect 15804 16600 15810 16612
rect 15930 16600 15936 16612
rect 15988 16600 15994 16652
rect 19521 16643 19579 16649
rect 19521 16609 19533 16643
rect 19567 16640 19579 16643
rect 20070 16640 20076 16652
rect 19567 16612 20076 16640
rect 19567 16609 19579 16612
rect 19521 16603 19579 16609
rect 20070 16600 20076 16612
rect 20128 16600 20134 16652
rect 20162 16600 20168 16652
rect 20220 16600 20226 16652
rect 20438 16600 20444 16652
rect 20496 16640 20502 16652
rect 20714 16640 20720 16652
rect 20496 16612 20720 16640
rect 20496 16600 20502 16612
rect 20714 16600 20720 16612
rect 20772 16600 20778 16652
rect 22002 16600 22008 16652
rect 22060 16640 22066 16652
rect 24578 16640 24584 16652
rect 22060 16612 22508 16640
rect 24539 16612 24584 16640
rect 22060 16600 22066 16612
rect 13541 16575 13599 16581
rect 13541 16541 13553 16575
rect 13587 16541 13599 16575
rect 14274 16572 14280 16584
rect 14235 16544 14280 16572
rect 13541 16535 13599 16541
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 16206 16572 16212 16584
rect 15686 16544 16212 16572
rect 16206 16532 16212 16544
rect 16264 16532 16270 16584
rect 16666 16532 16672 16584
rect 16724 16572 16730 16584
rect 16853 16575 16911 16581
rect 16853 16572 16865 16575
rect 16724 16544 16865 16572
rect 16724 16532 16730 16544
rect 16853 16541 16865 16544
rect 16899 16541 16911 16575
rect 16853 16535 16911 16541
rect 16942 16532 16948 16584
rect 17000 16572 17006 16584
rect 17494 16572 17500 16584
rect 17000 16544 17045 16572
rect 17455 16544 17500 16572
rect 17000 16532 17006 16544
rect 17494 16532 17500 16544
rect 17552 16572 17558 16584
rect 18598 16572 18604 16584
rect 17552 16544 18604 16572
rect 17552 16532 17558 16544
rect 18598 16532 18604 16544
rect 18656 16532 18662 16584
rect 18877 16575 18935 16581
rect 18877 16541 18889 16575
rect 18923 16572 18935 16575
rect 19334 16572 19340 16584
rect 18923 16544 19340 16572
rect 18923 16541 18935 16544
rect 18877 16535 18935 16541
rect 19334 16532 19340 16544
rect 19392 16532 19398 16584
rect 22480 16581 22508 16612
rect 24578 16600 24584 16612
rect 24636 16600 24642 16652
rect 24765 16643 24823 16649
rect 24765 16609 24777 16643
rect 24811 16640 24823 16643
rect 26142 16640 26148 16652
rect 24811 16612 26148 16640
rect 24811 16609 24823 16612
rect 24765 16603 24823 16609
rect 26142 16600 26148 16612
rect 26200 16600 26206 16652
rect 22465 16575 22523 16581
rect 22465 16541 22477 16575
rect 22511 16541 22523 16575
rect 22465 16535 22523 16541
rect 25225 16575 25283 16581
rect 25225 16541 25237 16575
rect 25271 16572 25283 16575
rect 27614 16572 27620 16584
rect 25271 16544 27620 16572
rect 25271 16541 25283 16544
rect 25225 16535 25283 16541
rect 27614 16532 27620 16544
rect 27672 16532 27678 16584
rect 38010 16572 38016 16584
rect 37971 16544 38016 16572
rect 38010 16532 38016 16544
rect 38068 16532 38074 16584
rect 10962 16504 10968 16516
rect 10521 16476 10968 16504
rect 10962 16464 10968 16476
rect 11020 16464 11026 16516
rect 12250 16504 12256 16516
rect 12190 16476 12256 16504
rect 12250 16464 12256 16476
rect 12308 16464 12314 16516
rect 12802 16464 12808 16516
rect 12860 16504 12866 16516
rect 13633 16507 13691 16513
rect 13633 16504 13645 16507
rect 12860 16476 13645 16504
rect 12860 16464 12866 16476
rect 13633 16473 13645 16476
rect 13679 16473 13691 16507
rect 13633 16467 13691 16473
rect 14553 16507 14611 16513
rect 14553 16473 14565 16507
rect 14599 16504 14611 16507
rect 14642 16504 14648 16516
rect 14599 16476 14648 16504
rect 14599 16473 14611 16476
rect 14553 16467 14611 16473
rect 14642 16464 14648 16476
rect 14700 16464 14706 16516
rect 16298 16464 16304 16516
rect 16356 16504 16362 16516
rect 17589 16507 17647 16513
rect 17589 16504 17601 16507
rect 16356 16476 17601 16504
rect 16356 16464 16362 16476
rect 17589 16473 17601 16476
rect 17635 16473 17647 16507
rect 17589 16467 17647 16473
rect 19606 16507 19664 16513
rect 19606 16473 19618 16507
rect 19652 16504 19664 16507
rect 19702 16504 19708 16516
rect 19652 16476 19708 16504
rect 19652 16473 19664 16476
rect 19606 16467 19664 16473
rect 19702 16464 19708 16476
rect 19760 16464 19766 16516
rect 20438 16464 20444 16516
rect 20496 16504 20502 16516
rect 20533 16507 20591 16513
rect 20533 16504 20545 16507
rect 20496 16476 20545 16504
rect 20496 16464 20502 16476
rect 20533 16473 20545 16476
rect 20579 16473 20591 16507
rect 28626 16504 28632 16516
rect 20533 16467 20591 16473
rect 22066 16476 28632 16504
rect 7484 16408 8424 16436
rect 8570 16396 8576 16448
rect 8628 16436 8634 16448
rect 9692 16436 9720 16464
rect 11054 16436 11060 16448
rect 8628 16408 8673 16436
rect 9692 16408 11060 16436
rect 8628 16396 8634 16408
rect 11054 16396 11060 16408
rect 11112 16396 11118 16448
rect 11146 16396 11152 16448
rect 11204 16436 11210 16448
rect 11974 16436 11980 16448
rect 11204 16408 11980 16436
rect 11204 16396 11210 16408
rect 11974 16396 11980 16408
rect 12032 16396 12038 16448
rect 12437 16439 12495 16445
rect 12437 16405 12449 16439
rect 12483 16436 12495 16439
rect 12526 16436 12532 16448
rect 12483 16408 12532 16436
rect 12483 16405 12495 16408
rect 12437 16399 12495 16405
rect 12526 16396 12532 16408
rect 12584 16396 12590 16448
rect 15930 16396 15936 16448
rect 15988 16436 15994 16448
rect 16025 16439 16083 16445
rect 16025 16436 16037 16439
rect 15988 16408 16037 16436
rect 15988 16396 15994 16408
rect 16025 16405 16037 16408
rect 16071 16436 16083 16439
rect 18690 16436 18696 16448
rect 16071 16408 18696 16436
rect 16071 16405 16083 16408
rect 16025 16399 16083 16405
rect 18690 16396 18696 16408
rect 18748 16396 18754 16448
rect 19518 16396 19524 16448
rect 19576 16436 19582 16448
rect 22066 16436 22094 16476
rect 28626 16464 28632 16476
rect 28684 16464 28690 16516
rect 22554 16436 22560 16448
rect 19576 16408 22094 16436
rect 22515 16408 22560 16436
rect 19576 16396 19582 16408
rect 22554 16396 22560 16408
rect 22612 16396 22618 16448
rect 38194 16436 38200 16448
rect 38155 16408 38200 16436
rect 38194 16396 38200 16408
rect 38252 16396 38258 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 1118 16192 1124 16244
rect 1176 16232 1182 16244
rect 1176 16204 4108 16232
rect 1176 16192 1182 16204
rect 4080 16164 4108 16204
rect 4448 16204 4752 16232
rect 4448 16164 4476 16204
rect 4080 16136 4476 16164
rect 4525 16167 4583 16173
rect 4525 16133 4537 16167
rect 4571 16164 4583 16167
rect 4614 16164 4620 16176
rect 4571 16136 4620 16164
rect 4571 16133 4583 16136
rect 4525 16127 4583 16133
rect 4614 16124 4620 16136
rect 4672 16124 4678 16176
rect 4724 16164 4752 16204
rect 5534 16192 5540 16244
rect 5592 16232 5598 16244
rect 5997 16235 6055 16241
rect 5997 16232 6009 16235
rect 5592 16204 6009 16232
rect 5592 16192 5598 16204
rect 5997 16201 6009 16204
rect 6043 16201 6055 16235
rect 5997 16195 6055 16201
rect 6086 16192 6092 16244
rect 6144 16232 6150 16244
rect 6362 16232 6368 16244
rect 6144 16204 6368 16232
rect 6144 16192 6150 16204
rect 6362 16192 6368 16204
rect 6420 16192 6426 16244
rect 6641 16235 6699 16241
rect 6641 16201 6653 16235
rect 6687 16232 6699 16235
rect 8386 16232 8392 16244
rect 6687 16204 8392 16232
rect 6687 16201 6699 16204
rect 6641 16195 6699 16201
rect 8386 16192 8392 16204
rect 8444 16192 8450 16244
rect 10413 16235 10471 16241
rect 10413 16201 10425 16235
rect 10459 16232 10471 16235
rect 11606 16232 11612 16244
rect 10459 16204 11612 16232
rect 10459 16201 10471 16204
rect 10413 16195 10471 16201
rect 11606 16192 11612 16204
rect 11664 16192 11670 16244
rect 13354 16192 13360 16244
rect 13412 16232 13418 16244
rect 16209 16235 16267 16241
rect 13412 16204 15148 16232
rect 13412 16192 13418 16204
rect 4724 16136 5014 16164
rect 8694 16136 12434 16164
rect 4246 16096 4252 16108
rect 3450 16068 4108 16096
rect 4207 16068 4252 16096
rect 1578 15988 1584 16040
rect 1636 16028 1642 16040
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1636 16000 2053 16028
rect 1636 15988 1642 16000
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 2866 15988 2872 16040
rect 2924 16028 2930 16040
rect 4080 16028 4108 16068
rect 4246 16056 4252 16068
rect 4304 16056 4310 16108
rect 6549 16099 6607 16105
rect 6549 16065 6561 16099
rect 6595 16065 6607 16099
rect 6549 16059 6607 16065
rect 4982 16028 4988 16040
rect 2924 16000 3924 16028
rect 4080 16000 4988 16028
rect 2924 15988 2930 16000
rect 2304 15895 2362 15901
rect 2304 15861 2316 15895
rect 2350 15892 2362 15895
rect 3326 15892 3332 15904
rect 2350 15864 3332 15892
rect 2350 15861 2362 15864
rect 2304 15855 2362 15861
rect 3326 15852 3332 15864
rect 3384 15852 3390 15904
rect 3602 15852 3608 15904
rect 3660 15892 3666 15904
rect 3789 15895 3847 15901
rect 3789 15892 3801 15895
rect 3660 15864 3801 15892
rect 3660 15852 3666 15864
rect 3789 15861 3801 15864
rect 3835 15861 3847 15895
rect 3896 15892 3924 16000
rect 4982 15988 4988 16000
rect 5040 15988 5046 16040
rect 5166 15988 5172 16040
rect 5224 16028 5230 16040
rect 5994 16028 6000 16040
rect 5224 16000 6000 16028
rect 5224 15988 5230 16000
rect 5994 15988 6000 16000
rect 6052 15988 6058 16040
rect 6564 16028 6592 16059
rect 6638 16056 6644 16108
rect 6696 16096 6702 16108
rect 7193 16099 7251 16105
rect 7193 16096 7205 16099
rect 6696 16068 7205 16096
rect 6696 16056 6702 16068
rect 7193 16065 7205 16068
rect 7239 16065 7251 16099
rect 7193 16059 7251 16065
rect 8754 16056 8760 16108
rect 8812 16096 8818 16108
rect 9677 16099 9735 16105
rect 9677 16096 9689 16099
rect 8812 16068 9689 16096
rect 8812 16056 8818 16068
rect 9677 16065 9689 16068
rect 9723 16065 9735 16099
rect 9677 16059 9735 16065
rect 10134 16056 10140 16108
rect 10192 16096 10198 16108
rect 10321 16099 10379 16105
rect 10321 16096 10333 16099
rect 10192 16068 10333 16096
rect 10192 16056 10198 16068
rect 10321 16065 10333 16068
rect 10367 16065 10379 16099
rect 10962 16096 10968 16108
rect 10923 16068 10968 16096
rect 10321 16059 10379 16065
rect 10962 16056 10968 16068
rect 11020 16056 11026 16108
rect 11054 16056 11060 16108
rect 11112 16096 11118 16108
rect 12161 16099 12219 16105
rect 12161 16096 12173 16099
rect 11112 16068 12173 16096
rect 11112 16056 11118 16068
rect 12161 16065 12173 16068
rect 12207 16065 12219 16099
rect 12406 16096 12434 16136
rect 13814 16124 13820 16176
rect 13872 16164 13878 16176
rect 13872 16136 13917 16164
rect 13872 16124 13878 16136
rect 14458 16124 14464 16176
rect 14516 16124 14522 16176
rect 15120 16164 15148 16204
rect 16209 16201 16221 16235
rect 16255 16232 16267 16235
rect 16390 16232 16396 16244
rect 16255 16204 16396 16232
rect 16255 16201 16267 16204
rect 16209 16195 16267 16201
rect 16390 16192 16396 16204
rect 16448 16192 16454 16244
rect 20070 16232 20076 16244
rect 17880 16204 20076 16232
rect 17880 16173 17908 16204
rect 20070 16192 20076 16204
rect 20128 16192 20134 16244
rect 20809 16235 20867 16241
rect 20809 16201 20821 16235
rect 20855 16232 20867 16235
rect 21082 16232 21088 16244
rect 20855 16204 21088 16232
rect 20855 16201 20867 16204
rect 20809 16195 20867 16201
rect 21082 16192 21088 16204
rect 21140 16192 21146 16244
rect 21192 16204 25912 16232
rect 17129 16167 17187 16173
rect 17129 16164 17141 16167
rect 15120 16136 17141 16164
rect 17129 16133 17141 16136
rect 17175 16133 17187 16167
rect 17129 16127 17187 16133
rect 17865 16167 17923 16173
rect 17865 16133 17877 16167
rect 17911 16133 17923 16167
rect 17865 16127 17923 16133
rect 17957 16167 18015 16173
rect 17957 16133 17969 16167
rect 18003 16164 18015 16167
rect 19429 16167 19487 16173
rect 19429 16164 19441 16167
rect 18003 16136 19441 16164
rect 18003 16133 18015 16136
rect 17957 16127 18015 16133
rect 19429 16133 19441 16136
rect 19475 16133 19487 16167
rect 19429 16127 19487 16133
rect 12802 16096 12808 16108
rect 12406 16068 12808 16096
rect 12161 16059 12219 16065
rect 12802 16056 12808 16068
rect 12860 16056 12866 16108
rect 16117 16099 16175 16105
rect 16117 16065 16129 16099
rect 16163 16065 16175 16099
rect 16117 16059 16175 16065
rect 16853 16099 16911 16105
rect 16853 16065 16865 16099
rect 16899 16096 16911 16099
rect 17310 16096 17316 16108
rect 16899 16068 17316 16096
rect 16899 16065 16911 16068
rect 16853 16059 16911 16065
rect 7098 16028 7104 16040
rect 6564 16000 7104 16028
rect 7098 15988 7104 16000
rect 7156 15988 7162 16040
rect 7469 16031 7527 16037
rect 7469 15997 7481 16031
rect 7515 16028 7527 16031
rect 8662 16028 8668 16040
rect 7515 16000 8668 16028
rect 7515 15997 7527 16000
rect 7469 15991 7527 15997
rect 8662 15988 8668 16000
rect 8720 15988 8726 16040
rect 8846 15988 8852 16040
rect 8904 16028 8910 16040
rect 9217 16031 9275 16037
rect 9217 16028 9229 16031
rect 8904 16000 9229 16028
rect 8904 15988 8910 16000
rect 9217 15997 9229 16000
rect 9263 16028 9275 16031
rect 9950 16028 9956 16040
rect 9263 16000 9956 16028
rect 9263 15997 9275 16000
rect 9217 15991 9275 15997
rect 9950 15988 9956 16000
rect 10008 15988 10014 16040
rect 10594 15988 10600 16040
rect 10652 16028 10658 16040
rect 12897 16031 12955 16037
rect 12897 16028 12909 16031
rect 10652 16000 12909 16028
rect 10652 15988 10658 16000
rect 12897 15997 12909 16000
rect 12943 16028 12955 16031
rect 13541 16031 13599 16037
rect 13541 16028 13553 16031
rect 12943 16000 13553 16028
rect 12943 15997 12955 16000
rect 12897 15991 12955 15997
rect 13541 15997 13553 16000
rect 13587 16028 13599 16031
rect 14274 16028 14280 16040
rect 13587 16000 14280 16028
rect 13587 15997 13599 16000
rect 13541 15991 13599 15997
rect 14274 15988 14280 16000
rect 14332 15988 14338 16040
rect 16132 16028 16160 16059
rect 17310 16056 17316 16068
rect 17368 16056 17374 16108
rect 18966 16056 18972 16108
rect 19024 16096 19030 16108
rect 19337 16099 19395 16105
rect 19337 16096 19349 16099
rect 19024 16068 19349 16096
rect 19024 16056 19030 16068
rect 19337 16065 19349 16068
rect 19383 16065 19395 16099
rect 19978 16096 19984 16108
rect 19939 16068 19984 16096
rect 19337 16059 19395 16065
rect 19978 16056 19984 16068
rect 20036 16056 20042 16108
rect 20717 16099 20775 16105
rect 20717 16065 20729 16099
rect 20763 16096 20775 16099
rect 20806 16096 20812 16108
rect 20763 16068 20812 16096
rect 20763 16065 20775 16068
rect 20717 16059 20775 16065
rect 20806 16056 20812 16068
rect 20864 16056 20870 16108
rect 18506 16028 18512 16040
rect 16132 16000 17632 16028
rect 18467 16000 18512 16028
rect 13262 15960 13268 15972
rect 5552 15932 6776 15960
rect 5552 15892 5580 15932
rect 3896 15864 5580 15892
rect 6748 15892 6776 15932
rect 8496 15932 13268 15960
rect 8496 15892 8524 15932
rect 13262 15920 13268 15932
rect 13320 15920 13326 15972
rect 15102 15920 15108 15972
rect 15160 15960 15166 15972
rect 16574 15960 16580 15972
rect 15160 15932 16580 15960
rect 15160 15920 15166 15932
rect 16574 15920 16580 15932
rect 16632 15920 16638 15972
rect 6748 15864 8524 15892
rect 9769 15895 9827 15901
rect 3789 15855 3847 15861
rect 9769 15861 9781 15895
rect 9815 15892 9827 15895
rect 10962 15892 10968 15904
rect 9815 15864 10968 15892
rect 9815 15861 9827 15864
rect 9769 15855 9827 15861
rect 10962 15852 10968 15864
rect 11020 15852 11026 15904
rect 11057 15895 11115 15901
rect 11057 15861 11069 15895
rect 11103 15892 11115 15895
rect 15010 15892 15016 15904
rect 11103 15864 15016 15892
rect 11103 15861 11115 15864
rect 11057 15855 11115 15861
rect 15010 15852 15016 15864
rect 15068 15852 15074 15904
rect 15286 15892 15292 15904
rect 15247 15864 15292 15892
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 17604 15892 17632 16000
rect 18506 15988 18512 16000
rect 18564 15988 18570 16040
rect 18690 15988 18696 16040
rect 18748 16028 18754 16040
rect 21192 16028 21220 16204
rect 21634 16124 21640 16176
rect 21692 16164 21698 16176
rect 22189 16167 22247 16173
rect 22189 16164 22201 16167
rect 21692 16136 22201 16164
rect 21692 16124 21698 16136
rect 22189 16133 22201 16136
rect 22235 16133 22247 16167
rect 22189 16127 22247 16133
rect 22462 16124 22468 16176
rect 22520 16164 22526 16176
rect 23106 16164 23112 16176
rect 22520 16136 23112 16164
rect 22520 16124 22526 16136
rect 23106 16124 23112 16136
rect 23164 16124 23170 16176
rect 25884 16096 25912 16204
rect 26142 16192 26148 16244
rect 26200 16232 26206 16244
rect 27249 16235 27307 16241
rect 27249 16232 27261 16235
rect 26200 16204 27261 16232
rect 26200 16192 26206 16204
rect 27249 16201 27261 16204
rect 27295 16201 27307 16235
rect 27249 16195 27307 16201
rect 28442 16164 28448 16176
rect 27172 16136 28448 16164
rect 27172 16105 27200 16136
rect 28442 16124 28448 16136
rect 28500 16124 28506 16176
rect 28534 16124 28540 16176
rect 28592 16164 28598 16176
rect 28592 16136 35894 16164
rect 28592 16124 28598 16136
rect 27157 16099 27215 16105
rect 27157 16096 27169 16099
rect 25884 16068 27169 16096
rect 27157 16065 27169 16068
rect 27203 16065 27215 16099
rect 27157 16059 27215 16065
rect 27614 16056 27620 16108
rect 27672 16096 27678 16108
rect 27893 16099 27951 16105
rect 27893 16096 27905 16099
rect 27672 16068 27905 16096
rect 27672 16056 27678 16068
rect 27893 16065 27905 16068
rect 27939 16065 27951 16099
rect 28718 16096 28724 16108
rect 28679 16068 28724 16096
rect 27893 16059 27951 16065
rect 28718 16056 28724 16068
rect 28776 16056 28782 16108
rect 35866 16096 35894 16136
rect 37274 16096 37280 16108
rect 35866 16068 37280 16096
rect 37274 16056 37280 16068
rect 37332 16056 37338 16108
rect 38286 16096 38292 16108
rect 38247 16068 38292 16096
rect 38286 16056 38292 16068
rect 38344 16056 38350 16108
rect 18748 16000 21220 16028
rect 22097 16031 22155 16037
rect 18748 15988 18754 16000
rect 22097 15997 22109 16031
rect 22143 16028 22155 16031
rect 27985 16031 28043 16037
rect 22143 16000 23060 16028
rect 22143 15997 22155 16000
rect 22097 15991 22155 15997
rect 20073 15963 20131 15969
rect 20073 15929 20085 15963
rect 20119 15960 20131 15963
rect 22278 15960 22284 15972
rect 20119 15932 22284 15960
rect 20119 15929 20131 15932
rect 20073 15923 20131 15929
rect 22278 15920 22284 15932
rect 22336 15920 22342 15972
rect 23032 15960 23060 16000
rect 27985 15997 27997 16031
rect 28031 16028 28043 16031
rect 30374 16028 30380 16040
rect 28031 16000 30380 16028
rect 28031 15997 28043 16000
rect 27985 15991 28043 15997
rect 30374 15988 30380 16000
rect 30432 15988 30438 16040
rect 38010 16028 38016 16040
rect 35866 16000 38016 16028
rect 26234 15960 26240 15972
rect 23032 15932 26240 15960
rect 26234 15920 26240 15932
rect 26292 15920 26298 15972
rect 28537 15963 28595 15969
rect 28537 15929 28549 15963
rect 28583 15960 28595 15963
rect 35866 15960 35894 16000
rect 38010 15988 38016 16000
rect 38068 15988 38074 16040
rect 28583 15932 35894 15960
rect 28583 15929 28595 15932
rect 28537 15923 28595 15929
rect 20162 15892 20168 15904
rect 17604 15864 20168 15892
rect 20162 15852 20168 15864
rect 20220 15852 20226 15904
rect 29730 15852 29736 15904
rect 29788 15892 29794 15904
rect 38105 15895 38163 15901
rect 38105 15892 38117 15895
rect 29788 15864 38117 15892
rect 29788 15852 29794 15864
rect 38105 15861 38117 15864
rect 38151 15861 38163 15895
rect 38105 15855 38163 15861
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 3602 15648 3608 15700
rect 3660 15688 3666 15700
rect 9122 15688 9128 15700
rect 3660 15660 6855 15688
rect 9083 15660 9128 15688
rect 3660 15648 3666 15660
rect 3252 15592 3464 15620
rect 1857 15555 1915 15561
rect 1857 15521 1869 15555
rect 1903 15552 1915 15555
rect 3252 15552 3280 15592
rect 1903 15524 3280 15552
rect 3329 15555 3387 15561
rect 1903 15521 1915 15524
rect 1857 15515 1915 15521
rect 3329 15521 3341 15555
rect 3375 15521 3387 15555
rect 3436 15552 3464 15592
rect 3510 15580 3516 15632
rect 3568 15620 3574 15632
rect 3568 15592 4292 15620
rect 3568 15580 3574 15592
rect 3786 15552 3792 15564
rect 3436 15524 3792 15552
rect 3329 15515 3387 15521
rect 1578 15484 1584 15496
rect 1539 15456 1584 15484
rect 1578 15444 1584 15456
rect 1636 15444 1642 15496
rect 3344 15484 3372 15515
rect 3786 15512 3792 15524
rect 3844 15512 3850 15564
rect 4062 15512 4068 15564
rect 4120 15552 4126 15564
rect 4157 15555 4215 15561
rect 4157 15552 4169 15555
rect 4120 15524 4169 15552
rect 4120 15512 4126 15524
rect 4157 15521 4169 15524
rect 4203 15521 4215 15555
rect 4264 15552 4292 15592
rect 5626 15580 5632 15632
rect 5684 15620 5690 15632
rect 6730 15620 6736 15632
rect 5684 15592 6736 15620
rect 5684 15580 5690 15592
rect 6730 15580 6736 15592
rect 6788 15580 6794 15632
rect 4433 15555 4491 15561
rect 4433 15552 4445 15555
rect 4264 15524 4445 15552
rect 4157 15515 4215 15521
rect 4433 15521 4445 15524
rect 4479 15521 4491 15555
rect 4433 15515 4491 15521
rect 4798 15512 4804 15564
rect 4856 15552 4862 15564
rect 5905 15555 5963 15561
rect 4856 15524 5580 15552
rect 4856 15512 4862 15524
rect 3970 15484 3976 15496
rect 3344 15456 3976 15484
rect 3970 15444 3976 15456
rect 4028 15444 4034 15496
rect 5552 15470 5580 15524
rect 5905 15521 5917 15555
rect 5951 15552 5963 15555
rect 6270 15552 6276 15564
rect 5951 15524 6276 15552
rect 5951 15521 5963 15524
rect 5905 15515 5963 15521
rect 6270 15512 6276 15524
rect 6328 15512 6334 15564
rect 6827 15552 6855 15660
rect 9122 15648 9128 15660
rect 9180 15648 9186 15700
rect 12526 15688 12532 15700
rect 12360 15660 12532 15688
rect 8846 15580 8852 15632
rect 8904 15620 8910 15632
rect 10410 15620 10416 15632
rect 8904 15592 10416 15620
rect 8904 15580 8910 15592
rect 10410 15580 10416 15592
rect 10468 15580 10474 15632
rect 12360 15620 12388 15660
rect 12526 15648 12532 15660
rect 12584 15648 12590 15700
rect 12986 15688 12992 15700
rect 12947 15660 12992 15688
rect 12986 15648 12992 15660
rect 13044 15648 13050 15700
rect 19150 15688 19156 15700
rect 15396 15660 19156 15688
rect 11992 15592 12388 15620
rect 7009 15555 7067 15561
rect 7009 15552 7021 15555
rect 6827 15524 7021 15552
rect 7009 15521 7021 15524
rect 7055 15521 7067 15555
rect 7009 15515 7067 15521
rect 7098 15512 7104 15564
rect 7156 15552 7162 15564
rect 10134 15552 10140 15564
rect 7156 15524 10140 15552
rect 7156 15512 7162 15524
rect 10134 15512 10140 15524
rect 10192 15512 10198 15564
rect 10873 15555 10931 15561
rect 10873 15521 10885 15555
rect 10919 15552 10931 15555
rect 11992 15552 12020 15592
rect 12434 15580 12440 15632
rect 12492 15620 12498 15632
rect 15396 15620 15424 15660
rect 19150 15648 19156 15660
rect 19208 15688 19214 15700
rect 20438 15688 20444 15700
rect 19208 15660 20444 15688
rect 19208 15648 19214 15660
rect 20438 15648 20444 15660
rect 20496 15648 20502 15700
rect 21085 15691 21143 15697
rect 21085 15657 21097 15691
rect 21131 15688 21143 15691
rect 21634 15688 21640 15700
rect 21131 15660 21640 15688
rect 21131 15657 21143 15660
rect 21085 15651 21143 15657
rect 21634 15648 21640 15660
rect 21692 15648 21698 15700
rect 12492 15592 14504 15620
rect 12492 15580 12498 15592
rect 10919 15524 12020 15552
rect 10919 15521 10931 15524
rect 10873 15515 10931 15521
rect 12066 15512 12072 15564
rect 12124 15512 12130 15564
rect 12342 15552 12348 15564
rect 12303 15524 12348 15552
rect 12342 15512 12348 15524
rect 12400 15512 12406 15564
rect 12802 15512 12808 15564
rect 12860 15552 12866 15564
rect 12860 15524 14412 15552
rect 12860 15512 12866 15524
rect 6730 15484 6736 15496
rect 6691 15456 6736 15484
rect 6730 15444 6736 15456
rect 6788 15444 6794 15496
rect 9306 15484 9312 15496
rect 9267 15456 9312 15484
rect 9306 15444 9312 15456
rect 9364 15444 9370 15496
rect 9769 15487 9827 15493
rect 9769 15453 9781 15487
rect 9815 15484 9827 15487
rect 9858 15484 9864 15496
rect 9815 15456 9864 15484
rect 9815 15453 9827 15456
rect 9769 15447 9827 15453
rect 9858 15444 9864 15456
rect 9916 15444 9922 15496
rect 10594 15484 10600 15496
rect 10555 15456 10600 15484
rect 10594 15444 10600 15456
rect 10652 15444 10658 15496
rect 12084 15484 12112 15512
rect 12897 15487 12955 15493
rect 12897 15484 12909 15487
rect 12084 15456 12909 15484
rect 12897 15453 12909 15456
rect 12943 15453 12955 15487
rect 12897 15447 12955 15453
rect 13262 15444 13268 15496
rect 13320 15484 13326 15496
rect 13541 15487 13599 15493
rect 13541 15484 13553 15487
rect 13320 15456 13553 15484
rect 13320 15444 13326 15456
rect 13541 15453 13553 15456
rect 13587 15453 13599 15487
rect 13541 15447 13599 15453
rect 2130 15376 2136 15428
rect 2188 15416 2194 15428
rect 2188 15388 2346 15416
rect 2188 15376 2194 15388
rect 7466 15376 7472 15428
rect 7524 15376 7530 15428
rect 12618 15416 12624 15428
rect 12098 15388 12624 15416
rect 12618 15376 12624 15388
rect 12676 15376 12682 15428
rect 13633 15419 13691 15425
rect 13633 15416 13645 15419
rect 12912 15388 13645 15416
rect 7190 15308 7196 15360
rect 7248 15348 7254 15360
rect 8481 15351 8539 15357
rect 8481 15348 8493 15351
rect 7248 15320 8493 15348
rect 7248 15308 7254 15320
rect 8481 15317 8493 15320
rect 8527 15317 8539 15351
rect 8481 15311 8539 15317
rect 9861 15351 9919 15357
rect 9861 15317 9873 15351
rect 9907 15348 9919 15351
rect 9950 15348 9956 15360
rect 9907 15320 9956 15348
rect 9907 15317 9919 15320
rect 9861 15311 9919 15317
rect 9950 15308 9956 15320
rect 10008 15308 10014 15360
rect 10870 15308 10876 15360
rect 10928 15348 10934 15360
rect 12912 15348 12940 15388
rect 13633 15385 13645 15388
rect 13679 15385 13691 15419
rect 14384 15416 14412 15524
rect 14476 15493 14504 15592
rect 15212 15592 15424 15620
rect 15212 15561 15240 15592
rect 15470 15580 15476 15632
rect 15528 15620 15534 15632
rect 15528 15592 16160 15620
rect 15528 15580 15534 15592
rect 16132 15561 16160 15592
rect 16298 15580 16304 15632
rect 16356 15620 16362 15632
rect 19242 15620 19248 15632
rect 16356 15592 19248 15620
rect 16356 15580 16362 15592
rect 19242 15580 19248 15592
rect 19300 15580 19306 15632
rect 20070 15580 20076 15632
rect 20128 15620 20134 15632
rect 29825 15623 29883 15629
rect 29825 15620 29837 15623
rect 20128 15592 29837 15620
rect 20128 15580 20134 15592
rect 29825 15589 29837 15592
rect 29871 15589 29883 15623
rect 29825 15583 29883 15589
rect 15197 15555 15255 15561
rect 15197 15521 15209 15555
rect 15243 15521 15255 15555
rect 15197 15515 15255 15521
rect 16117 15555 16175 15561
rect 16117 15521 16129 15555
rect 16163 15552 16175 15555
rect 16390 15552 16396 15564
rect 16163 15524 16396 15552
rect 16163 15521 16175 15524
rect 16117 15515 16175 15521
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 16574 15512 16580 15564
rect 16632 15552 16638 15564
rect 18966 15552 18972 15564
rect 16632 15524 18972 15552
rect 16632 15512 16638 15524
rect 18966 15512 18972 15524
rect 19024 15512 19030 15564
rect 19058 15512 19064 15564
rect 19116 15552 19122 15564
rect 20165 15555 20223 15561
rect 20165 15552 20177 15555
rect 19116 15524 20177 15552
rect 19116 15512 19122 15524
rect 20165 15521 20177 15524
rect 20211 15521 20223 15555
rect 20165 15515 20223 15521
rect 20622 15512 20628 15564
rect 20680 15552 20686 15564
rect 21729 15555 21787 15561
rect 21729 15552 21741 15555
rect 20680 15524 21741 15552
rect 20680 15512 20686 15524
rect 21729 15521 21741 15524
rect 21775 15521 21787 15555
rect 21729 15515 21787 15521
rect 22741 15555 22799 15561
rect 22741 15521 22753 15555
rect 22787 15552 22799 15555
rect 24854 15552 24860 15564
rect 22787 15524 24860 15552
rect 22787 15521 22799 15524
rect 22741 15515 22799 15521
rect 24854 15512 24860 15524
rect 24912 15552 24918 15564
rect 28534 15552 28540 15564
rect 24912 15524 28540 15552
rect 24912 15512 24918 15524
rect 28534 15512 28540 15524
rect 28592 15512 28598 15564
rect 14461 15487 14519 15493
rect 14461 15453 14473 15487
rect 14507 15484 14519 15487
rect 14550 15484 14556 15496
rect 14507 15456 14556 15484
rect 14507 15453 14519 15456
rect 14461 15447 14519 15453
rect 14550 15444 14556 15456
rect 14608 15444 14614 15496
rect 16761 15487 16819 15493
rect 16761 15453 16773 15487
rect 16807 15484 16819 15487
rect 17310 15484 17316 15496
rect 16807 15456 17316 15484
rect 16807 15453 16819 15456
rect 16761 15447 16819 15453
rect 17310 15444 17316 15456
rect 17368 15484 17374 15496
rect 18046 15484 18052 15496
rect 17368 15456 18052 15484
rect 17368 15444 17374 15456
rect 18046 15444 18052 15456
rect 18104 15444 18110 15496
rect 19429 15487 19487 15493
rect 19429 15453 19441 15487
rect 19475 15453 19487 15487
rect 19429 15447 19487 15453
rect 14384 15388 15240 15416
rect 13633 15379 13691 15385
rect 10928 15320 12940 15348
rect 10928 15308 10934 15320
rect 12986 15308 12992 15360
rect 13044 15348 13050 15360
rect 14458 15348 14464 15360
rect 13044 15320 14464 15348
rect 13044 15308 13050 15320
rect 14458 15308 14464 15320
rect 14516 15308 14522 15360
rect 14553 15351 14611 15357
rect 14553 15317 14565 15351
rect 14599 15348 14611 15351
rect 14734 15348 14740 15360
rect 14599 15320 14740 15348
rect 14599 15317 14611 15320
rect 14553 15311 14611 15317
rect 14734 15308 14740 15320
rect 14792 15308 14798 15360
rect 15212 15348 15240 15388
rect 15286 15376 15292 15428
rect 15344 15416 15350 15428
rect 15344 15388 15389 15416
rect 15344 15376 15350 15388
rect 16666 15376 16672 15428
rect 16724 15416 16730 15428
rect 16942 15416 16948 15428
rect 16724 15388 16948 15416
rect 16724 15376 16730 15388
rect 16942 15376 16948 15388
rect 17000 15416 17006 15428
rect 17037 15419 17095 15425
rect 17037 15416 17049 15419
rect 17000 15388 17049 15416
rect 17000 15376 17006 15388
rect 17037 15385 17049 15388
rect 17083 15385 17095 15419
rect 18230 15416 18236 15428
rect 18191 15388 18236 15416
rect 17037 15379 17095 15385
rect 18230 15376 18236 15388
rect 18288 15376 18294 15428
rect 18325 15419 18383 15425
rect 18325 15385 18337 15419
rect 18371 15385 18383 15419
rect 18325 15379 18383 15385
rect 18877 15419 18935 15425
rect 18877 15385 18889 15419
rect 18923 15416 18935 15419
rect 18966 15416 18972 15428
rect 18923 15388 18972 15416
rect 18923 15385 18935 15388
rect 18877 15379 18935 15385
rect 18138 15348 18144 15360
rect 15212 15320 18144 15348
rect 18138 15308 18144 15320
rect 18196 15308 18202 15360
rect 18340 15348 18368 15379
rect 18966 15376 18972 15388
rect 19024 15376 19030 15428
rect 19444 15416 19472 15447
rect 19886 15444 19892 15496
rect 19944 15484 19950 15496
rect 20073 15487 20131 15493
rect 20073 15484 20085 15487
rect 19944 15456 20085 15484
rect 19944 15444 19950 15456
rect 20073 15453 20085 15456
rect 20119 15453 20131 15487
rect 20073 15447 20131 15453
rect 20254 15444 20260 15496
rect 20312 15484 20318 15496
rect 20993 15487 21051 15493
rect 20312 15456 20852 15484
rect 20312 15444 20318 15456
rect 20824 15416 20852 15456
rect 20993 15453 21005 15487
rect 21039 15484 21051 15487
rect 21174 15484 21180 15496
rect 21039 15456 21180 15484
rect 21039 15453 21051 15456
rect 20993 15447 21051 15453
rect 21174 15444 21180 15456
rect 21232 15444 21238 15496
rect 27062 15444 27068 15496
rect 27120 15484 27126 15496
rect 27801 15487 27859 15493
rect 27801 15484 27813 15487
rect 27120 15456 27813 15484
rect 27120 15444 27126 15456
rect 27801 15453 27813 15456
rect 27847 15453 27859 15487
rect 29730 15484 29736 15496
rect 29691 15456 29736 15484
rect 27801 15447 27859 15453
rect 29730 15444 29736 15456
rect 29788 15444 29794 15496
rect 21821 15419 21879 15425
rect 21821 15416 21833 15419
rect 19444 15388 20760 15416
rect 20824 15388 21833 15416
rect 19521 15351 19579 15357
rect 19521 15348 19533 15351
rect 18340 15320 19533 15348
rect 19521 15317 19533 15320
rect 19567 15317 19579 15351
rect 20732 15348 20760 15388
rect 21821 15385 21833 15388
rect 21867 15385 21879 15419
rect 21821 15379 21879 15385
rect 23382 15348 23388 15360
rect 20732 15320 23388 15348
rect 19521 15311 19579 15317
rect 23382 15308 23388 15320
rect 23440 15308 23446 15360
rect 27617 15351 27675 15357
rect 27617 15317 27629 15351
rect 27663 15348 27675 15351
rect 27982 15348 27988 15360
rect 27663 15320 27988 15348
rect 27663 15317 27675 15320
rect 27617 15311 27675 15317
rect 27982 15308 27988 15320
rect 28040 15308 28046 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 2682 15104 2688 15156
rect 2740 15144 2746 15156
rect 3326 15144 3332 15156
rect 2740 15116 3004 15144
rect 3287 15116 3332 15144
rect 2740 15104 2746 15116
rect 2976 14994 3004 15116
rect 3326 15104 3332 15116
rect 3384 15104 3390 15156
rect 5534 15144 5540 15156
rect 5495 15116 5540 15144
rect 5534 15104 5540 15116
rect 5592 15144 5598 15156
rect 6086 15144 6092 15156
rect 5592 15116 6092 15144
rect 5592 15104 5598 15116
rect 6086 15104 6092 15116
rect 6144 15104 6150 15156
rect 8573 15147 8631 15153
rect 8573 15113 8585 15147
rect 8619 15144 8631 15147
rect 9030 15144 9036 15156
rect 8619 15116 9036 15144
rect 8619 15113 8631 15116
rect 8573 15107 8631 15113
rect 9030 15104 9036 15116
rect 9088 15104 9094 15156
rect 9490 15104 9496 15156
rect 9548 15144 9554 15156
rect 9548 15116 13952 15144
rect 9548 15104 9554 15116
rect 4062 15076 4068 15088
rect 4023 15048 4068 15076
rect 4062 15036 4068 15048
rect 4120 15036 4126 15088
rect 9398 15036 9404 15088
rect 9456 15076 9462 15088
rect 9456 15048 9798 15076
rect 9456 15036 9462 15048
rect 11882 15036 11888 15088
rect 11940 15076 11946 15088
rect 12526 15076 12532 15088
rect 11940 15048 12532 15076
rect 11940 15036 11946 15048
rect 12526 15036 12532 15048
rect 12584 15036 12590 15088
rect 13924 15076 13952 15116
rect 15286 15104 15292 15156
rect 15344 15144 15350 15156
rect 15565 15147 15623 15153
rect 15565 15144 15577 15147
rect 15344 15116 15577 15144
rect 15344 15104 15350 15116
rect 15565 15113 15577 15116
rect 15611 15113 15623 15147
rect 15565 15107 15623 15113
rect 18874 15104 18880 15156
rect 18932 15144 18938 15156
rect 19150 15144 19156 15156
rect 18932 15116 19156 15144
rect 18932 15104 18938 15116
rect 19150 15104 19156 15116
rect 19208 15104 19214 15156
rect 19334 15144 19340 15156
rect 19295 15116 19340 15144
rect 19334 15104 19340 15116
rect 19392 15104 19398 15156
rect 16209 15079 16267 15085
rect 13924 15048 15516 15076
rect 6178 15008 6184 15020
rect 5198 14980 6184 15008
rect 6178 14968 6184 14980
rect 6236 14968 6242 15020
rect 8202 14968 8208 15020
rect 8260 14968 8266 15020
rect 12066 14968 12072 15020
rect 12124 15008 12130 15020
rect 12161 15011 12219 15017
rect 12161 15008 12173 15011
rect 12124 14980 12173 15008
rect 12124 14968 12130 14980
rect 12161 14977 12173 14980
rect 12207 14977 12219 15011
rect 12161 14971 12219 14977
rect 13538 14968 13544 15020
rect 13596 14968 13602 15020
rect 13722 14968 13728 15020
rect 13780 15008 13786 15020
rect 15488 15017 15516 15048
rect 16209 15045 16221 15079
rect 16255 15076 16267 15079
rect 17037 15079 17095 15085
rect 17037 15076 17049 15079
rect 16255 15048 17049 15076
rect 16255 15045 16267 15048
rect 16209 15039 16267 15045
rect 17037 15045 17049 15048
rect 17083 15045 17095 15079
rect 17037 15039 17095 15045
rect 17788 15048 21312 15076
rect 14829 15011 14887 15017
rect 14829 15008 14841 15011
rect 13780 14980 14841 15008
rect 13780 14968 13786 14980
rect 14829 14977 14841 14980
rect 14875 14977 14887 15011
rect 14829 14971 14887 14977
rect 15473 15011 15531 15017
rect 15473 14977 15485 15011
rect 15519 14977 15531 15011
rect 15473 14971 15531 14977
rect 15838 14968 15844 15020
rect 15896 15008 15902 15020
rect 16117 15011 16175 15017
rect 16117 15008 16129 15011
rect 15896 14980 16129 15008
rect 15896 14968 15902 14980
rect 16117 14977 16129 14980
rect 16163 14977 16175 15011
rect 16117 14971 16175 14977
rect 1578 14940 1584 14952
rect 1539 14912 1584 14940
rect 1578 14900 1584 14912
rect 1636 14900 1642 14952
rect 1854 14940 1860 14952
rect 1688 14912 1860 14940
rect 1210 14832 1216 14884
rect 1268 14872 1274 14884
rect 1688 14872 1716 14912
rect 1854 14900 1860 14912
rect 1912 14900 1918 14952
rect 3786 14940 3792 14952
rect 3747 14912 3792 14940
rect 3786 14900 3792 14912
rect 3844 14900 3850 14952
rect 6822 14940 6828 14952
rect 6783 14912 6828 14940
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 7101 14943 7159 14949
rect 7101 14909 7113 14943
rect 7147 14940 7159 14943
rect 7650 14940 7656 14952
rect 7147 14912 7656 14940
rect 7147 14909 7159 14912
rect 7101 14903 7159 14909
rect 7650 14900 7656 14912
rect 7708 14900 7714 14952
rect 9030 14940 9036 14952
rect 8991 14912 9036 14940
rect 9030 14900 9036 14912
rect 9088 14900 9094 14952
rect 9398 14900 9404 14952
rect 9456 14940 9462 14952
rect 9456 14912 10364 14940
rect 9456 14900 9462 14912
rect 1268 14844 1716 14872
rect 1268 14832 1274 14844
rect 8478 14832 8484 14884
rect 8536 14872 8542 14884
rect 10336 14872 10364 14912
rect 10502 14900 10508 14952
rect 10560 14940 10566 14952
rect 12437 14943 12495 14949
rect 12437 14940 12449 14943
rect 10560 14912 12449 14940
rect 10560 14900 10566 14912
rect 12437 14909 12449 14912
rect 12483 14940 12495 14943
rect 16945 14943 17003 14949
rect 12483 14912 15240 14940
rect 12483 14909 12495 14912
rect 12437 14903 12495 14909
rect 10781 14875 10839 14881
rect 10781 14872 10793 14875
rect 8536 14844 9168 14872
rect 10336 14844 10793 14872
rect 8536 14832 8542 14844
rect 9140 14804 9168 14844
rect 10781 14841 10793 14844
rect 10827 14841 10839 14875
rect 10781 14835 10839 14841
rect 13909 14875 13967 14881
rect 13909 14841 13921 14875
rect 13955 14872 13967 14875
rect 14182 14872 14188 14884
rect 13955 14844 14188 14872
rect 13955 14841 13967 14844
rect 13909 14835 13967 14841
rect 14182 14832 14188 14844
rect 14240 14832 14246 14884
rect 14366 14832 14372 14884
rect 14424 14872 14430 14884
rect 15102 14872 15108 14884
rect 14424 14844 15108 14872
rect 14424 14832 14430 14844
rect 15102 14832 15108 14844
rect 15160 14832 15166 14884
rect 15212 14872 15240 14912
rect 16945 14909 16957 14943
rect 16991 14940 17003 14943
rect 17586 14940 17592 14952
rect 16991 14912 17592 14940
rect 16991 14909 17003 14912
rect 16945 14903 17003 14909
rect 17586 14900 17592 14912
rect 17644 14900 17650 14952
rect 17788 14872 17816 15048
rect 21284 15020 21312 15048
rect 18046 14968 18052 15020
rect 18104 15008 18110 15020
rect 18417 15011 18475 15017
rect 18417 15008 18429 15011
rect 18104 14980 18429 15008
rect 18104 14968 18110 14980
rect 18417 14977 18429 14980
rect 18463 15008 18475 15011
rect 18874 15008 18880 15020
rect 18463 14980 18880 15008
rect 18463 14977 18475 14980
rect 18417 14971 18475 14977
rect 18874 14968 18880 14980
rect 18932 14968 18938 15020
rect 19334 14968 19340 15020
rect 19392 15008 19398 15020
rect 19521 15011 19579 15017
rect 19521 15008 19533 15011
rect 19392 14980 19533 15008
rect 19392 14968 19398 14980
rect 19521 14977 19533 14980
rect 19567 14977 19579 15011
rect 19521 14971 19579 14977
rect 20165 15011 20223 15017
rect 20165 14977 20177 15011
rect 20211 14977 20223 15011
rect 20165 14971 20223 14977
rect 17862 14900 17868 14952
rect 17920 14940 17926 14952
rect 18598 14940 18604 14952
rect 17920 14912 17965 14940
rect 18559 14912 18604 14940
rect 17920 14900 17926 14912
rect 18598 14900 18604 14912
rect 18656 14900 18662 14952
rect 18690 14900 18696 14952
rect 18748 14940 18754 14952
rect 20180 14940 20208 14971
rect 20438 14968 20444 15020
rect 20496 15008 20502 15020
rect 20625 15011 20683 15017
rect 20625 15008 20637 15011
rect 20496 14980 20637 15008
rect 20496 14968 20502 14980
rect 20625 14977 20637 14980
rect 20671 14977 20683 15011
rect 20625 14971 20683 14977
rect 21266 14968 21272 15020
rect 21324 15008 21330 15020
rect 22189 15011 22247 15017
rect 22189 15008 22201 15011
rect 21324 14980 22201 15008
rect 21324 14968 21330 14980
rect 22189 14977 22201 14980
rect 22235 14977 22247 15011
rect 27982 15008 27988 15020
rect 27943 14980 27988 15008
rect 22189 14971 22247 14977
rect 27982 14968 27988 14980
rect 28040 14968 28046 15020
rect 18748 14912 20208 14940
rect 25685 14943 25743 14949
rect 18748 14900 18754 14912
rect 25685 14909 25697 14943
rect 25731 14940 25743 14943
rect 25958 14940 25964 14952
rect 25731 14912 25964 14940
rect 25731 14909 25743 14912
rect 25685 14903 25743 14909
rect 25958 14900 25964 14912
rect 26016 14900 26022 14952
rect 15212 14844 17816 14872
rect 18414 14832 18420 14884
rect 18472 14872 18478 14884
rect 20717 14875 20775 14881
rect 20717 14872 20729 14875
rect 18472 14844 20729 14872
rect 18472 14832 18478 14844
rect 20717 14841 20729 14844
rect 20763 14841 20775 14875
rect 20717 14835 20775 14841
rect 9290 14807 9348 14813
rect 9290 14804 9302 14807
rect 9140 14776 9302 14804
rect 9290 14773 9302 14776
rect 9336 14773 9348 14807
rect 9290 14767 9348 14773
rect 9398 14764 9404 14816
rect 9456 14804 9462 14816
rect 10686 14804 10692 14816
rect 9456 14776 10692 14804
rect 9456 14764 9462 14776
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 11790 14764 11796 14816
rect 11848 14804 11854 14816
rect 12066 14804 12072 14816
rect 11848 14776 12072 14804
rect 11848 14764 11854 14776
rect 12066 14764 12072 14776
rect 12124 14764 12130 14816
rect 12526 14764 12532 14816
rect 12584 14804 12590 14816
rect 13170 14804 13176 14816
rect 12584 14776 13176 14804
rect 12584 14764 12590 14776
rect 13170 14764 13176 14776
rect 13228 14804 13234 14816
rect 13722 14804 13728 14816
rect 13228 14776 13728 14804
rect 13228 14764 13234 14776
rect 13722 14764 13728 14776
rect 13780 14764 13786 14816
rect 14458 14764 14464 14816
rect 14516 14804 14522 14816
rect 14921 14807 14979 14813
rect 14921 14804 14933 14807
rect 14516 14776 14933 14804
rect 14516 14764 14522 14776
rect 14921 14773 14933 14776
rect 14967 14773 14979 14807
rect 14921 14767 14979 14773
rect 17770 14764 17776 14816
rect 17828 14804 17834 14816
rect 18782 14804 18788 14816
rect 17828 14776 18788 14804
rect 17828 14764 17834 14776
rect 18782 14764 18788 14776
rect 18840 14764 18846 14816
rect 19610 14764 19616 14816
rect 19668 14804 19674 14816
rect 19981 14807 20039 14813
rect 19981 14804 19993 14807
rect 19668 14776 19993 14804
rect 19668 14764 19674 14776
rect 19981 14773 19993 14776
rect 20027 14773 20039 14807
rect 19981 14767 20039 14773
rect 22005 14807 22063 14813
rect 22005 14773 22017 14807
rect 22051 14804 22063 14807
rect 22094 14804 22100 14816
rect 22051 14776 22100 14804
rect 22051 14773 22063 14776
rect 22005 14767 22063 14773
rect 22094 14764 22100 14776
rect 22152 14764 22158 14816
rect 26142 14764 26148 14816
rect 26200 14804 26206 14816
rect 27801 14807 27859 14813
rect 27801 14804 27813 14807
rect 26200 14776 27813 14804
rect 26200 14764 26206 14776
rect 27801 14773 27813 14776
rect 27847 14773 27859 14807
rect 27801 14767 27859 14773
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 3329 14603 3387 14609
rect 3329 14569 3341 14603
rect 3375 14600 3387 14603
rect 3418 14600 3424 14612
rect 3375 14572 3424 14600
rect 3375 14569 3387 14572
rect 3329 14563 3387 14569
rect 3418 14560 3424 14572
rect 3476 14560 3482 14612
rect 4798 14560 4804 14612
rect 4856 14600 4862 14612
rect 5166 14600 5172 14612
rect 4856 14572 5172 14600
rect 4856 14560 4862 14572
rect 5166 14560 5172 14572
rect 5224 14560 5230 14612
rect 5534 14600 5540 14612
rect 5495 14572 5540 14600
rect 5534 14560 5540 14572
rect 5592 14560 5598 14612
rect 6178 14600 6184 14612
rect 6139 14572 6184 14600
rect 6178 14560 6184 14572
rect 6236 14560 6242 14612
rect 9388 14603 9446 14609
rect 9388 14569 9400 14603
rect 9434 14600 9446 14603
rect 12342 14600 12348 14612
rect 9434 14572 12348 14600
rect 9434 14569 9446 14572
rect 9388 14563 9446 14569
rect 12342 14560 12348 14572
rect 12400 14560 12406 14612
rect 13078 14560 13084 14612
rect 13136 14600 13142 14612
rect 14540 14603 14598 14609
rect 14540 14600 14552 14603
rect 13136 14572 14552 14600
rect 13136 14560 13142 14572
rect 14540 14569 14552 14572
rect 14586 14600 14598 14603
rect 14918 14600 14924 14612
rect 14586 14572 14924 14600
rect 14586 14569 14598 14572
rect 14540 14563 14598 14569
rect 14918 14560 14924 14572
rect 14976 14560 14982 14612
rect 16022 14600 16028 14612
rect 15983 14572 16028 14600
rect 16022 14560 16028 14572
rect 16080 14560 16086 14612
rect 17862 14560 17868 14612
rect 17920 14600 17926 14612
rect 21913 14603 21971 14609
rect 21913 14600 21925 14603
rect 17920 14572 21925 14600
rect 17920 14560 17926 14572
rect 21913 14569 21925 14572
rect 21959 14569 21971 14603
rect 21913 14563 21971 14569
rect 25501 14603 25559 14609
rect 25501 14569 25513 14603
rect 25547 14600 25559 14603
rect 26050 14600 26056 14612
rect 25547 14572 26056 14600
rect 25547 14569 25559 14572
rect 25501 14563 25559 14569
rect 26050 14560 26056 14572
rect 26108 14600 26114 14612
rect 26329 14603 26387 14609
rect 26329 14600 26341 14603
rect 26108 14572 26341 14600
rect 26108 14560 26114 14572
rect 26329 14569 26341 14572
rect 26375 14569 26387 14603
rect 26329 14563 26387 14569
rect 4614 14492 4620 14544
rect 4672 14532 4678 14544
rect 11422 14532 11428 14544
rect 4672 14504 6132 14532
rect 11383 14504 11428 14532
rect 4672 14492 4678 14504
rect 1578 14464 1584 14476
rect 1491 14436 1584 14464
rect 1578 14424 1584 14436
rect 1636 14464 1642 14476
rect 2866 14464 2872 14476
rect 1636 14436 2872 14464
rect 1636 14424 1642 14436
rect 2866 14424 2872 14436
rect 2924 14464 2930 14476
rect 3786 14464 3792 14476
rect 2924 14436 3792 14464
rect 2924 14424 2930 14436
rect 3786 14424 3792 14436
rect 3844 14464 3850 14476
rect 4709 14467 4767 14473
rect 4709 14464 4721 14467
rect 3844 14436 4721 14464
rect 3844 14424 3850 14436
rect 4709 14433 4721 14436
rect 4755 14433 4767 14467
rect 4709 14427 4767 14433
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14396 4031 14399
rect 4062 14396 4068 14408
rect 4019 14368 4068 14396
rect 4019 14365 4031 14368
rect 3973 14359 4031 14365
rect 4062 14356 4068 14368
rect 4120 14396 4126 14408
rect 5074 14396 5080 14408
rect 4120 14368 5080 14396
rect 4120 14356 4126 14368
rect 5074 14356 5080 14368
rect 5132 14356 5138 14408
rect 5166 14356 5172 14408
rect 5224 14396 5230 14408
rect 6104 14405 6132 14504
rect 11422 14492 11428 14504
rect 11480 14492 11486 14544
rect 12158 14532 12164 14544
rect 11532 14504 12164 14532
rect 6638 14424 6644 14476
rect 6696 14464 6702 14476
rect 6733 14467 6791 14473
rect 6733 14464 6745 14467
rect 6696 14436 6745 14464
rect 6696 14424 6702 14436
rect 6733 14433 6745 14436
rect 6779 14433 6791 14467
rect 6733 14427 6791 14433
rect 7009 14467 7067 14473
rect 7009 14433 7021 14467
rect 7055 14464 7067 14467
rect 7098 14464 7104 14476
rect 7055 14436 7104 14464
rect 7055 14433 7067 14436
rect 7009 14427 7067 14433
rect 7098 14424 7104 14436
rect 7156 14424 7162 14476
rect 9030 14424 9036 14476
rect 9088 14464 9094 14476
rect 9125 14467 9183 14473
rect 9125 14464 9137 14467
rect 9088 14436 9137 14464
rect 9088 14424 9094 14436
rect 9125 14433 9137 14436
rect 9171 14464 9183 14467
rect 10594 14464 10600 14476
rect 9171 14436 10600 14464
rect 9171 14433 9183 14436
rect 9125 14427 9183 14433
rect 10594 14424 10600 14436
rect 10652 14424 10658 14476
rect 10873 14467 10931 14473
rect 10873 14433 10885 14467
rect 10919 14464 10931 14467
rect 11532 14464 11560 14504
rect 12158 14492 12164 14504
rect 12216 14492 12222 14544
rect 13262 14532 13268 14544
rect 12268 14504 13268 14532
rect 10919 14436 11560 14464
rect 10919 14433 10931 14436
rect 10873 14427 10931 14433
rect 6089 14399 6147 14405
rect 5224 14368 5672 14396
rect 5224 14356 5230 14368
rect 1857 14331 1915 14337
rect 1857 14297 1869 14331
rect 1903 14328 1915 14331
rect 1946 14328 1952 14340
rect 1903 14300 1952 14328
rect 1903 14297 1915 14300
rect 1857 14291 1915 14297
rect 1946 14288 1952 14300
rect 2004 14288 2010 14340
rect 3082 14300 3464 14328
rect 3436 14260 3464 14300
rect 3510 14288 3516 14340
rect 3568 14328 3574 14340
rect 5445 14331 5503 14337
rect 5445 14328 5457 14331
rect 3568 14300 5457 14328
rect 3568 14288 3574 14300
rect 5445 14297 5457 14300
rect 5491 14297 5503 14331
rect 5445 14291 5503 14297
rect 5258 14260 5264 14272
rect 3436 14232 5264 14260
rect 5258 14220 5264 14232
rect 5316 14220 5322 14272
rect 5644 14260 5672 14368
rect 6089 14365 6101 14399
rect 6135 14365 6147 14399
rect 11330 14396 11336 14408
rect 11291 14368 11336 14396
rect 6089 14359 6147 14365
rect 6104 14328 6132 14359
rect 11330 14356 11336 14368
rect 11388 14356 11394 14408
rect 11974 14396 11980 14408
rect 11887 14368 11980 14396
rect 11974 14356 11980 14368
rect 12032 14396 12038 14408
rect 12268 14396 12296 14504
rect 13262 14492 13268 14504
rect 13320 14492 13326 14544
rect 18690 14532 18696 14544
rect 15580 14504 18696 14532
rect 12526 14424 12532 14476
rect 12584 14464 12590 14476
rect 15580 14464 15608 14504
rect 18690 14492 18696 14504
rect 18748 14492 18754 14544
rect 19429 14535 19487 14541
rect 19429 14501 19441 14535
rect 19475 14501 19487 14535
rect 19429 14495 19487 14501
rect 12584 14436 15608 14464
rect 16761 14467 16819 14473
rect 12584 14424 12590 14436
rect 16761 14433 16773 14467
rect 16807 14464 16819 14467
rect 19444 14464 19472 14495
rect 21358 14492 21364 14544
rect 21416 14532 21422 14544
rect 21416 14504 31754 14532
rect 21416 14492 21422 14504
rect 25958 14464 25964 14476
rect 16807 14436 19472 14464
rect 25919 14436 25964 14464
rect 16807 14433 16819 14436
rect 16761 14427 16819 14433
rect 25958 14424 25964 14436
rect 26016 14424 26022 14476
rect 26142 14464 26148 14476
rect 26103 14436 26148 14464
rect 26142 14424 26148 14436
rect 26200 14424 26206 14476
rect 31726 14464 31754 14504
rect 37274 14464 37280 14476
rect 31726 14436 37280 14464
rect 37274 14424 37280 14436
rect 37332 14424 37338 14476
rect 12032 14368 12296 14396
rect 12032 14356 12038 14368
rect 12342 14356 12348 14408
rect 12400 14396 12406 14408
rect 13541 14399 13599 14405
rect 13541 14396 13553 14399
rect 12400 14368 13553 14396
rect 12400 14356 12406 14368
rect 13541 14365 13553 14368
rect 13587 14396 13599 14399
rect 14277 14399 14335 14405
rect 13587 14368 14228 14396
rect 13587 14365 13599 14368
rect 13541 14359 13599 14365
rect 7282 14328 7288 14340
rect 6104 14300 7288 14328
rect 7282 14288 7288 14300
rect 7340 14288 7346 14340
rect 7466 14288 7472 14340
rect 7524 14288 7530 14340
rect 8294 14288 8300 14340
rect 8352 14328 8358 14340
rect 13078 14328 13084 14340
rect 8352 14300 9890 14328
rect 11532 14300 13084 14328
rect 8352 14288 8358 14300
rect 7650 14260 7656 14272
rect 5644 14232 7656 14260
rect 7650 14220 7656 14232
rect 7708 14220 7714 14272
rect 8481 14263 8539 14269
rect 8481 14229 8493 14263
rect 8527 14260 8539 14263
rect 11532 14260 11560 14300
rect 13078 14288 13084 14300
rect 13136 14288 13142 14340
rect 8527 14232 11560 14260
rect 8527 14229 8539 14232
rect 8481 14223 8539 14229
rect 11606 14220 11612 14272
rect 11664 14260 11670 14272
rect 12069 14263 12127 14269
rect 12069 14260 12081 14263
rect 11664 14232 12081 14260
rect 11664 14220 11670 14232
rect 12069 14229 12081 14232
rect 12115 14229 12127 14263
rect 13630 14260 13636 14272
rect 13591 14232 13636 14260
rect 12069 14223 12127 14229
rect 13630 14220 13636 14232
rect 13688 14220 13694 14272
rect 14200 14260 14228 14368
rect 14277 14365 14289 14399
rect 14323 14365 14335 14399
rect 14277 14359 14335 14365
rect 16577 14399 16635 14405
rect 16577 14365 16589 14399
rect 16623 14365 16635 14399
rect 19610 14396 19616 14408
rect 19571 14368 19616 14396
rect 16577 14359 16635 14365
rect 14292 14328 14320 14359
rect 14550 14328 14556 14340
rect 14292 14300 14556 14328
rect 14550 14288 14556 14300
rect 14608 14288 14614 14340
rect 15010 14288 15016 14340
rect 15068 14288 15074 14340
rect 16592 14328 16620 14359
rect 19610 14356 19616 14368
rect 19668 14356 19674 14408
rect 21266 14396 21272 14408
rect 21227 14368 21272 14396
rect 21266 14356 21272 14368
rect 21324 14356 21330 14408
rect 22094 14356 22100 14408
rect 22152 14396 22158 14408
rect 22152 14368 22197 14396
rect 22152 14356 22158 14368
rect 22278 14356 22284 14408
rect 22336 14396 22342 14408
rect 24857 14399 24915 14405
rect 24857 14396 24869 14399
rect 22336 14368 24869 14396
rect 22336 14356 22342 14368
rect 24857 14365 24869 14368
rect 24903 14365 24915 14399
rect 24857 14359 24915 14365
rect 25041 14399 25099 14405
rect 25041 14365 25053 14399
rect 25087 14365 25099 14399
rect 27062 14396 27068 14408
rect 27023 14368 27068 14396
rect 25041 14359 25099 14365
rect 17770 14328 17776 14340
rect 16592 14300 17776 14328
rect 17770 14288 17776 14300
rect 17828 14288 17834 14340
rect 17865 14331 17923 14337
rect 17865 14297 17877 14331
rect 17911 14328 17923 14331
rect 18138 14328 18144 14340
rect 17911 14300 18144 14328
rect 17911 14297 17923 14300
rect 17865 14291 17923 14297
rect 18138 14288 18144 14300
rect 18196 14288 18202 14340
rect 18417 14331 18475 14337
rect 18417 14297 18429 14331
rect 18463 14328 18475 14331
rect 18966 14328 18972 14340
rect 18463 14300 18972 14328
rect 18463 14297 18475 14300
rect 18417 14291 18475 14297
rect 18966 14288 18972 14300
rect 19024 14328 19030 14340
rect 21634 14328 21640 14340
rect 19024 14300 21640 14328
rect 19024 14288 19030 14300
rect 21634 14288 21640 14300
rect 21692 14288 21698 14340
rect 25056 14328 25084 14359
rect 27062 14356 27068 14368
rect 27120 14356 27126 14408
rect 37918 14356 37924 14408
rect 37976 14396 37982 14408
rect 38013 14399 38071 14405
rect 38013 14396 38025 14399
rect 37976 14368 38025 14396
rect 37976 14356 37982 14368
rect 38013 14365 38025 14368
rect 38059 14365 38071 14399
rect 38013 14359 38071 14365
rect 27157 14331 27215 14337
rect 27157 14328 27169 14331
rect 25056 14300 27169 14328
rect 27157 14297 27169 14300
rect 27203 14297 27215 14331
rect 27157 14291 27215 14297
rect 16666 14260 16672 14272
rect 14200 14232 16672 14260
rect 16666 14220 16672 14232
rect 16724 14220 16730 14272
rect 17221 14263 17279 14269
rect 17221 14229 17233 14263
rect 17267 14260 17279 14263
rect 18046 14260 18052 14272
rect 17267 14232 18052 14260
rect 17267 14229 17279 14232
rect 17221 14223 17279 14229
rect 18046 14220 18052 14232
rect 18104 14220 18110 14272
rect 20438 14220 20444 14272
rect 20496 14260 20502 14272
rect 20625 14263 20683 14269
rect 20625 14260 20637 14263
rect 20496 14232 20637 14260
rect 20496 14220 20502 14232
rect 20625 14229 20637 14232
rect 20671 14229 20683 14263
rect 20625 14223 20683 14229
rect 20714 14220 20720 14272
rect 20772 14260 20778 14272
rect 21361 14263 21419 14269
rect 21361 14260 21373 14263
rect 20772 14232 21373 14260
rect 20772 14220 20778 14232
rect 21361 14229 21373 14232
rect 21407 14229 21419 14263
rect 38194 14260 38200 14272
rect 38155 14232 38200 14260
rect 21361 14223 21419 14229
rect 38194 14220 38200 14232
rect 38252 14220 38258 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 1765 14059 1823 14065
rect 1765 14025 1777 14059
rect 1811 14056 1823 14059
rect 2774 14056 2780 14068
rect 1811 14028 2780 14056
rect 1811 14025 1823 14028
rect 1765 14019 1823 14025
rect 2774 14016 2780 14028
rect 2832 14016 2838 14068
rect 4614 14056 4620 14068
rect 2884 14028 4620 14056
rect 2222 13988 2228 14000
rect 1596 13960 2228 13988
rect 1596 13929 1624 13960
rect 2222 13948 2228 13960
rect 2280 13948 2286 14000
rect 2314 13948 2320 14000
rect 2372 13988 2378 14000
rect 2884 13988 2912 14028
rect 4614 14016 4620 14028
rect 4672 14016 4678 14068
rect 5810 14056 5816 14068
rect 5771 14028 5816 14056
rect 5810 14016 5816 14028
rect 5868 14016 5874 14068
rect 6733 14059 6791 14065
rect 6733 14025 6745 14059
rect 6779 14056 6791 14059
rect 7006 14056 7012 14068
rect 6779 14028 7012 14056
rect 6779 14025 6791 14028
rect 6733 14019 6791 14025
rect 7006 14016 7012 14028
rect 7064 14016 7070 14068
rect 7374 14056 7380 14068
rect 7335 14028 7380 14056
rect 7374 14016 7380 14028
rect 7432 14016 7438 14068
rect 8021 14059 8079 14065
rect 8021 14025 8033 14059
rect 8067 14056 8079 14059
rect 8067 14028 10272 14056
rect 8067 14025 8079 14028
rect 8021 14019 8079 14025
rect 4706 13988 4712 14000
rect 2372 13960 2912 13988
rect 4370 13960 4712 13988
rect 2372 13948 2378 13960
rect 4706 13948 4712 13960
rect 4764 13948 4770 14000
rect 8846 13988 8852 14000
rect 8807 13960 8852 13988
rect 8846 13948 8852 13960
rect 8904 13948 8910 14000
rect 10244 13988 10272 14028
rect 10318 14016 10324 14068
rect 10376 14056 10382 14068
rect 10965 14059 11023 14065
rect 10376 14028 10421 14056
rect 10376 14016 10382 14028
rect 10965 14025 10977 14059
rect 11011 14056 11023 14059
rect 11514 14056 11520 14068
rect 11011 14028 11520 14056
rect 11011 14025 11023 14028
rect 10965 14019 11023 14025
rect 11514 14016 11520 14028
rect 11572 14016 11578 14068
rect 13906 14016 13912 14068
rect 13964 14056 13970 14068
rect 16942 14056 16948 14068
rect 13964 14028 16948 14056
rect 13964 14016 13970 14028
rect 16942 14016 16948 14028
rect 17000 14016 17006 14068
rect 18598 14056 18604 14068
rect 17512 14028 18604 14056
rect 13630 13988 13636 14000
rect 10244 13960 10456 13988
rect 13478 13960 13636 13988
rect 1581 13923 1639 13929
rect 1581 13889 1593 13923
rect 1627 13889 1639 13923
rect 2866 13920 2872 13932
rect 2827 13892 2872 13920
rect 1581 13883 1639 13889
rect 2866 13880 2872 13892
rect 2924 13880 2930 13932
rect 5074 13880 5080 13932
rect 5132 13920 5138 13932
rect 5721 13923 5779 13929
rect 5132 13892 5177 13920
rect 5132 13880 5138 13892
rect 5721 13889 5733 13923
rect 5767 13920 5779 13923
rect 5767 13892 6040 13920
rect 5767 13889 5779 13892
rect 5721 13883 5779 13889
rect 5169 13855 5227 13861
rect 5169 13821 5181 13855
rect 5215 13852 5227 13855
rect 5902 13852 5908 13864
rect 5215 13824 5908 13852
rect 5215 13821 5227 13824
rect 5169 13815 5227 13821
rect 5902 13812 5908 13824
rect 5960 13812 5966 13864
rect 6012 13784 6040 13892
rect 6086 13880 6092 13932
rect 6144 13920 6150 13932
rect 6641 13923 6699 13929
rect 6641 13920 6653 13923
rect 6144 13892 6653 13920
rect 6144 13880 6150 13892
rect 6641 13889 6653 13892
rect 6687 13889 6699 13923
rect 6641 13883 6699 13889
rect 6730 13880 6736 13932
rect 6788 13920 6794 13932
rect 7285 13923 7343 13929
rect 7285 13920 7297 13923
rect 6788 13892 7297 13920
rect 6788 13880 6794 13892
rect 7285 13889 7297 13892
rect 7331 13889 7343 13923
rect 7285 13883 7343 13889
rect 7650 13880 7656 13932
rect 7708 13920 7714 13932
rect 7929 13923 7987 13929
rect 7929 13920 7941 13923
rect 7708 13892 7941 13920
rect 7708 13880 7714 13892
rect 7929 13889 7941 13892
rect 7975 13889 7987 13923
rect 7929 13883 7987 13889
rect 9950 13880 9956 13932
rect 10008 13880 10014 13932
rect 6822 13812 6828 13864
rect 6880 13852 6886 13864
rect 8573 13855 8631 13861
rect 8573 13852 8585 13855
rect 6880 13824 8585 13852
rect 6880 13812 6886 13824
rect 8573 13821 8585 13824
rect 8619 13821 8631 13855
rect 8573 13815 8631 13821
rect 8846 13812 8852 13864
rect 8904 13852 8910 13864
rect 10428 13852 10456 13960
rect 13630 13948 13636 13960
rect 13688 13948 13694 14000
rect 14734 13988 14740 14000
rect 14695 13960 14740 13988
rect 14734 13948 14740 13960
rect 14792 13948 14798 14000
rect 15102 13948 15108 14000
rect 15160 13988 15166 14000
rect 15160 13960 16160 13988
rect 15160 13948 15166 13960
rect 10686 13880 10692 13932
rect 10744 13920 10750 13932
rect 10873 13923 10931 13929
rect 10873 13920 10885 13923
rect 10744 13892 10885 13920
rect 10744 13880 10750 13892
rect 10873 13889 10885 13892
rect 10919 13889 10931 13923
rect 10873 13883 10931 13889
rect 11698 13880 11704 13932
rect 11756 13920 11762 13932
rect 16132 13929 16160 13960
rect 16850 13948 16856 14000
rect 16908 13988 16914 14000
rect 17037 13991 17095 13997
rect 17037 13988 17049 13991
rect 16908 13960 17049 13988
rect 16908 13948 16914 13960
rect 17037 13957 17049 13960
rect 17083 13957 17095 13991
rect 17037 13951 17095 13957
rect 11977 13923 12035 13929
rect 11977 13920 11989 13923
rect 11756 13892 11989 13920
rect 11756 13880 11762 13892
rect 11977 13889 11989 13892
rect 12023 13889 12035 13923
rect 16117 13923 16175 13929
rect 11977 13883 12035 13889
rect 15580 13892 16068 13920
rect 12710 13852 12716 13864
rect 8904 13824 10180 13852
rect 10428 13824 12716 13852
rect 8904 13812 8910 13824
rect 7742 13784 7748 13796
rect 6012 13756 7748 13784
rect 7742 13744 7748 13756
rect 7800 13744 7806 13796
rect 8018 13744 8024 13796
rect 8076 13784 8082 13796
rect 10152 13784 10180 13824
rect 12710 13812 12716 13824
rect 12768 13812 12774 13864
rect 13446 13812 13452 13864
rect 13504 13852 13510 13864
rect 13725 13855 13783 13861
rect 13725 13852 13737 13855
rect 13504 13824 13737 13852
rect 13504 13812 13510 13824
rect 13725 13821 13737 13824
rect 13771 13821 13783 13855
rect 13725 13815 13783 13821
rect 14366 13812 14372 13864
rect 14424 13852 14430 13864
rect 14645 13855 14703 13861
rect 14645 13852 14657 13855
rect 14424 13824 14657 13852
rect 14424 13812 14430 13824
rect 14645 13821 14657 13824
rect 14691 13821 14703 13855
rect 14645 13815 14703 13821
rect 15194 13812 15200 13864
rect 15252 13852 15258 13864
rect 15580 13852 15608 13892
rect 15252 13824 15608 13852
rect 15657 13855 15715 13861
rect 15252 13812 15258 13824
rect 15657 13821 15669 13855
rect 15703 13852 15715 13855
rect 15930 13852 15936 13864
rect 15703 13824 15936 13852
rect 15703 13821 15715 13824
rect 15657 13815 15715 13821
rect 15930 13812 15936 13824
rect 15988 13812 15994 13864
rect 16040 13852 16068 13892
rect 16117 13889 16129 13923
rect 16163 13889 16175 13923
rect 16117 13883 16175 13889
rect 16666 13880 16672 13932
rect 16724 13920 16730 13932
rect 16945 13923 17003 13929
rect 16945 13920 16957 13923
rect 16724 13892 16957 13920
rect 16724 13880 16730 13892
rect 16945 13889 16957 13892
rect 16991 13920 17003 13923
rect 17512 13920 17540 14028
rect 18598 14016 18604 14028
rect 18656 14016 18662 14068
rect 20622 14056 20628 14068
rect 20272 14028 20628 14056
rect 17678 13988 17684 14000
rect 17639 13960 17684 13988
rect 17678 13948 17684 13960
rect 17736 13948 17742 14000
rect 17773 13991 17831 13997
rect 17773 13957 17785 13991
rect 17819 13988 17831 13991
rect 19797 13991 19855 13997
rect 19797 13988 19809 13991
rect 17819 13960 19809 13988
rect 17819 13957 17831 13960
rect 17773 13951 17831 13957
rect 19797 13957 19809 13960
rect 19843 13957 19855 13991
rect 19797 13951 19855 13957
rect 16991 13892 17540 13920
rect 18785 13923 18843 13929
rect 16991 13889 17003 13892
rect 16945 13883 17003 13889
rect 18785 13889 18797 13923
rect 18831 13920 18843 13923
rect 18874 13920 18880 13932
rect 18831 13892 18880 13920
rect 18831 13889 18843 13892
rect 18785 13883 18843 13889
rect 18874 13880 18880 13892
rect 18932 13880 18938 13932
rect 18966 13880 18972 13932
rect 19024 13920 19030 13932
rect 19061 13923 19119 13929
rect 19061 13920 19073 13923
rect 19024 13892 19073 13920
rect 19024 13880 19030 13892
rect 19061 13889 19073 13892
rect 19107 13889 19119 13923
rect 19061 13883 19119 13889
rect 19150 13880 19156 13932
rect 19208 13920 19214 13932
rect 19705 13923 19763 13929
rect 19705 13920 19717 13923
rect 19208 13892 19717 13920
rect 19208 13880 19214 13892
rect 19705 13889 19717 13892
rect 19751 13920 19763 13923
rect 20272 13920 20300 14028
rect 20622 14016 20628 14028
rect 20680 14016 20686 14068
rect 20438 13988 20444 14000
rect 20399 13960 20444 13988
rect 20438 13948 20444 13960
rect 20496 13948 20502 14000
rect 20533 13991 20591 13997
rect 20533 13957 20545 13991
rect 20579 13988 20591 13991
rect 20898 13988 20904 14000
rect 20579 13960 20904 13988
rect 20579 13957 20591 13960
rect 20533 13951 20591 13957
rect 20898 13948 20904 13960
rect 20956 13948 20962 14000
rect 21450 13988 21456 14000
rect 21411 13960 21456 13988
rect 21450 13948 21456 13960
rect 21508 13948 21514 14000
rect 19751 13892 20300 13920
rect 22005 13923 22063 13929
rect 19751 13889 19763 13892
rect 19705 13883 19763 13889
rect 22005 13889 22017 13923
rect 22051 13889 22063 13923
rect 22005 13883 22063 13889
rect 16040 13824 16896 13852
rect 11974 13784 11980 13796
rect 8076 13756 8708 13784
rect 10152 13756 11980 13784
rect 8076 13744 8082 13756
rect 3132 13719 3190 13725
rect 3132 13685 3144 13719
rect 3178 13716 3190 13719
rect 8570 13716 8576 13728
rect 3178 13688 8576 13716
rect 3178 13685 3190 13688
rect 3132 13679 3190 13685
rect 8570 13676 8576 13688
rect 8628 13676 8634 13728
rect 8680 13716 8708 13756
rect 11974 13744 11980 13756
rect 12032 13744 12038 13796
rect 16114 13784 16120 13796
rect 13556 13756 16120 13784
rect 10226 13716 10232 13728
rect 8680 13688 10232 13716
rect 10226 13676 10232 13688
rect 10284 13676 10290 13728
rect 12240 13719 12298 13725
rect 12240 13685 12252 13719
rect 12286 13716 12298 13719
rect 13556 13716 13584 13756
rect 16114 13744 16120 13756
rect 16172 13744 16178 13796
rect 16206 13744 16212 13796
rect 16264 13784 16270 13796
rect 16868 13784 16896 13824
rect 17144 13824 17724 13852
rect 17144 13784 17172 13824
rect 16264 13756 16309 13784
rect 16868 13756 17172 13784
rect 17696 13784 17724 13824
rect 17770 13812 17776 13864
rect 17828 13852 17834 13864
rect 17957 13855 18015 13861
rect 17957 13852 17969 13855
rect 17828 13824 17969 13852
rect 17828 13812 17834 13824
rect 17957 13821 17969 13824
rect 18003 13821 18015 13855
rect 21266 13852 21272 13864
rect 17957 13815 18015 13821
rect 18064 13824 21272 13852
rect 18064 13784 18092 13824
rect 21266 13812 21272 13824
rect 21324 13852 21330 13864
rect 22020 13852 22048 13883
rect 21324 13824 22048 13852
rect 21324 13812 21330 13824
rect 17696 13756 18092 13784
rect 16264 13744 16270 13756
rect 18230 13744 18236 13796
rect 18288 13784 18294 13796
rect 18690 13784 18696 13796
rect 18288 13756 18696 13784
rect 18288 13744 18294 13756
rect 18690 13744 18696 13756
rect 18748 13744 18754 13796
rect 12286 13688 13584 13716
rect 12286 13685 12298 13688
rect 12240 13679 12298 13685
rect 13630 13676 13636 13728
rect 13688 13716 13694 13728
rect 14642 13716 14648 13728
rect 13688 13688 14648 13716
rect 13688 13676 13694 13688
rect 14642 13676 14648 13688
rect 14700 13676 14706 13728
rect 16022 13676 16028 13728
rect 16080 13716 16086 13728
rect 20622 13716 20628 13728
rect 16080 13688 20628 13716
rect 16080 13676 16086 13688
rect 20622 13676 20628 13688
rect 20680 13676 20686 13728
rect 20990 13676 20996 13728
rect 21048 13716 21054 13728
rect 22097 13719 22155 13725
rect 22097 13716 22109 13719
rect 21048 13688 22109 13716
rect 21048 13676 21054 13688
rect 22097 13685 22109 13688
rect 22143 13685 22155 13719
rect 22097 13679 22155 13685
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 1302 13472 1308 13524
rect 1360 13512 1366 13524
rect 3329 13515 3387 13521
rect 3329 13512 3341 13515
rect 1360 13484 3341 13512
rect 1360 13472 1366 13484
rect 3329 13481 3341 13484
rect 3375 13481 3387 13515
rect 3329 13475 3387 13481
rect 3694 13472 3700 13524
rect 3752 13512 3758 13524
rect 6362 13512 6368 13524
rect 3752 13484 6368 13512
rect 3752 13472 3758 13484
rect 6362 13472 6368 13484
rect 6420 13472 6426 13524
rect 7926 13472 7932 13524
rect 7984 13512 7990 13524
rect 8113 13515 8171 13521
rect 8113 13512 8125 13515
rect 7984 13484 8125 13512
rect 7984 13472 7990 13484
rect 8113 13481 8125 13484
rect 8159 13481 8171 13515
rect 8113 13475 8171 13481
rect 9756 13515 9814 13521
rect 9756 13481 9768 13515
rect 9802 13512 9814 13515
rect 9802 13484 11836 13512
rect 9802 13481 9814 13484
rect 9756 13475 9814 13481
rect 3970 13444 3976 13456
rect 3436 13416 3976 13444
rect 1857 13379 1915 13385
rect 1857 13345 1869 13379
rect 1903 13376 1915 13379
rect 3436 13376 3464 13416
rect 3970 13404 3976 13416
rect 4028 13404 4034 13456
rect 5813 13447 5871 13453
rect 5813 13413 5825 13447
rect 5859 13444 5871 13447
rect 6270 13444 6276 13456
rect 5859 13416 6276 13444
rect 5859 13413 5871 13416
rect 5813 13407 5871 13413
rect 1903 13348 3464 13376
rect 1903 13345 1915 13348
rect 1857 13339 1915 13345
rect 3510 13336 3516 13388
rect 3568 13376 3574 13388
rect 5828 13376 5856 13407
rect 6270 13404 6276 13416
rect 6328 13404 6334 13456
rect 11238 13444 11244 13456
rect 11199 13416 11244 13444
rect 11238 13404 11244 13416
rect 11296 13404 11302 13456
rect 9493 13379 9551 13385
rect 9493 13376 9505 13379
rect 3568 13348 5856 13376
rect 6380 13348 9505 13376
rect 3568 13336 3574 13348
rect 6380 13320 6408 13348
rect 9493 13345 9505 13348
rect 9539 13376 9551 13379
rect 9766 13376 9772 13388
rect 9539 13348 9772 13376
rect 9539 13345 9551 13348
rect 9493 13339 9551 13345
rect 9766 13336 9772 13348
rect 9824 13376 9830 13388
rect 11701 13379 11759 13385
rect 11701 13376 11713 13379
rect 9824 13348 11713 13376
rect 9824 13336 9830 13348
rect 11701 13345 11713 13348
rect 11747 13345 11759 13379
rect 11808 13376 11836 13484
rect 11974 13472 11980 13524
rect 12032 13512 12038 13524
rect 12032 13484 13216 13512
rect 12032 13472 12038 13484
rect 12342 13376 12348 13388
rect 11808 13348 12348 13376
rect 11701 13339 11759 13345
rect 12342 13336 12348 13348
rect 12400 13336 12406 13388
rect 1578 13308 1584 13320
rect 1539 13280 1584 13308
rect 1578 13268 1584 13280
rect 1636 13268 1642 13320
rect 3786 13268 3792 13320
rect 3844 13308 3850 13320
rect 4065 13311 4123 13317
rect 4065 13308 4077 13311
rect 3844 13280 4077 13308
rect 3844 13268 3850 13280
rect 4065 13277 4077 13280
rect 4111 13277 4123 13311
rect 6362 13308 6368 13320
rect 6323 13280 6368 13308
rect 4065 13271 4123 13277
rect 6362 13268 6368 13280
rect 6420 13268 6426 13320
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 13188 13308 13216 13484
rect 16482 13472 16488 13524
rect 16540 13512 16546 13524
rect 16540 13484 20392 13512
rect 16540 13472 16546 13484
rect 13262 13404 13268 13456
rect 13320 13444 13326 13456
rect 20254 13444 20260 13456
rect 13320 13416 16896 13444
rect 13320 13404 13326 13416
rect 14550 13336 14556 13388
rect 14608 13376 14614 13388
rect 16577 13379 16635 13385
rect 16577 13376 16589 13379
rect 14608 13348 16589 13376
rect 14608 13336 14614 13348
rect 16577 13345 16589 13348
rect 16623 13345 16635 13379
rect 16577 13339 16635 13345
rect 11296 13280 11560 13308
rect 13188 13280 13860 13308
rect 11296 13268 11302 13280
rect 3970 13240 3976 13252
rect 3082 13212 3976 13240
rect 3970 13200 3976 13212
rect 4028 13200 4034 13252
rect 4338 13240 4344 13252
rect 4299 13212 4344 13240
rect 4338 13200 4344 13212
rect 4396 13200 4402 13252
rect 4798 13200 4804 13252
rect 4856 13200 4862 13252
rect 6641 13243 6699 13249
rect 6641 13209 6653 13243
rect 6687 13240 6699 13243
rect 6914 13240 6920 13252
rect 6687 13212 6920 13240
rect 6687 13209 6699 13212
rect 6641 13203 6699 13209
rect 6914 13200 6920 13212
rect 6972 13200 6978 13252
rect 7098 13200 7104 13252
rect 7156 13200 7162 13252
rect 11532 13240 11560 13280
rect 11977 13243 12035 13249
rect 11977 13240 11989 13243
rect 7944 13212 10258 13240
rect 11532 13212 11989 13240
rect 934 13132 940 13184
rect 992 13172 998 13184
rect 5626 13172 5632 13184
rect 992 13144 5632 13172
rect 992 13132 998 13144
rect 5626 13132 5632 13144
rect 5684 13132 5690 13184
rect 6454 13132 6460 13184
rect 6512 13172 6518 13184
rect 7944 13172 7972 13212
rect 11977 13209 11989 13212
rect 12023 13209 12035 13243
rect 13538 13240 13544 13252
rect 13202 13212 13544 13240
rect 11977 13203 12035 13209
rect 13538 13200 13544 13212
rect 13596 13200 13602 13252
rect 13630 13200 13636 13252
rect 13688 13240 13694 13252
rect 13725 13243 13783 13249
rect 13725 13240 13737 13243
rect 13688 13212 13737 13240
rect 13688 13200 13694 13212
rect 13725 13209 13737 13212
rect 13771 13209 13783 13243
rect 13832 13240 13860 13280
rect 15470 13268 15476 13320
rect 15528 13308 15534 13320
rect 16758 13308 16764 13320
rect 15528 13280 16764 13308
rect 15528 13268 15534 13280
rect 16758 13268 16764 13280
rect 16816 13268 16822 13320
rect 14366 13240 14372 13252
rect 13832 13212 14372 13240
rect 13725 13203 13783 13209
rect 14366 13200 14372 13212
rect 14424 13200 14430 13252
rect 14458 13200 14464 13252
rect 14516 13240 14522 13252
rect 14516 13212 14561 13240
rect 14516 13200 14522 13212
rect 14826 13200 14832 13252
rect 14884 13240 14890 13252
rect 15381 13243 15439 13249
rect 15381 13240 15393 13243
rect 14884 13212 15393 13240
rect 14884 13200 14890 13212
rect 15381 13209 15393 13212
rect 15427 13209 15439 13243
rect 15381 13203 15439 13209
rect 15841 13243 15899 13249
rect 15841 13209 15853 13243
rect 15887 13209 15899 13243
rect 16868 13240 16896 13416
rect 18432 13416 20260 13444
rect 16942 13268 16948 13320
rect 17000 13308 17006 13320
rect 17221 13311 17279 13317
rect 17221 13308 17233 13311
rect 17000 13280 17233 13308
rect 17000 13268 17006 13280
rect 17221 13277 17233 13280
rect 17267 13308 17279 13311
rect 17310 13308 17316 13320
rect 17267 13280 17316 13308
rect 17267 13277 17279 13280
rect 17221 13271 17279 13277
rect 17310 13268 17316 13280
rect 17368 13268 17374 13320
rect 18432 13308 18460 13416
rect 20254 13404 20260 13416
rect 20312 13404 20318 13456
rect 20364 13444 20392 13484
rect 20622 13472 20628 13524
rect 20680 13512 20686 13524
rect 20717 13515 20775 13521
rect 20717 13512 20729 13515
rect 20680 13484 20729 13512
rect 20680 13472 20686 13484
rect 20717 13481 20729 13484
rect 20763 13481 20775 13515
rect 20717 13475 20775 13481
rect 22189 13515 22247 13521
rect 22189 13481 22201 13515
rect 22235 13512 22247 13515
rect 22278 13512 22284 13524
rect 22235 13484 22284 13512
rect 22235 13481 22247 13484
rect 22189 13475 22247 13481
rect 22278 13472 22284 13484
rect 22336 13472 22342 13524
rect 37642 13512 37648 13524
rect 25332 13484 37648 13512
rect 20364 13416 20668 13444
rect 18782 13336 18788 13388
rect 18840 13376 18846 13388
rect 19886 13376 19892 13388
rect 18840 13348 19892 13376
rect 18840 13336 18846 13348
rect 19886 13336 19892 13348
rect 19944 13336 19950 13388
rect 18601 13311 18659 13317
rect 18601 13308 18613 13311
rect 18432 13280 18613 13308
rect 18601 13277 18613 13280
rect 18647 13277 18659 13311
rect 18601 13271 18659 13277
rect 18690 13268 18696 13320
rect 18748 13308 18754 13320
rect 20640 13317 20668 13416
rect 20625 13311 20683 13317
rect 18748 13280 18793 13308
rect 18748 13268 18754 13280
rect 20625 13277 20637 13311
rect 20671 13277 20683 13311
rect 20625 13271 20683 13277
rect 22094 13268 22100 13320
rect 22152 13308 22158 13320
rect 25332 13308 25360 13484
rect 37642 13472 37648 13484
rect 37700 13472 37706 13524
rect 26418 13444 26424 13456
rect 26379 13416 26424 13444
rect 26418 13404 26424 13416
rect 26476 13404 26482 13456
rect 26050 13376 26056 13388
rect 26011 13348 26056 13376
rect 26050 13336 26056 13348
rect 26108 13336 26114 13388
rect 22152 13280 25360 13308
rect 26237 13311 26295 13317
rect 22152 13268 22158 13280
rect 26237 13277 26249 13311
rect 26283 13308 26295 13311
rect 27522 13308 27528 13320
rect 26283 13280 27528 13308
rect 26283 13277 26295 13280
rect 26237 13271 26295 13277
rect 27522 13268 27528 13280
rect 27580 13268 27586 13320
rect 30374 13268 30380 13320
rect 30432 13308 30438 13320
rect 34333 13311 34391 13317
rect 34333 13308 34345 13311
rect 30432 13280 34345 13308
rect 30432 13268 30438 13280
rect 34333 13277 34345 13280
rect 34379 13277 34391 13311
rect 34333 13271 34391 13277
rect 37274 13268 37280 13320
rect 37332 13308 37338 13320
rect 38013 13311 38071 13317
rect 38013 13308 38025 13311
rect 37332 13280 38025 13308
rect 37332 13268 37338 13280
rect 38013 13277 38025 13280
rect 38059 13277 38071 13311
rect 38013 13271 38071 13277
rect 18049 13243 18107 13249
rect 18049 13240 18061 13243
rect 16868 13212 18061 13240
rect 15841 13203 15899 13209
rect 18049 13209 18061 13212
rect 18095 13240 18107 13243
rect 19150 13240 19156 13252
rect 18095 13212 19156 13240
rect 18095 13209 18107 13212
rect 18049 13203 18107 13209
rect 6512 13144 7972 13172
rect 6512 13132 6518 13144
rect 11054 13132 11060 13184
rect 11112 13172 11118 13184
rect 15856 13172 15884 13203
rect 19150 13200 19156 13212
rect 19208 13200 19214 13252
rect 19518 13240 19524 13252
rect 19479 13212 19524 13240
rect 19518 13200 19524 13212
rect 19576 13200 19582 13252
rect 19613 13243 19671 13249
rect 19613 13209 19625 13243
rect 19659 13209 19671 13243
rect 19613 13203 19671 13209
rect 20165 13243 20223 13249
rect 20165 13209 20177 13243
rect 20211 13240 20223 13243
rect 20438 13240 20444 13252
rect 20211 13212 20444 13240
rect 20211 13209 20223 13212
rect 20165 13203 20223 13209
rect 16666 13172 16672 13184
rect 11112 13144 16672 13172
rect 11112 13132 11118 13144
rect 16666 13132 16672 13144
rect 16724 13132 16730 13184
rect 17954 13132 17960 13184
rect 18012 13172 18018 13184
rect 18782 13172 18788 13184
rect 18012 13144 18788 13172
rect 18012 13132 18018 13144
rect 18782 13132 18788 13144
rect 18840 13132 18846 13184
rect 19628 13172 19656 13203
rect 20438 13200 20444 13212
rect 20496 13200 20502 13252
rect 20990 13240 20996 13252
rect 20640 13212 20996 13240
rect 20640 13172 20668 13212
rect 20990 13200 20996 13212
rect 21048 13200 21054 13252
rect 19628 13144 20668 13172
rect 21266 13132 21272 13184
rect 21324 13172 21330 13184
rect 27706 13172 27712 13184
rect 21324 13144 27712 13172
rect 21324 13132 21330 13144
rect 27706 13132 27712 13144
rect 27764 13132 27770 13184
rect 34149 13175 34207 13181
rect 34149 13141 34161 13175
rect 34195 13172 34207 13175
rect 36906 13172 36912 13184
rect 34195 13144 36912 13172
rect 34195 13141 34207 13144
rect 34149 13135 34207 13141
rect 36906 13132 36912 13144
rect 36964 13132 36970 13184
rect 38194 13172 38200 13184
rect 38155 13144 38200 13172
rect 38194 13132 38200 13144
rect 38252 13132 38258 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 658 12928 664 12980
rect 716 12968 722 12980
rect 4798 12968 4804 12980
rect 716 12940 4804 12968
rect 716 12928 722 12940
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 5902 12928 5908 12980
rect 5960 12968 5966 12980
rect 9217 12971 9275 12977
rect 5960 12940 7604 12968
rect 5960 12928 5966 12940
rect 2866 12860 2872 12912
rect 2924 12860 2930 12912
rect 3418 12860 3424 12912
rect 3476 12900 3482 12912
rect 3476 12872 4646 12900
rect 3476 12860 3482 12872
rect 6362 12860 6368 12912
rect 6420 12900 6426 12912
rect 7576 12900 7604 12940
rect 9217 12937 9229 12971
rect 9263 12968 9275 12971
rect 9263 12940 10824 12968
rect 9263 12937 9275 12940
rect 9217 12931 9275 12937
rect 6420 12872 7512 12900
rect 7576 12872 8234 12900
rect 6420 12860 6426 12872
rect 3881 12835 3939 12841
rect 3881 12832 3893 12835
rect 3620 12804 3893 12832
rect 1578 12764 1584 12776
rect 1539 12736 1584 12764
rect 1578 12724 1584 12736
rect 1636 12724 1642 12776
rect 1857 12767 1915 12773
rect 1857 12733 1869 12767
rect 1903 12764 1915 12767
rect 3510 12764 3516 12776
rect 1903 12736 3516 12764
rect 1903 12733 1915 12736
rect 1857 12727 1915 12733
rect 3510 12724 3516 12736
rect 3568 12724 3574 12776
rect 3234 12656 3240 12708
rect 3292 12696 3298 12708
rect 3329 12699 3387 12705
rect 3329 12696 3341 12699
rect 3292 12668 3341 12696
rect 3292 12656 3298 12668
rect 3329 12665 3341 12668
rect 3375 12665 3387 12699
rect 3329 12659 3387 12665
rect 3620 12628 3648 12804
rect 3881 12801 3893 12804
rect 3927 12801 3939 12835
rect 3881 12795 3939 12801
rect 5626 12792 5632 12844
rect 5684 12832 5690 12844
rect 7484 12841 7512 12872
rect 9766 12860 9772 12912
rect 9824 12900 9830 12912
rect 10597 12903 10655 12909
rect 10597 12900 10609 12903
rect 9824 12872 10609 12900
rect 9824 12860 9830 12872
rect 10597 12869 10609 12872
rect 10643 12869 10655 12903
rect 10796 12900 10824 12940
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 20070 12968 20076 12980
rect 12492 12940 17356 12968
rect 12492 12928 12498 12940
rect 17328 12912 17356 12940
rect 17420 12940 20076 12968
rect 13078 12900 13084 12912
rect 10796 12872 13084 12900
rect 10597 12863 10655 12869
rect 13078 12860 13084 12872
rect 13136 12860 13142 12912
rect 13446 12900 13452 12912
rect 13280 12872 13452 12900
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 5684 12804 6561 12832
rect 5684 12792 5690 12804
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 7469 12835 7527 12841
rect 7469 12801 7481 12835
rect 7515 12801 7527 12835
rect 7469 12795 7527 12801
rect 9674 12792 9680 12844
rect 9732 12832 9738 12844
rect 9861 12835 9919 12841
rect 9861 12832 9873 12835
rect 9732 12804 9873 12832
rect 9732 12792 9738 12804
rect 9861 12801 9873 12804
rect 9907 12832 9919 12835
rect 11054 12832 11060 12844
rect 9907 12804 11060 12832
rect 9907 12801 9919 12804
rect 9861 12795 9919 12801
rect 11054 12792 11060 12804
rect 11112 12792 11118 12844
rect 11330 12792 11336 12844
rect 11388 12832 11394 12844
rect 11701 12835 11759 12841
rect 11701 12832 11713 12835
rect 11388 12804 11713 12832
rect 11388 12792 11394 12804
rect 11701 12801 11713 12804
rect 11747 12801 11759 12835
rect 12618 12832 12624 12844
rect 12579 12804 12624 12832
rect 11701 12795 11759 12801
rect 12618 12792 12624 12804
rect 12676 12792 12682 12844
rect 12986 12792 12992 12844
rect 13044 12832 13050 12844
rect 13280 12841 13308 12872
rect 13446 12860 13452 12872
rect 13504 12860 13510 12912
rect 15470 12900 15476 12912
rect 14766 12872 15476 12900
rect 15470 12860 15476 12872
rect 15528 12860 15534 12912
rect 15654 12900 15660 12912
rect 15615 12872 15660 12900
rect 15654 12860 15660 12872
rect 15712 12860 15718 12912
rect 15749 12903 15807 12909
rect 15749 12869 15761 12903
rect 15795 12900 15807 12903
rect 17126 12900 17132 12912
rect 15795 12872 17132 12900
rect 15795 12869 15807 12872
rect 15749 12863 15807 12869
rect 17126 12860 17132 12872
rect 17184 12860 17190 12912
rect 17310 12900 17316 12912
rect 17223 12872 17316 12900
rect 17310 12860 17316 12872
rect 17368 12860 17374 12912
rect 13265 12835 13323 12841
rect 13044 12804 13216 12832
rect 13044 12792 13050 12804
rect 3694 12724 3700 12776
rect 3752 12764 3758 12776
rect 4157 12767 4215 12773
rect 4157 12764 4169 12767
rect 3752 12736 4169 12764
rect 3752 12724 3758 12736
rect 4157 12733 4169 12736
rect 4203 12733 4215 12767
rect 4157 12727 4215 12733
rect 4246 12724 4252 12776
rect 4304 12764 4310 12776
rect 7745 12767 7803 12773
rect 4304 12736 6868 12764
rect 4304 12724 4310 12736
rect 5626 12696 5632 12708
rect 5587 12668 5632 12696
rect 5626 12656 5632 12668
rect 5684 12656 5690 12708
rect 4614 12628 4620 12640
rect 3620 12600 4620 12628
rect 4614 12588 4620 12600
rect 4672 12588 4678 12640
rect 5166 12588 5172 12640
rect 5224 12628 5230 12640
rect 6733 12631 6791 12637
rect 6733 12628 6745 12631
rect 5224 12600 6745 12628
rect 5224 12588 5230 12600
rect 6733 12597 6745 12600
rect 6779 12597 6791 12631
rect 6840 12628 6868 12736
rect 7745 12733 7757 12767
rect 7791 12764 7803 12767
rect 10318 12764 10324 12776
rect 7791 12736 10324 12764
rect 7791 12733 7803 12736
rect 7745 12727 7803 12733
rect 10318 12724 10324 12736
rect 10376 12724 10382 12776
rect 10410 12724 10416 12776
rect 10468 12764 10474 12776
rect 11974 12764 11980 12776
rect 10468 12736 11980 12764
rect 10468 12724 10474 12736
rect 11974 12724 11980 12736
rect 12032 12724 12038 12776
rect 13188 12764 13216 12804
rect 13265 12801 13277 12835
rect 13311 12801 13323 12835
rect 13265 12795 13323 12801
rect 14826 12792 14832 12844
rect 14884 12832 14890 12844
rect 15286 12832 15292 12844
rect 14884 12804 15292 12832
rect 14884 12792 14890 12804
rect 15286 12792 15292 12804
rect 15344 12792 15350 12844
rect 16942 12832 16948 12844
rect 16903 12804 16948 12832
rect 16942 12792 16948 12804
rect 17000 12792 17006 12844
rect 13541 12767 13599 12773
rect 13541 12764 13553 12767
rect 13188 12736 13553 12764
rect 13541 12733 13553 12736
rect 13587 12733 13599 12767
rect 13541 12727 13599 12733
rect 13630 12724 13636 12776
rect 13688 12764 13694 12776
rect 16114 12764 16120 12776
rect 13688 12736 16120 12764
rect 13688 12724 13694 12736
rect 16114 12724 16120 12736
rect 16172 12724 16178 12776
rect 16301 12767 16359 12773
rect 16301 12733 16313 12767
rect 16347 12764 16359 12767
rect 17310 12764 17316 12776
rect 16347 12736 17316 12764
rect 16347 12733 16359 12736
rect 16301 12727 16359 12733
rect 17310 12724 17316 12736
rect 17368 12724 17374 12776
rect 11882 12696 11888 12708
rect 10521 12668 11888 12696
rect 10226 12628 10232 12640
rect 6840 12600 10232 12628
rect 6733 12591 6791 12597
rect 10226 12588 10232 12600
rect 10284 12588 10290 12640
rect 10318 12588 10324 12640
rect 10376 12628 10382 12640
rect 10521 12628 10549 12668
rect 11882 12656 11888 12668
rect 11940 12696 11946 12708
rect 11940 12668 13400 12696
rect 11940 12656 11946 12668
rect 11790 12628 11796 12640
rect 10376 12600 10549 12628
rect 11751 12600 11796 12628
rect 10376 12588 10382 12600
rect 11790 12588 11796 12600
rect 11848 12588 11854 12640
rect 11974 12588 11980 12640
rect 12032 12628 12038 12640
rect 12618 12628 12624 12640
rect 12032 12600 12624 12628
rect 12032 12588 12038 12600
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 12713 12631 12771 12637
rect 12713 12597 12725 12631
rect 12759 12628 12771 12631
rect 13262 12628 13268 12640
rect 12759 12600 13268 12628
rect 12759 12597 12771 12600
rect 12713 12591 12771 12597
rect 13262 12588 13268 12600
rect 13320 12588 13326 12640
rect 13372 12628 13400 12668
rect 16206 12656 16212 12708
rect 16264 12696 16270 12708
rect 17420 12696 17448 12940
rect 20070 12928 20076 12940
rect 20128 12928 20134 12980
rect 20898 12968 20904 12980
rect 20272 12940 20760 12968
rect 20859 12940 20904 12968
rect 17586 12860 17592 12912
rect 17644 12900 17650 12912
rect 17770 12900 17776 12912
rect 17644 12872 17776 12900
rect 17644 12860 17650 12872
rect 17770 12860 17776 12872
rect 17828 12860 17834 12912
rect 18141 12903 18199 12909
rect 18141 12900 18153 12903
rect 17972 12872 18153 12900
rect 16264 12668 17448 12696
rect 17972 12696 18000 12872
rect 18141 12869 18153 12872
rect 18187 12869 18199 12903
rect 18141 12863 18199 12869
rect 18233 12903 18291 12909
rect 18233 12869 18245 12903
rect 18279 12900 18291 12903
rect 18414 12900 18420 12912
rect 18279 12872 18420 12900
rect 18279 12869 18291 12872
rect 18233 12863 18291 12869
rect 18414 12860 18420 12872
rect 18472 12860 18478 12912
rect 19797 12903 19855 12909
rect 19797 12869 19809 12903
rect 19843 12900 19855 12903
rect 20272 12900 20300 12940
rect 19843 12872 20300 12900
rect 20732 12900 20760 12940
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 27522 12968 27528 12980
rect 27483 12940 27528 12968
rect 27522 12928 27528 12940
rect 27580 12928 27586 12980
rect 22094 12900 22100 12912
rect 20732 12872 22100 12900
rect 19843 12869 19855 12872
rect 19797 12863 19855 12869
rect 22094 12860 22100 12872
rect 22152 12860 22158 12912
rect 22373 12903 22431 12909
rect 22373 12869 22385 12903
rect 22419 12900 22431 12903
rect 22830 12900 22836 12912
rect 22419 12872 22836 12900
rect 22419 12869 22431 12872
rect 22373 12863 22431 12869
rect 22830 12860 22836 12872
rect 22888 12860 22894 12912
rect 20809 12835 20867 12841
rect 20809 12801 20821 12835
rect 20855 12801 20867 12835
rect 20809 12795 20867 12801
rect 22189 12835 22247 12841
rect 22189 12801 22201 12835
rect 22235 12832 22247 12835
rect 23566 12832 23572 12844
rect 22235 12804 23572 12832
rect 22235 12801 22247 12804
rect 22189 12795 22247 12801
rect 18414 12764 18420 12776
rect 18375 12736 18420 12764
rect 18414 12724 18420 12736
rect 18472 12724 18478 12776
rect 19518 12724 19524 12776
rect 19576 12764 19582 12776
rect 19705 12767 19763 12773
rect 19705 12764 19717 12767
rect 19576 12736 19717 12764
rect 19576 12724 19582 12736
rect 19705 12733 19717 12736
rect 19751 12733 19763 12767
rect 19705 12727 19763 12733
rect 20349 12767 20407 12773
rect 20349 12733 20361 12767
rect 20395 12764 20407 12767
rect 20438 12764 20444 12776
rect 20395 12736 20444 12764
rect 20395 12733 20407 12736
rect 20349 12727 20407 12733
rect 20438 12724 20444 12736
rect 20496 12724 20502 12776
rect 19886 12696 19892 12708
rect 17972 12668 19892 12696
rect 16264 12656 16270 12668
rect 19886 12656 19892 12668
rect 19944 12656 19950 12708
rect 20070 12656 20076 12708
rect 20128 12696 20134 12708
rect 20824 12696 20852 12795
rect 23566 12792 23572 12804
rect 23624 12792 23630 12844
rect 27709 12835 27767 12841
rect 27709 12801 27721 12835
rect 27755 12832 27767 12835
rect 28350 12832 28356 12844
rect 27755 12804 28212 12832
rect 28311 12804 28356 12832
rect 27755 12801 27767 12804
rect 27709 12795 27767 12801
rect 22646 12696 22652 12708
rect 20128 12668 20852 12696
rect 22066 12668 22652 12696
rect 20128 12656 20134 12668
rect 15013 12631 15071 12637
rect 15013 12628 15025 12631
rect 13372 12600 15025 12628
rect 15013 12597 15025 12600
rect 15059 12597 15071 12631
rect 15013 12591 15071 12597
rect 15930 12588 15936 12640
rect 15988 12628 15994 12640
rect 18414 12628 18420 12640
rect 15988 12600 18420 12628
rect 15988 12588 15994 12600
rect 18414 12588 18420 12600
rect 18472 12588 18478 12640
rect 18598 12588 18604 12640
rect 18656 12628 18662 12640
rect 22066 12628 22094 12668
rect 22646 12656 22652 12668
rect 22704 12656 22710 12708
rect 28184 12705 28212 12804
rect 28350 12792 28356 12804
rect 28408 12792 28414 12844
rect 38102 12832 38108 12844
rect 38063 12804 38108 12832
rect 38102 12792 38108 12804
rect 38160 12792 38166 12844
rect 28169 12699 28227 12705
rect 28169 12665 28181 12699
rect 28215 12665 28227 12699
rect 28169 12659 28227 12665
rect 38194 12628 38200 12640
rect 18656 12600 22094 12628
rect 38155 12600 38200 12628
rect 18656 12588 18662 12600
rect 38194 12588 38200 12600
rect 38252 12588 38258 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 1026 12384 1032 12436
rect 1084 12424 1090 12436
rect 3510 12424 3516 12436
rect 1084 12396 3516 12424
rect 1084 12384 1090 12396
rect 3510 12384 3516 12396
rect 3568 12424 3574 12436
rect 3568 12396 3648 12424
rect 3568 12384 3574 12396
rect 3234 12316 3240 12368
rect 3292 12356 3298 12368
rect 3329 12359 3387 12365
rect 3329 12356 3341 12359
rect 3292 12328 3341 12356
rect 3292 12316 3298 12328
rect 3329 12325 3341 12328
rect 3375 12325 3387 12359
rect 3620 12356 3648 12396
rect 3694 12384 3700 12436
rect 3752 12424 3758 12436
rect 5166 12424 5172 12436
rect 3752 12396 5172 12424
rect 3752 12384 3758 12396
rect 5166 12384 5172 12396
rect 5224 12384 5230 12436
rect 7285 12427 7343 12433
rect 7285 12393 7297 12427
rect 7331 12424 7343 12427
rect 7742 12424 7748 12436
rect 7331 12396 7748 12424
rect 7331 12393 7343 12396
rect 7285 12387 7343 12393
rect 7742 12384 7748 12396
rect 7800 12384 7806 12436
rect 8938 12384 8944 12436
rect 8996 12424 9002 12436
rect 9217 12427 9275 12433
rect 9217 12424 9229 12427
rect 8996 12396 9229 12424
rect 8996 12384 9002 12396
rect 9217 12393 9229 12396
rect 9263 12393 9275 12427
rect 9217 12387 9275 12393
rect 9306 12384 9312 12436
rect 9364 12424 9370 12436
rect 11517 12427 11575 12433
rect 11517 12424 11529 12427
rect 9364 12396 11529 12424
rect 9364 12384 9370 12396
rect 11517 12393 11529 12396
rect 11563 12393 11575 12427
rect 11517 12387 11575 12393
rect 12240 12427 12298 12433
rect 12240 12393 12252 12427
rect 12286 12424 12298 12427
rect 12286 12396 13492 12424
rect 12286 12393 12298 12396
rect 12240 12387 12298 12393
rect 3970 12356 3976 12368
rect 3620 12328 3976 12356
rect 3329 12319 3387 12325
rect 3970 12316 3976 12328
rect 4028 12316 4034 12368
rect 7558 12316 7564 12368
rect 7616 12356 7622 12368
rect 7929 12359 7987 12365
rect 7929 12356 7941 12359
rect 7616 12328 7941 12356
rect 7616 12316 7622 12328
rect 7929 12325 7941 12328
rect 7975 12325 7987 12359
rect 13464 12356 13492 12396
rect 13538 12384 13544 12436
rect 13596 12424 13602 12436
rect 13725 12427 13783 12433
rect 13725 12424 13737 12427
rect 13596 12396 13737 12424
rect 13596 12384 13602 12396
rect 13725 12393 13737 12396
rect 13771 12393 13783 12427
rect 16025 12427 16083 12433
rect 16025 12424 16037 12427
rect 13725 12387 13783 12393
rect 14384 12396 16037 12424
rect 14384 12356 14412 12396
rect 16025 12393 16037 12396
rect 16071 12424 16083 12427
rect 16206 12424 16212 12436
rect 16071 12396 16212 12424
rect 16071 12393 16083 12396
rect 16025 12387 16083 12393
rect 16206 12384 16212 12396
rect 16264 12384 16270 12436
rect 16574 12384 16580 12436
rect 16632 12424 16638 12436
rect 16850 12424 16856 12436
rect 16632 12396 16856 12424
rect 16632 12384 16638 12396
rect 16850 12384 16856 12396
rect 16908 12424 16914 12436
rect 18598 12424 18604 12436
rect 16908 12396 18604 12424
rect 16908 12384 16914 12396
rect 18598 12384 18604 12396
rect 18656 12384 18662 12436
rect 19426 12384 19432 12436
rect 19484 12424 19490 12436
rect 20438 12424 20444 12436
rect 19484 12396 20444 12424
rect 19484 12384 19490 12396
rect 20438 12384 20444 12396
rect 20496 12384 20502 12436
rect 13464 12328 14412 12356
rect 7929 12319 7987 12325
rect 15654 12316 15660 12368
rect 15712 12356 15718 12368
rect 15712 12328 24992 12356
rect 15712 12316 15718 12328
rect 1394 12248 1400 12300
rect 1452 12288 1458 12300
rect 1857 12291 1915 12297
rect 1857 12288 1869 12291
rect 1452 12260 1869 12288
rect 1452 12248 1458 12260
rect 1857 12257 1869 12260
rect 1903 12257 1915 12291
rect 1857 12251 1915 12257
rect 3786 12248 3792 12300
rect 3844 12288 3850 12300
rect 4709 12291 4767 12297
rect 4709 12288 4721 12291
rect 3844 12260 4721 12288
rect 3844 12248 3850 12260
rect 4709 12257 4721 12260
rect 4755 12257 4767 12291
rect 4709 12251 4767 12257
rect 5537 12291 5595 12297
rect 5537 12257 5549 12291
rect 5583 12288 5595 12291
rect 6270 12288 6276 12300
rect 5583 12260 6276 12288
rect 5583 12257 5595 12260
rect 5537 12251 5595 12257
rect 1578 12220 1584 12232
rect 1539 12192 1584 12220
rect 1578 12180 1584 12192
rect 1636 12180 1642 12232
rect 4614 12180 4620 12232
rect 4672 12220 4678 12232
rect 5552 12220 5580 12251
rect 6270 12248 6276 12260
rect 6328 12248 6334 12300
rect 11606 12288 11612 12300
rect 7760 12260 11612 12288
rect 7760 12220 7788 12260
rect 11606 12248 11612 12260
rect 11664 12248 11670 12300
rect 11698 12248 11704 12300
rect 11756 12288 11762 12300
rect 11977 12291 12035 12297
rect 11977 12288 11989 12291
rect 11756 12260 11989 12288
rect 11756 12248 11762 12260
rect 11977 12257 11989 12260
rect 12023 12288 12035 12291
rect 12986 12288 12992 12300
rect 12023 12260 12992 12288
rect 12023 12257 12035 12260
rect 11977 12251 12035 12257
rect 12986 12248 12992 12260
rect 13044 12288 13050 12300
rect 13446 12288 13452 12300
rect 13044 12260 13452 12288
rect 13044 12248 13050 12260
rect 13446 12248 13452 12260
rect 13504 12288 13510 12300
rect 14277 12291 14335 12297
rect 14277 12288 14289 12291
rect 13504 12260 14289 12288
rect 13504 12248 13510 12260
rect 14277 12257 14289 12260
rect 14323 12288 14335 12291
rect 14550 12288 14556 12300
rect 14323 12260 14556 12288
rect 14323 12257 14335 12260
rect 14277 12251 14335 12257
rect 14550 12248 14556 12260
rect 14608 12248 14614 12300
rect 16577 12291 16635 12297
rect 16577 12257 16589 12291
rect 16623 12288 16635 12291
rect 17034 12288 17040 12300
rect 16623 12260 17040 12288
rect 16623 12257 16635 12260
rect 16577 12251 16635 12257
rect 17034 12248 17040 12260
rect 17092 12248 17098 12300
rect 17773 12291 17831 12297
rect 17773 12257 17785 12291
rect 17819 12288 17831 12291
rect 19518 12288 19524 12300
rect 17819 12260 19524 12288
rect 17819 12257 17831 12260
rect 17773 12251 17831 12257
rect 19518 12248 19524 12260
rect 19576 12248 19582 12300
rect 20901 12291 20959 12297
rect 20901 12288 20913 12291
rect 19628 12260 20913 12288
rect 4672 12192 5580 12220
rect 6946 12192 7788 12220
rect 4672 12180 4678 12192
rect 7834 12180 7840 12232
rect 7892 12220 7898 12232
rect 8202 12220 8208 12232
rect 7892 12192 8208 12220
rect 7892 12180 7898 12192
rect 8202 12180 8208 12192
rect 8260 12180 8266 12232
rect 8662 12180 8668 12232
rect 8720 12220 8726 12232
rect 9030 12220 9036 12232
rect 8720 12192 9036 12220
rect 8720 12180 8726 12192
rect 9030 12180 9036 12192
rect 9088 12220 9094 12232
rect 9125 12223 9183 12229
rect 9125 12220 9137 12223
rect 9088 12192 9137 12220
rect 9088 12180 9094 12192
rect 9125 12189 9137 12192
rect 9171 12189 9183 12223
rect 9125 12183 9183 12189
rect 9674 12180 9680 12232
rect 9732 12220 9738 12232
rect 9769 12223 9827 12229
rect 9769 12220 9781 12223
rect 9732 12192 9781 12220
rect 9732 12180 9738 12192
rect 9769 12189 9781 12192
rect 9815 12189 9827 12223
rect 19426 12220 19432 12232
rect 19387 12192 19432 12220
rect 9769 12183 9827 12189
rect 19426 12180 19432 12192
rect 19484 12180 19490 12232
rect 3142 12152 3148 12164
rect 3082 12124 3148 12152
rect 3142 12112 3148 12124
rect 3200 12112 3206 12164
rect 3973 12155 4031 12161
rect 3973 12121 3985 12155
rect 4019 12152 4031 12155
rect 4062 12152 4068 12164
rect 4019 12124 4068 12152
rect 4019 12121 4031 12124
rect 3973 12115 4031 12121
rect 4062 12112 4068 12124
rect 4120 12112 4126 12164
rect 5813 12155 5871 12161
rect 5813 12121 5825 12155
rect 5859 12121 5871 12155
rect 5813 12115 5871 12121
rect 2774 12044 2780 12096
rect 2832 12084 2838 12096
rect 3234 12084 3240 12096
rect 2832 12056 3240 12084
rect 2832 12044 2838 12056
rect 3234 12044 3240 12056
rect 3292 12044 3298 12096
rect 4154 12044 4160 12096
rect 4212 12084 4218 12096
rect 4982 12084 4988 12096
rect 4212 12056 4988 12084
rect 4212 12044 4218 12056
rect 4982 12044 4988 12056
rect 5040 12044 5046 12096
rect 5828 12084 5856 12115
rect 7742 12112 7748 12164
rect 7800 12152 7806 12164
rect 9490 12152 9496 12164
rect 7800 12124 9496 12152
rect 7800 12112 7806 12124
rect 9490 12112 9496 12124
rect 9548 12112 9554 12164
rect 10045 12155 10103 12161
rect 10045 12121 10057 12155
rect 10091 12121 10103 12155
rect 11790 12152 11796 12164
rect 11270 12124 11796 12152
rect 10045 12115 10103 12121
rect 7926 12084 7932 12096
rect 5828 12056 7932 12084
rect 7926 12044 7932 12056
rect 7984 12044 7990 12096
rect 9858 12044 9864 12096
rect 9916 12084 9922 12096
rect 10060 12084 10088 12115
rect 11790 12112 11796 12124
rect 11848 12112 11854 12164
rect 12526 12112 12532 12164
rect 12584 12152 12590 12164
rect 14550 12152 14556 12164
rect 12584 12124 12742 12152
rect 14511 12124 14556 12152
rect 12584 12112 12590 12124
rect 14550 12112 14556 12124
rect 14608 12112 14614 12164
rect 16574 12152 16580 12164
rect 15778 12124 16580 12152
rect 16574 12112 16580 12124
rect 16632 12112 16638 12164
rect 16669 12155 16727 12161
rect 16669 12121 16681 12155
rect 16715 12121 16727 12155
rect 17218 12152 17224 12164
rect 17179 12124 17224 12152
rect 16669 12115 16727 12121
rect 10962 12084 10968 12096
rect 9916 12056 10968 12084
rect 9916 12044 9922 12056
rect 10962 12044 10968 12056
rect 11020 12044 11026 12096
rect 11514 12044 11520 12096
rect 11572 12084 11578 12096
rect 13078 12084 13084 12096
rect 11572 12056 13084 12084
rect 11572 12044 11578 12056
rect 13078 12044 13084 12056
rect 13136 12044 13142 12096
rect 13262 12044 13268 12096
rect 13320 12084 13326 12096
rect 15562 12084 15568 12096
rect 13320 12056 15568 12084
rect 13320 12044 13326 12056
rect 15562 12044 15568 12056
rect 15620 12044 15626 12096
rect 16114 12044 16120 12096
rect 16172 12084 16178 12096
rect 16684 12084 16712 12115
rect 17218 12112 17224 12124
rect 17276 12112 17282 12164
rect 17862 12112 17868 12164
rect 17920 12152 17926 12164
rect 18414 12152 18420 12164
rect 17920 12124 17965 12152
rect 18375 12124 18420 12152
rect 17920 12112 17926 12124
rect 18414 12112 18420 12124
rect 18472 12112 18478 12164
rect 18598 12112 18604 12164
rect 18656 12152 18662 12164
rect 19628 12152 19656 12260
rect 20901 12257 20913 12260
rect 20947 12257 20959 12291
rect 20901 12251 20959 12257
rect 24486 12248 24492 12300
rect 24544 12288 24550 12300
rect 24857 12291 24915 12297
rect 24857 12288 24869 12291
rect 24544 12260 24869 12288
rect 24544 12248 24550 12260
rect 24857 12257 24869 12260
rect 24903 12257 24915 12291
rect 24857 12251 24915 12257
rect 22002 12180 22008 12232
rect 22060 12220 22066 12232
rect 22097 12223 22155 12229
rect 22097 12220 22109 12223
rect 22060 12192 22109 12220
rect 22060 12180 22066 12192
rect 22097 12189 22109 12192
rect 22143 12189 22155 12223
rect 24964 12220 24992 12328
rect 25041 12291 25099 12297
rect 25041 12257 25053 12291
rect 25087 12288 25099 12291
rect 26973 12291 27031 12297
rect 26973 12288 26985 12291
rect 25087 12260 26985 12288
rect 25087 12257 25099 12260
rect 25041 12251 25099 12257
rect 26973 12257 26985 12260
rect 27019 12257 27031 12291
rect 26973 12251 27031 12257
rect 26881 12223 26939 12229
rect 26881 12220 26893 12223
rect 24964 12192 26893 12220
rect 22097 12183 22155 12189
rect 26881 12189 26893 12192
rect 26927 12220 26939 12223
rect 28350 12220 28356 12232
rect 26927 12192 28356 12220
rect 26927 12189 26939 12192
rect 26881 12183 26939 12189
rect 28350 12180 28356 12192
rect 28408 12180 28414 12232
rect 18656 12124 19656 12152
rect 18656 12112 18662 12124
rect 19886 12112 19892 12164
rect 19944 12152 19950 12164
rect 20622 12152 20628 12164
rect 19944 12124 20628 12152
rect 19944 12112 19950 12124
rect 20622 12112 20628 12124
rect 20680 12112 20686 12164
rect 20717 12155 20775 12161
rect 20717 12121 20729 12155
rect 20763 12152 20775 12155
rect 22554 12152 22560 12164
rect 20763 12124 22560 12152
rect 20763 12121 20775 12124
rect 20717 12115 20775 12121
rect 22554 12112 22560 12124
rect 22612 12112 22618 12164
rect 16172 12056 16712 12084
rect 16172 12044 16178 12056
rect 16758 12044 16764 12096
rect 16816 12084 16822 12096
rect 21266 12084 21272 12096
rect 16816 12056 21272 12084
rect 16816 12044 16822 12056
rect 21266 12044 21272 12056
rect 21324 12044 21330 12096
rect 21818 12044 21824 12096
rect 21876 12084 21882 12096
rect 22189 12087 22247 12093
rect 22189 12084 22201 12087
rect 21876 12056 22201 12084
rect 21876 12044 21882 12056
rect 22189 12053 22201 12056
rect 22235 12053 22247 12087
rect 22189 12047 22247 12053
rect 25501 12087 25559 12093
rect 25501 12053 25513 12087
rect 25547 12084 25559 12087
rect 26234 12084 26240 12096
rect 25547 12056 26240 12084
rect 25547 12053 25559 12056
rect 25501 12047 25559 12053
rect 26234 12044 26240 12056
rect 26292 12044 26298 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 3786 11880 3792 11892
rect 2056 11852 3792 11880
rect 1578 11704 1584 11756
rect 1636 11744 1642 11756
rect 2056 11753 2084 11852
rect 3786 11840 3792 11852
rect 3844 11840 3850 11892
rect 4798 11880 4804 11892
rect 4172 11852 4804 11880
rect 4172 11812 4200 11852
rect 4798 11840 4804 11852
rect 4856 11840 4862 11892
rect 6641 11883 6699 11889
rect 6641 11849 6653 11883
rect 6687 11880 6699 11883
rect 7006 11880 7012 11892
rect 6687 11852 7012 11880
rect 6687 11849 6699 11852
rect 6641 11843 6699 11849
rect 7006 11840 7012 11852
rect 7064 11840 7070 11892
rect 9950 11880 9956 11892
rect 7484 11852 9956 11880
rect 4614 11812 4620 11824
rect 3542 11784 4200 11812
rect 4264 11784 4620 11812
rect 4264 11753 4292 11784
rect 4614 11772 4620 11784
rect 4672 11772 4678 11824
rect 6822 11812 6828 11824
rect 5750 11784 6828 11812
rect 6822 11772 6828 11784
rect 6880 11772 6886 11824
rect 7484 11821 7512 11852
rect 9950 11840 9956 11852
rect 10008 11840 10014 11892
rect 12434 11880 12440 11892
rect 11348 11852 12440 11880
rect 7469 11815 7527 11821
rect 7469 11781 7481 11815
rect 7515 11781 7527 11815
rect 9214 11812 9220 11824
rect 8694 11784 9220 11812
rect 7469 11775 7527 11781
rect 9214 11772 9220 11784
rect 9272 11772 9278 11824
rect 9674 11812 9680 11824
rect 9416 11784 9680 11812
rect 2041 11747 2099 11753
rect 2041 11744 2053 11747
rect 1636 11716 2053 11744
rect 1636 11704 1642 11716
rect 2041 11713 2053 11716
rect 2087 11713 2099 11747
rect 2041 11707 2099 11713
rect 4249 11747 4307 11753
rect 4249 11713 4261 11747
rect 4295 11713 4307 11747
rect 4249 11707 4307 11713
rect 6454 11704 6460 11756
rect 6512 11744 6518 11756
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 6512 11716 6561 11744
rect 6512 11704 6518 11716
rect 6549 11713 6561 11716
rect 6595 11744 6607 11747
rect 6638 11744 6644 11756
rect 6595 11716 6644 11744
rect 6595 11713 6607 11716
rect 6549 11707 6607 11713
rect 6638 11704 6644 11716
rect 6696 11704 6702 11756
rect 9416 11753 9444 11784
rect 9674 11772 9680 11784
rect 9732 11772 9738 11824
rect 10134 11772 10140 11824
rect 10192 11772 10198 11824
rect 9401 11747 9459 11753
rect 9401 11713 9413 11747
rect 9447 11713 9459 11747
rect 9401 11707 9459 11713
rect 2317 11679 2375 11685
rect 2317 11645 2329 11679
rect 2363 11676 2375 11679
rect 4154 11676 4160 11688
rect 2363 11648 4160 11676
rect 2363 11645 2375 11648
rect 2317 11639 2375 11645
rect 4154 11636 4160 11648
rect 4212 11636 4218 11688
rect 4525 11679 4583 11685
rect 4525 11645 4537 11679
rect 4571 11676 4583 11679
rect 5534 11676 5540 11688
rect 4571 11648 5540 11676
rect 4571 11645 4583 11648
rect 4525 11639 4583 11645
rect 5534 11636 5540 11648
rect 5592 11636 5598 11688
rect 5810 11636 5816 11688
rect 5868 11676 5874 11688
rect 6086 11676 6092 11688
rect 5868 11648 6092 11676
rect 5868 11636 5874 11648
rect 6086 11636 6092 11648
rect 6144 11636 6150 11688
rect 7098 11636 7104 11688
rect 7156 11676 7162 11688
rect 7193 11679 7251 11685
rect 7193 11676 7205 11679
rect 7156 11648 7205 11676
rect 7156 11636 7162 11648
rect 7193 11645 7205 11648
rect 7239 11645 7251 11679
rect 7193 11639 7251 11645
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11676 9735 11679
rect 11348 11676 11376 11852
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 12912 11852 13124 11880
rect 11606 11772 11612 11824
rect 11664 11812 11670 11824
rect 12912 11812 12940 11852
rect 11664 11784 12296 11812
rect 11664 11772 11670 11784
rect 11701 11747 11759 11753
rect 11701 11713 11713 11747
rect 11747 11744 11759 11747
rect 11790 11744 11796 11756
rect 11747 11716 11796 11744
rect 11747 11713 11759 11716
rect 11701 11707 11759 11713
rect 11790 11704 11796 11716
rect 11848 11744 11854 11756
rect 12158 11744 12164 11756
rect 11848 11716 12164 11744
rect 11848 11704 11854 11716
rect 12158 11704 12164 11716
rect 12216 11704 12222 11756
rect 12268 11744 12296 11784
rect 12452 11784 12940 11812
rect 13096 11812 13124 11852
rect 13262 11840 13268 11892
rect 13320 11880 13326 11892
rect 13320 11852 16436 11880
rect 13320 11840 13326 11852
rect 13096 11784 13754 11812
rect 12452 11753 12480 11784
rect 14826 11772 14832 11824
rect 14884 11812 14890 11824
rect 15013 11815 15071 11821
rect 15013 11812 15025 11815
rect 14884 11784 15025 11812
rect 14884 11772 14890 11784
rect 15013 11781 15025 11784
rect 15059 11781 15071 11815
rect 15654 11812 15660 11824
rect 15013 11775 15071 11781
rect 15113 11784 15660 11812
rect 12345 11747 12403 11753
rect 12345 11744 12357 11747
rect 12268 11716 12357 11744
rect 12345 11713 12357 11716
rect 12391 11713 12403 11747
rect 12345 11707 12403 11713
rect 12437 11747 12495 11753
rect 12437 11713 12449 11747
rect 12483 11713 12495 11747
rect 12986 11744 12992 11756
rect 12947 11716 12992 11744
rect 12437 11707 12495 11713
rect 12986 11704 12992 11716
rect 13044 11704 13050 11756
rect 9723 11648 11376 11676
rect 9723 11645 9735 11648
rect 9677 11639 9735 11645
rect 12710 11636 12716 11688
rect 12768 11676 12774 11688
rect 13265 11679 13323 11685
rect 13265 11676 13277 11679
rect 12768 11648 13277 11676
rect 12768 11636 12774 11648
rect 13265 11645 13277 11648
rect 13311 11676 13323 11679
rect 15113 11676 15141 11784
rect 15654 11772 15660 11784
rect 15712 11772 15718 11824
rect 15749 11815 15807 11821
rect 15749 11781 15761 11815
rect 15795 11812 15807 11815
rect 16022 11812 16028 11824
rect 15795 11784 16028 11812
rect 15795 11781 15807 11784
rect 15749 11775 15807 11781
rect 16022 11772 16028 11784
rect 16080 11772 16086 11824
rect 16298 11812 16304 11824
rect 16259 11784 16304 11812
rect 16298 11772 16304 11784
rect 16356 11772 16362 11824
rect 16408 11812 16436 11852
rect 16574 11840 16580 11892
rect 16632 11880 16638 11892
rect 16632 11852 18184 11880
rect 16632 11840 16638 11852
rect 16758 11812 16764 11824
rect 16408 11784 16764 11812
rect 16758 11772 16764 11784
rect 16816 11772 16822 11824
rect 16942 11772 16948 11824
rect 17000 11812 17006 11824
rect 17037 11815 17095 11821
rect 17037 11812 17049 11815
rect 17000 11784 17049 11812
rect 17000 11772 17006 11784
rect 17037 11781 17049 11784
rect 17083 11781 17095 11815
rect 17586 11812 17592 11824
rect 17547 11784 17592 11812
rect 17037 11775 17095 11781
rect 17586 11772 17592 11784
rect 17644 11772 17650 11824
rect 18156 11812 18184 11852
rect 20438 11840 20444 11892
rect 20496 11880 20502 11892
rect 20533 11883 20591 11889
rect 20533 11880 20545 11883
rect 20496 11852 20545 11880
rect 20496 11840 20502 11852
rect 20533 11849 20545 11852
rect 20579 11849 20591 11883
rect 20533 11843 20591 11849
rect 23014 11840 23020 11892
rect 23072 11880 23078 11892
rect 28718 11880 28724 11892
rect 23072 11852 28724 11880
rect 23072 11840 23078 11852
rect 28718 11840 28724 11852
rect 28776 11840 28782 11892
rect 21177 11815 21235 11821
rect 21177 11812 21189 11815
rect 18156 11784 21189 11812
rect 21177 11781 21189 11784
rect 21223 11781 21235 11815
rect 21177 11775 21235 11781
rect 21266 11772 21272 11824
rect 21324 11812 21330 11824
rect 22189 11815 22247 11821
rect 22189 11812 22201 11815
rect 21324 11784 22201 11812
rect 21324 11772 21330 11784
rect 22189 11781 22201 11784
rect 22235 11781 22247 11815
rect 22189 11775 22247 11781
rect 18049 11747 18107 11753
rect 18049 11713 18061 11747
rect 18095 11744 18107 11747
rect 18969 11747 19027 11753
rect 18969 11744 18981 11747
rect 18095 11716 18981 11744
rect 18095 11713 18107 11716
rect 18049 11707 18107 11713
rect 18969 11713 18981 11716
rect 19015 11713 19027 11747
rect 20441 11747 20499 11753
rect 20441 11744 20453 11747
rect 18969 11707 19027 11713
rect 19076 11716 20453 11744
rect 13311 11648 15141 11676
rect 13311 11645 13323 11648
rect 13265 11639 13323 11645
rect 15654 11636 15660 11688
rect 15712 11676 15718 11688
rect 16574 11676 16580 11688
rect 15712 11648 16580 11676
rect 15712 11636 15718 11648
rect 16574 11636 16580 11648
rect 16632 11636 16638 11688
rect 16945 11679 17003 11685
rect 16945 11645 16957 11679
rect 16991 11645 17003 11679
rect 16945 11639 17003 11645
rect 9398 11608 9404 11620
rect 8496 11580 9404 11608
rect 1854 11500 1860 11552
rect 1912 11540 1918 11552
rect 3789 11543 3847 11549
rect 3789 11540 3801 11543
rect 1912 11512 3801 11540
rect 1912 11500 1918 11512
rect 3789 11509 3801 11512
rect 3835 11509 3847 11543
rect 3789 11503 3847 11509
rect 5997 11543 6055 11549
rect 5997 11509 6009 11543
rect 6043 11540 6055 11543
rect 6086 11540 6092 11552
rect 6043 11512 6092 11540
rect 6043 11509 6055 11512
rect 5997 11503 6055 11509
rect 6086 11500 6092 11512
rect 6144 11540 6150 11552
rect 8496 11540 8524 11580
rect 9398 11568 9404 11580
rect 9456 11568 9462 11620
rect 11149 11611 11207 11617
rect 11149 11577 11161 11611
rect 11195 11608 11207 11611
rect 12158 11608 12164 11620
rect 11195 11580 12164 11608
rect 11195 11577 11207 11580
rect 11149 11571 11207 11577
rect 12158 11568 12164 11580
rect 12216 11568 12222 11620
rect 14642 11568 14648 11620
rect 14700 11608 14706 11620
rect 16960 11608 16988 11639
rect 17034 11636 17040 11688
rect 17092 11676 17098 11688
rect 17862 11676 17868 11688
rect 17092 11648 17868 11676
rect 17092 11636 17098 11648
rect 17862 11636 17868 11648
rect 17920 11676 17926 11688
rect 18064 11676 18092 11707
rect 17920 11648 18092 11676
rect 18233 11679 18291 11685
rect 17920 11636 17926 11648
rect 18233 11645 18245 11679
rect 18279 11645 18291 11679
rect 18233 11639 18291 11645
rect 14700 11580 16988 11608
rect 14700 11568 14706 11580
rect 18248 11552 18276 11639
rect 18598 11636 18604 11688
rect 18656 11676 18662 11688
rect 19076 11676 19104 11716
rect 20441 11713 20453 11716
rect 20487 11713 20499 11747
rect 20441 11707 20499 11713
rect 21085 11747 21143 11753
rect 21085 11713 21097 11747
rect 21131 11713 21143 11747
rect 23566 11744 23572 11756
rect 23479 11716 23572 11744
rect 21085 11707 21143 11713
rect 18656 11648 19104 11676
rect 19153 11679 19211 11685
rect 18656 11636 18662 11648
rect 19153 11645 19165 11679
rect 19199 11645 19211 11679
rect 19153 11639 19211 11645
rect 18690 11568 18696 11620
rect 18748 11608 18754 11620
rect 19168 11608 19196 11639
rect 19242 11636 19248 11688
rect 19300 11676 19306 11688
rect 21100 11676 21128 11707
rect 23566 11704 23572 11716
rect 23624 11744 23630 11756
rect 24118 11744 24124 11756
rect 23624 11716 24124 11744
rect 23624 11704 23630 11716
rect 24118 11704 24124 11716
rect 24176 11704 24182 11756
rect 21174 11676 21180 11688
rect 19300 11648 21180 11676
rect 19300 11636 19306 11648
rect 21174 11636 21180 11648
rect 21232 11636 21238 11688
rect 22097 11679 22155 11685
rect 22097 11645 22109 11679
rect 22143 11676 22155 11679
rect 22278 11676 22284 11688
rect 22143 11648 22284 11676
rect 22143 11645 22155 11648
rect 22097 11639 22155 11645
rect 22278 11636 22284 11648
rect 22336 11636 22342 11688
rect 22370 11636 22376 11688
rect 22428 11676 22434 11688
rect 22428 11648 22473 11676
rect 22428 11636 22434 11648
rect 18748 11580 19196 11608
rect 18748 11568 18754 11580
rect 20622 11568 20628 11620
rect 20680 11608 20686 11620
rect 25958 11608 25964 11620
rect 20680 11580 25964 11608
rect 20680 11568 20686 11580
rect 25958 11568 25964 11580
rect 26016 11568 26022 11620
rect 8938 11540 8944 11552
rect 6144 11512 8524 11540
rect 8899 11512 8944 11540
rect 6144 11500 6150 11512
rect 8938 11500 8944 11512
rect 8996 11500 9002 11552
rect 9490 11500 9496 11552
rect 9548 11540 9554 11552
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 9548 11512 11805 11540
rect 9548 11500 9554 11512
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 18230 11540 18236 11552
rect 18143 11512 18236 11540
rect 11793 11503 11851 11509
rect 18230 11500 18236 11512
rect 18288 11540 18294 11552
rect 21266 11540 21272 11552
rect 18288 11512 21272 11540
rect 18288 11500 18294 11512
rect 21266 11500 21272 11512
rect 21324 11500 21330 11552
rect 21726 11500 21732 11552
rect 21784 11540 21790 11552
rect 23198 11540 23204 11552
rect 21784 11512 23204 11540
rect 21784 11500 21790 11512
rect 23198 11500 23204 11512
rect 23256 11500 23262 11552
rect 23658 11540 23664 11552
rect 23619 11512 23664 11540
rect 23658 11500 23664 11512
rect 23716 11500 23722 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 3329 11339 3387 11345
rect 3329 11305 3341 11339
rect 3375 11336 3387 11339
rect 3418 11336 3424 11348
rect 3375 11308 3424 11336
rect 3375 11305 3387 11308
rect 3329 11299 3387 11305
rect 3418 11296 3424 11308
rect 3476 11296 3482 11348
rect 4604 11339 4662 11345
rect 4604 11305 4616 11339
rect 4650 11336 4662 11339
rect 5994 11336 6000 11348
rect 4650 11308 6000 11336
rect 4650 11305 4662 11308
rect 4604 11299 4662 11305
rect 5994 11296 6000 11308
rect 6052 11296 6058 11348
rect 6638 11296 6644 11348
rect 6696 11336 6702 11348
rect 6812 11339 6870 11345
rect 6812 11336 6824 11339
rect 6696 11308 6824 11336
rect 6696 11296 6702 11308
rect 6812 11305 6824 11308
rect 6858 11336 6870 11339
rect 8294 11336 8300 11348
rect 6858 11308 8300 11336
rect 6858 11305 6870 11308
rect 6812 11299 6870 11305
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 9214 11336 9220 11348
rect 9175 11308 9220 11336
rect 9214 11296 9220 11308
rect 9272 11296 9278 11348
rect 11606 11336 11612 11348
rect 9324 11308 11612 11336
rect 8938 11268 8944 11280
rect 7852 11240 8944 11268
rect 1578 11200 1584 11212
rect 1539 11172 1584 11200
rect 1578 11160 1584 11172
rect 1636 11160 1642 11212
rect 1857 11203 1915 11209
rect 1857 11169 1869 11203
rect 1903 11200 1915 11203
rect 2314 11200 2320 11212
rect 1903 11172 2320 11200
rect 1903 11169 1915 11172
rect 1857 11163 1915 11169
rect 2314 11160 2320 11172
rect 2372 11160 2378 11212
rect 4341 11203 4399 11209
rect 4341 11169 4353 11203
rect 4387 11200 4399 11203
rect 4614 11200 4620 11212
rect 4387 11172 4620 11200
rect 4387 11169 4399 11172
rect 4341 11163 4399 11169
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 6270 11160 6276 11212
rect 6328 11200 6334 11212
rect 6549 11203 6607 11209
rect 6549 11200 6561 11203
rect 6328 11172 6561 11200
rect 6328 11160 6334 11172
rect 6549 11169 6561 11172
rect 6595 11200 6607 11203
rect 6914 11200 6920 11212
rect 6595 11172 6920 11200
rect 6595 11169 6607 11172
rect 6549 11163 6607 11169
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 7282 11160 7288 11212
rect 7340 11200 7346 11212
rect 7852 11200 7880 11240
rect 8938 11228 8944 11240
rect 8996 11228 9002 11280
rect 9324 11200 9352 11308
rect 11606 11296 11612 11308
rect 11664 11296 11670 11348
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 14182 11336 14188 11348
rect 12492 11308 14188 11336
rect 12492 11296 12498 11308
rect 14182 11296 14188 11308
rect 14240 11296 14246 11348
rect 14550 11336 14556 11348
rect 14384 11308 14556 11336
rect 9766 11268 9772 11280
rect 7340 11172 7880 11200
rect 7944 11172 9352 11200
rect 9600 11240 9772 11268
rect 7340 11160 7346 11172
rect 7944 11118 7972 11172
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11132 9183 11135
rect 9600 11132 9628 11240
rect 9766 11228 9772 11240
rect 9824 11228 9830 11280
rect 11514 11268 11520 11280
rect 11475 11240 11520 11268
rect 11514 11228 11520 11240
rect 11572 11228 11578 11280
rect 13725 11271 13783 11277
rect 13725 11237 13737 11271
rect 13771 11268 13783 11271
rect 14384 11268 14412 11308
rect 14550 11296 14556 11308
rect 14608 11296 14614 11348
rect 15562 11296 15568 11348
rect 15620 11336 15626 11348
rect 16025 11339 16083 11345
rect 16025 11336 16037 11339
rect 15620 11308 16037 11336
rect 15620 11296 15626 11308
rect 16025 11305 16037 11308
rect 16071 11305 16083 11339
rect 16025 11299 16083 11305
rect 16132 11308 20852 11336
rect 13771 11240 14412 11268
rect 13771 11237 13783 11240
rect 13725 11231 13783 11237
rect 15746 11228 15752 11280
rect 15804 11268 15810 11280
rect 16132 11268 16160 11308
rect 18230 11268 18236 11280
rect 15804 11240 16160 11268
rect 16684 11240 18236 11268
rect 15804 11228 15810 11240
rect 11974 11200 11980 11212
rect 9784 11172 11980 11200
rect 9784 11144 9812 11172
rect 11974 11160 11980 11172
rect 12032 11160 12038 11212
rect 12250 11160 12256 11212
rect 12308 11200 12314 11212
rect 16684 11209 16712 11240
rect 18230 11228 18236 11240
rect 18288 11228 18294 11280
rect 18414 11228 18420 11280
rect 18472 11268 18478 11280
rect 20073 11271 20131 11277
rect 20073 11268 20085 11271
rect 18472 11240 20085 11268
rect 18472 11228 18478 11240
rect 20073 11237 20085 11240
rect 20119 11237 20131 11271
rect 20073 11231 20131 11237
rect 16669 11203 16727 11209
rect 12308 11172 15700 11200
rect 12308 11160 12314 11172
rect 9766 11132 9772 11144
rect 9171 11104 9628 11132
rect 9727 11104 9772 11132
rect 9171 11101 9183 11104
rect 9125 11095 9183 11101
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 14274 11132 14280 11144
rect 14235 11104 14280 11132
rect 14274 11092 14280 11104
rect 14332 11092 14338 11144
rect 15672 11118 15700 11172
rect 16669 11169 16681 11203
rect 16715 11169 16727 11203
rect 16669 11163 16727 11169
rect 17681 11203 17739 11209
rect 17681 11169 17693 11203
rect 17727 11200 17739 11203
rect 17954 11200 17960 11212
rect 17727 11172 17960 11200
rect 17727 11169 17739 11172
rect 17681 11163 17739 11169
rect 17954 11160 17960 11172
rect 18012 11160 18018 11212
rect 19334 11200 19340 11212
rect 18156 11172 19340 11200
rect 17862 11092 17868 11144
rect 17920 11132 17926 11144
rect 18156 11141 18184 11172
rect 19334 11160 19340 11172
rect 19392 11160 19398 11212
rect 19610 11160 19616 11212
rect 19668 11200 19674 11212
rect 20714 11200 20720 11212
rect 19668 11172 20720 11200
rect 19668 11160 19674 11172
rect 20714 11160 20720 11172
rect 20772 11160 20778 11212
rect 18141 11135 18199 11141
rect 18141 11132 18153 11135
rect 17920 11104 18153 11132
rect 17920 11092 17926 11104
rect 18141 11101 18153 11104
rect 18187 11101 18199 11135
rect 19058 11132 19064 11144
rect 18141 11095 18199 11101
rect 18340 11104 19064 11132
rect 4890 11064 4896 11076
rect 3082 11036 4896 11064
rect 4890 11024 4896 11036
rect 4948 11024 4954 11076
rect 5994 11064 6000 11076
rect 5842 11036 6000 11064
rect 5994 11024 6000 11036
rect 6052 11024 6058 11076
rect 8573 11067 8631 11073
rect 8573 11033 8585 11067
rect 8619 11064 8631 11067
rect 9030 11064 9036 11076
rect 8619 11036 9036 11064
rect 8619 11033 8631 11036
rect 8573 11027 8631 11033
rect 9030 11024 9036 11036
rect 9088 11064 9094 11076
rect 10042 11064 10048 11076
rect 9088 11036 9904 11064
rect 10003 11036 10048 11064
rect 9088 11024 9094 11036
rect 5350 10956 5356 11008
rect 5408 10996 5414 11008
rect 6089 10999 6147 11005
rect 6089 10996 6101 10999
rect 5408 10968 6101 10996
rect 5408 10956 5414 10968
rect 6089 10965 6101 10968
rect 6135 10996 6147 10999
rect 6730 10996 6736 11008
rect 6135 10968 6736 10996
rect 6135 10965 6147 10968
rect 6089 10959 6147 10965
rect 6730 10956 6736 10968
rect 6788 10956 6794 11008
rect 9876 10996 9904 11036
rect 10042 11024 10048 11036
rect 10100 11024 10106 11076
rect 12158 11064 12164 11076
rect 11270 11036 12164 11064
rect 12158 11024 12164 11036
rect 12216 11024 12222 11076
rect 12253 11067 12311 11073
rect 12253 11033 12265 11067
rect 12299 11064 12311 11067
rect 12342 11064 12348 11076
rect 12299 11036 12348 11064
rect 12299 11033 12311 11036
rect 12253 11027 12311 11033
rect 12342 11024 12348 11036
rect 12400 11024 12406 11076
rect 13538 11064 13544 11076
rect 13478 11036 13544 11064
rect 13538 11024 13544 11036
rect 13596 11024 13602 11076
rect 14182 11024 14188 11076
rect 14240 11064 14246 11076
rect 14553 11067 14611 11073
rect 14553 11064 14565 11067
rect 14240 11036 14565 11064
rect 14240 11024 14246 11036
rect 14553 11033 14565 11036
rect 14599 11033 14611 11067
rect 14553 11027 14611 11033
rect 16761 11067 16819 11073
rect 16761 11033 16773 11067
rect 16807 11064 16819 11067
rect 18340 11064 18368 11104
rect 19058 11092 19064 11104
rect 19116 11092 19122 11144
rect 20162 11092 20168 11144
rect 20220 11132 20226 11144
rect 20438 11132 20444 11144
rect 20220 11104 20444 11132
rect 20220 11092 20226 11104
rect 20438 11092 20444 11104
rect 20496 11092 20502 11144
rect 20622 11132 20628 11144
rect 20583 11104 20628 11132
rect 20622 11092 20628 11104
rect 20680 11092 20686 11144
rect 20824 11132 20852 11308
rect 21174 11296 21180 11348
rect 21232 11336 21238 11348
rect 23106 11336 23112 11348
rect 21232 11308 23112 11336
rect 21232 11296 21238 11308
rect 23106 11296 23112 11308
rect 23164 11296 23170 11348
rect 23290 11336 23296 11348
rect 23251 11308 23296 11336
rect 23290 11296 23296 11308
rect 23348 11296 23354 11348
rect 20990 11160 20996 11212
rect 21048 11200 21054 11212
rect 21818 11200 21824 11212
rect 21048 11172 21824 11200
rect 21048 11160 21054 11172
rect 21818 11160 21824 11172
rect 21876 11160 21882 11212
rect 37366 11160 37372 11212
rect 37424 11200 37430 11212
rect 37737 11203 37795 11209
rect 37737 11200 37749 11203
rect 37424 11172 37749 11200
rect 37424 11160 37430 11172
rect 37737 11169 37749 11172
rect 37783 11169 37795 11203
rect 37737 11163 37795 11169
rect 21269 11135 21327 11141
rect 21269 11132 21281 11135
rect 20824 11104 21281 11132
rect 21269 11101 21281 11104
rect 21315 11101 21327 11135
rect 21910 11132 21916 11144
rect 21871 11104 21916 11132
rect 21269 11095 21327 11101
rect 21910 11092 21916 11104
rect 21968 11132 21974 11144
rect 22557 11135 22615 11141
rect 22557 11132 22569 11135
rect 21968 11104 22569 11132
rect 21968 11092 21974 11104
rect 22557 11101 22569 11104
rect 22603 11132 22615 11135
rect 22830 11132 22836 11144
rect 22603 11104 22836 11132
rect 22603 11101 22615 11104
rect 22557 11095 22615 11101
rect 22830 11092 22836 11104
rect 22888 11092 22894 11144
rect 23198 11132 23204 11144
rect 23159 11104 23204 11132
rect 23198 11092 23204 11104
rect 23256 11092 23262 11144
rect 26053 11135 26111 11141
rect 26053 11101 26065 11135
rect 26099 11132 26111 11135
rect 26234 11132 26240 11144
rect 26099 11104 26240 11132
rect 26099 11101 26111 11104
rect 26053 11095 26111 11101
rect 26234 11092 26240 11104
rect 26292 11092 26298 11144
rect 37182 11092 37188 11144
rect 37240 11132 37246 11144
rect 37461 11135 37519 11141
rect 37461 11132 37473 11135
rect 37240 11104 37473 11132
rect 37240 11092 37246 11104
rect 37461 11101 37473 11104
rect 37507 11101 37519 11135
rect 37461 11095 37519 11101
rect 16807 11036 18368 11064
rect 18417 11067 18475 11073
rect 16807 11033 16819 11036
rect 16761 11027 16819 11033
rect 18417 11033 18429 11067
rect 18463 11064 18475 11067
rect 18690 11064 18696 11076
rect 18463 11036 18696 11064
rect 18463 11033 18475 11036
rect 18417 11027 18475 11033
rect 18690 11024 18696 11036
rect 18748 11024 18754 11076
rect 19521 11067 19579 11073
rect 19521 11033 19533 11067
rect 19567 11033 19579 11067
rect 19521 11027 19579 11033
rect 11422 10996 11428 11008
rect 9876 10968 11428 10996
rect 11422 10956 11428 10968
rect 11480 10956 11486 11008
rect 11606 10956 11612 11008
rect 11664 10996 11670 11008
rect 12434 10996 12440 11008
rect 11664 10968 12440 10996
rect 11664 10956 11670 10968
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 12894 10956 12900 11008
rect 12952 10996 12958 11008
rect 13998 10996 14004 11008
rect 12952 10968 14004 10996
rect 12952 10956 12958 10968
rect 13998 10956 14004 10968
rect 14056 10956 14062 11008
rect 17034 10956 17040 11008
rect 17092 10996 17098 11008
rect 18506 10996 18512 11008
rect 17092 10968 18512 10996
rect 17092 10956 17098 10968
rect 18506 10956 18512 10968
rect 18564 10956 18570 11008
rect 18874 10956 18880 11008
rect 18932 10996 18938 11008
rect 19536 10996 19564 11027
rect 19610 11024 19616 11076
rect 19668 11064 19674 11076
rect 19668 11036 19713 11064
rect 19668 11024 19674 11036
rect 20254 11024 20260 11076
rect 20312 11064 20318 11076
rect 22005 11067 22063 11073
rect 22005 11064 22017 11067
rect 20312 11036 22017 11064
rect 20312 11024 20318 11036
rect 22005 11033 22017 11036
rect 22051 11033 22063 11067
rect 26142 11064 26148 11076
rect 26103 11036 26148 11064
rect 22005 11027 22063 11033
rect 26142 11024 26148 11036
rect 26200 11024 26206 11076
rect 20622 10996 20628 11008
rect 18932 10968 20628 10996
rect 18932 10956 18938 10968
rect 20622 10956 20628 10968
rect 20680 10956 20686 11008
rect 20717 10999 20775 11005
rect 20717 10965 20729 10999
rect 20763 10996 20775 10999
rect 20898 10996 20904 11008
rect 20763 10968 20904 10996
rect 20763 10965 20775 10968
rect 20717 10959 20775 10965
rect 20898 10956 20904 10968
rect 20956 10956 20962 11008
rect 21358 10996 21364 11008
rect 21319 10968 21364 10996
rect 21358 10956 21364 10968
rect 21416 10956 21422 11008
rect 22646 10996 22652 11008
rect 22607 10968 22652 10996
rect 22646 10956 22652 10968
rect 22704 10956 22710 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 1762 10752 1768 10804
rect 1820 10792 1826 10804
rect 1949 10795 2007 10801
rect 1949 10792 1961 10795
rect 1820 10764 1961 10792
rect 1820 10752 1826 10764
rect 1949 10761 1961 10764
rect 1995 10761 2007 10795
rect 2590 10792 2596 10804
rect 2551 10764 2596 10792
rect 1949 10755 2007 10761
rect 2590 10752 2596 10764
rect 2648 10752 2654 10804
rect 3050 10752 3056 10804
rect 3108 10792 3114 10804
rect 3237 10795 3295 10801
rect 3237 10792 3249 10795
rect 3108 10764 3249 10792
rect 3108 10752 3114 10764
rect 3237 10761 3249 10764
rect 3283 10761 3295 10795
rect 5534 10792 5540 10804
rect 5495 10764 5540 10792
rect 3237 10755 3295 10761
rect 5534 10752 5540 10764
rect 5592 10752 5598 10804
rect 9766 10792 9772 10804
rect 6748 10764 9772 10792
rect 3602 10724 3608 10736
rect 2516 10696 3608 10724
rect 2516 10665 2544 10696
rect 3602 10684 3608 10696
rect 3660 10684 3666 10736
rect 5442 10724 5448 10736
rect 5290 10696 5448 10724
rect 5442 10684 5448 10696
rect 5500 10684 5506 10736
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10625 1915 10659
rect 1857 10619 1915 10625
rect 2501 10659 2559 10665
rect 2501 10625 2513 10659
rect 2547 10625 2559 10659
rect 2501 10619 2559 10625
rect 1872 10588 1900 10619
rect 2590 10616 2596 10668
rect 2648 10656 2654 10668
rect 3145 10659 3203 10665
rect 3145 10656 3157 10659
rect 2648 10628 3157 10656
rect 2648 10616 2654 10628
rect 3145 10625 3157 10628
rect 3191 10625 3203 10659
rect 3786 10656 3792 10668
rect 3747 10628 3792 10656
rect 3145 10619 3203 10625
rect 3786 10616 3792 10628
rect 3844 10616 3850 10668
rect 6748 10665 6776 10764
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 11793 10795 11851 10801
rect 11793 10761 11805 10795
rect 11839 10792 11851 10795
rect 12250 10792 12256 10804
rect 11839 10764 12256 10792
rect 11839 10761 11851 10764
rect 11793 10755 11851 10761
rect 12250 10752 12256 10764
rect 12308 10752 12314 10804
rect 12437 10795 12495 10801
rect 12437 10761 12449 10795
rect 12483 10792 12495 10795
rect 12526 10792 12532 10804
rect 12483 10764 12532 10792
rect 12483 10761 12495 10764
rect 12437 10755 12495 10761
rect 12526 10752 12532 10764
rect 12584 10752 12590 10804
rect 17497 10795 17555 10801
rect 12912 10764 17080 10792
rect 6914 10684 6920 10736
rect 6972 10724 6978 10736
rect 7282 10724 7288 10736
rect 6972 10696 7288 10724
rect 6972 10684 6978 10696
rect 7282 10684 7288 10696
rect 7340 10684 7346 10736
rect 9490 10724 9496 10736
rect 8234 10696 9496 10724
rect 9490 10684 9496 10696
rect 9548 10684 9554 10736
rect 9582 10684 9588 10736
rect 9640 10724 9646 10736
rect 10594 10724 10600 10736
rect 9640 10696 10600 10724
rect 9640 10684 9646 10696
rect 10594 10684 10600 10696
rect 10652 10684 10658 10736
rect 10689 10727 10747 10733
rect 10689 10693 10701 10727
rect 10735 10724 10747 10727
rect 11054 10724 11060 10736
rect 10735 10696 11060 10724
rect 10735 10693 10747 10696
rect 10689 10687 10747 10693
rect 11054 10684 11060 10696
rect 11112 10684 11118 10736
rect 12066 10684 12072 10736
rect 12124 10724 12130 10736
rect 12710 10724 12716 10736
rect 12124 10696 12716 10724
rect 12124 10684 12130 10696
rect 12710 10684 12716 10696
rect 12768 10684 12774 10736
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10625 6791 10659
rect 6733 10619 6791 10625
rect 8294 10616 8300 10668
rect 8352 10656 8358 10668
rect 8941 10659 8999 10665
rect 8941 10656 8953 10659
rect 8352 10628 8953 10656
rect 8352 10616 8358 10628
rect 8941 10625 8953 10628
rect 8987 10625 8999 10659
rect 8941 10619 8999 10625
rect 11330 10616 11336 10668
rect 11388 10656 11394 10668
rect 11693 10657 11751 10663
rect 11388 10654 11652 10656
rect 11693 10654 11705 10657
rect 11388 10628 11705 10654
rect 11388 10616 11394 10628
rect 11624 10626 11705 10628
rect 11693 10623 11705 10626
rect 11739 10623 11751 10657
rect 11693 10617 11751 10623
rect 11882 10616 11888 10668
rect 11940 10656 11946 10668
rect 12345 10659 12403 10665
rect 12345 10656 12357 10659
rect 11940 10628 12357 10656
rect 11940 10616 11946 10628
rect 12345 10625 12357 10628
rect 12391 10625 12403 10659
rect 12345 10619 12403 10625
rect 3694 10588 3700 10600
rect 1872 10560 3700 10588
rect 3694 10548 3700 10560
rect 3752 10548 3758 10600
rect 4065 10591 4123 10597
rect 4065 10557 4077 10591
rect 4111 10588 4123 10591
rect 5258 10588 5264 10600
rect 4111 10560 5264 10588
rect 4111 10557 4123 10560
rect 4065 10551 4123 10557
rect 5258 10548 5264 10560
rect 5316 10548 5322 10600
rect 7009 10591 7067 10597
rect 7009 10557 7021 10591
rect 7055 10588 7067 10591
rect 10686 10588 10692 10600
rect 7055 10560 10692 10588
rect 7055 10557 7067 10560
rect 7009 10551 7067 10557
rect 10686 10548 10692 10560
rect 10744 10548 10750 10600
rect 9122 10520 9128 10532
rect 8496 10492 9128 10520
rect 5810 10412 5816 10464
rect 5868 10452 5874 10464
rect 8294 10452 8300 10464
rect 5868 10424 8300 10452
rect 5868 10412 5874 10424
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 8496 10461 8524 10492
rect 9122 10480 9128 10492
rect 9180 10520 9186 10532
rect 12618 10520 12624 10532
rect 9180 10492 12624 10520
rect 9180 10480 9186 10492
rect 12618 10480 12624 10492
rect 12676 10480 12682 10532
rect 8481 10455 8539 10461
rect 8481 10421 8493 10455
rect 8527 10421 8539 10455
rect 8481 10415 8539 10421
rect 11882 10412 11888 10464
rect 11940 10452 11946 10464
rect 12912 10452 12940 10764
rect 13170 10684 13176 10736
rect 13228 10724 13234 10736
rect 13265 10727 13323 10733
rect 13265 10724 13277 10727
rect 13228 10696 13277 10724
rect 13228 10684 13234 10696
rect 13265 10693 13277 10696
rect 13311 10693 13323 10727
rect 13265 10687 13323 10693
rect 15654 10684 15660 10736
rect 15712 10724 15718 10736
rect 15749 10727 15807 10733
rect 15749 10724 15761 10727
rect 15712 10696 15761 10724
rect 15712 10684 15718 10696
rect 15749 10693 15761 10696
rect 15795 10693 15807 10727
rect 15749 10687 15807 10693
rect 14366 10616 14372 10668
rect 14424 10616 14430 10668
rect 16942 10656 16948 10668
rect 16776 10628 16948 10656
rect 12989 10591 13047 10597
rect 12989 10557 13001 10591
rect 13035 10557 13047 10591
rect 12989 10551 13047 10557
rect 11940 10424 12940 10452
rect 13004 10452 13032 10551
rect 13722 10548 13728 10600
rect 13780 10588 13786 10600
rect 15010 10588 15016 10600
rect 13780 10560 14320 10588
rect 14971 10560 15016 10588
rect 13780 10548 13786 10560
rect 14292 10520 14320 10560
rect 15010 10548 15016 10560
rect 15068 10548 15074 10600
rect 15657 10591 15715 10597
rect 15657 10557 15669 10591
rect 15703 10588 15715 10591
rect 16776 10588 16804 10628
rect 16942 10616 16948 10628
rect 17000 10616 17006 10668
rect 17052 10665 17080 10764
rect 17497 10761 17509 10795
rect 17543 10792 17555 10795
rect 17954 10792 17960 10804
rect 17543 10764 17960 10792
rect 17543 10761 17555 10764
rect 17497 10755 17555 10761
rect 17954 10752 17960 10764
rect 18012 10752 18018 10804
rect 21358 10792 21364 10804
rect 18156 10764 21364 10792
rect 18156 10733 18184 10764
rect 21358 10752 21364 10764
rect 21416 10752 21422 10804
rect 23750 10792 23756 10804
rect 22664 10764 23756 10792
rect 18141 10727 18199 10733
rect 18141 10693 18153 10727
rect 18187 10693 18199 10727
rect 18141 10687 18199 10693
rect 18414 10684 18420 10736
rect 18472 10724 18478 10736
rect 19705 10727 19763 10733
rect 19705 10724 19717 10727
rect 18472 10696 19717 10724
rect 18472 10684 18478 10696
rect 19705 10693 19717 10696
rect 19751 10693 19763 10727
rect 20898 10724 20904 10736
rect 20859 10696 20904 10724
rect 19705 10687 19763 10693
rect 20898 10684 20904 10696
rect 20956 10684 20962 10736
rect 21174 10684 21180 10736
rect 21232 10724 21238 10736
rect 22664 10724 22692 10764
rect 23750 10752 23756 10764
rect 23808 10752 23814 10804
rect 23566 10724 23572 10736
rect 21232 10696 22692 10724
rect 21232 10684 21238 10696
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10625 17095 10659
rect 17037 10619 17095 10625
rect 22005 10659 22063 10665
rect 22005 10625 22017 10659
rect 22051 10656 22063 10659
rect 22186 10656 22192 10668
rect 22051 10628 22192 10656
rect 22051 10625 22063 10628
rect 22005 10619 22063 10625
rect 22186 10616 22192 10628
rect 22244 10616 22250 10668
rect 22664 10665 22692 10696
rect 23492 10696 23572 10724
rect 23492 10665 23520 10696
rect 23566 10684 23572 10696
rect 23624 10684 23630 10736
rect 22649 10659 22707 10665
rect 22649 10625 22661 10659
rect 22695 10625 22707 10659
rect 22649 10619 22707 10625
rect 23477 10659 23535 10665
rect 23477 10625 23489 10659
rect 23523 10625 23535 10659
rect 24670 10656 24676 10668
rect 24631 10628 24676 10656
rect 23477 10619 23535 10625
rect 24670 10616 24676 10628
rect 24728 10616 24734 10668
rect 15703 10560 16804 10588
rect 16853 10591 16911 10597
rect 15703 10557 15715 10560
rect 15657 10551 15715 10557
rect 16853 10557 16865 10591
rect 16899 10557 16911 10591
rect 16853 10551 16911 10557
rect 18049 10591 18107 10597
rect 18049 10557 18061 10591
rect 18095 10588 18107 10591
rect 18322 10588 18328 10600
rect 18095 10560 18328 10588
rect 18095 10557 18107 10560
rect 18049 10551 18107 10557
rect 15562 10520 15568 10532
rect 14292 10492 15568 10520
rect 15562 10480 15568 10492
rect 15620 10480 15626 10532
rect 16209 10523 16267 10529
rect 16209 10489 16221 10523
rect 16255 10489 16267 10523
rect 16868 10520 16896 10551
rect 18322 10548 18328 10560
rect 18380 10548 18386 10600
rect 19061 10591 19119 10597
rect 19061 10557 19073 10591
rect 19107 10588 19119 10591
rect 19150 10588 19156 10600
rect 19107 10560 19156 10588
rect 19107 10557 19119 10560
rect 19061 10551 19119 10557
rect 19150 10548 19156 10560
rect 19208 10548 19214 10600
rect 19613 10591 19671 10597
rect 19613 10557 19625 10591
rect 19659 10588 19671 10591
rect 20809 10591 20867 10597
rect 19659 10560 20300 10588
rect 19659 10557 19671 10560
rect 19613 10551 19671 10557
rect 19628 10520 19656 10551
rect 20162 10520 20168 10532
rect 16868 10492 19656 10520
rect 20123 10492 20168 10520
rect 16209 10483 16267 10489
rect 13814 10452 13820 10464
rect 13004 10424 13820 10452
rect 11940 10412 11946 10424
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 16224 10452 16252 10483
rect 20162 10480 20168 10492
rect 20220 10480 20226 10532
rect 20272 10520 20300 10560
rect 20809 10557 20821 10591
rect 20855 10588 20867 10591
rect 20855 10560 21496 10588
rect 20855 10557 20867 10560
rect 20809 10551 20867 10557
rect 20990 10520 20996 10532
rect 20272 10492 20996 10520
rect 20990 10480 20996 10492
rect 21048 10480 21054 10532
rect 21082 10480 21088 10532
rect 21140 10520 21146 10532
rect 21358 10520 21364 10532
rect 21140 10492 21364 10520
rect 21140 10480 21146 10492
rect 21358 10480 21364 10492
rect 21416 10480 21422 10532
rect 21468 10520 21496 10560
rect 21726 10548 21732 10600
rect 21784 10588 21790 10600
rect 23569 10591 23627 10597
rect 23569 10588 23581 10591
rect 21784 10560 23581 10588
rect 21784 10548 21790 10560
rect 23569 10557 23581 10560
rect 23615 10557 23627 10591
rect 23569 10551 23627 10557
rect 22738 10520 22744 10532
rect 21468 10492 22600 10520
rect 22699 10492 22744 10520
rect 16758 10452 16764 10464
rect 16224 10424 16764 10452
rect 16758 10412 16764 10424
rect 16816 10452 16822 10464
rect 17218 10452 17224 10464
rect 16816 10424 17224 10452
rect 16816 10412 16822 10424
rect 17218 10412 17224 10424
rect 17276 10412 17282 10464
rect 19058 10412 19064 10464
rect 19116 10452 19122 10464
rect 22097 10455 22155 10461
rect 22097 10452 22109 10455
rect 19116 10424 22109 10452
rect 19116 10412 19122 10424
rect 22097 10421 22109 10424
rect 22143 10421 22155 10455
rect 22572 10452 22600 10492
rect 22738 10480 22744 10492
rect 22796 10480 22802 10532
rect 23658 10452 23664 10464
rect 22572 10424 23664 10452
rect 22097 10415 22155 10421
rect 23658 10412 23664 10424
rect 23716 10412 23722 10464
rect 24489 10455 24547 10461
rect 24489 10421 24501 10455
rect 24535 10452 24547 10455
rect 26050 10452 26056 10464
rect 24535 10424 26056 10452
rect 24535 10421 24547 10424
rect 24489 10415 24547 10421
rect 26050 10412 26056 10424
rect 26108 10412 26114 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 2590 10248 2596 10260
rect 2551 10220 2596 10248
rect 2590 10208 2596 10220
rect 2648 10208 2654 10260
rect 3329 10251 3387 10257
rect 3329 10217 3341 10251
rect 3375 10248 3387 10251
rect 4706 10248 4712 10260
rect 3375 10220 4712 10248
rect 3375 10217 3387 10220
rect 3329 10211 3387 10217
rect 4706 10208 4712 10220
rect 4764 10208 4770 10260
rect 5721 10251 5779 10257
rect 5721 10217 5733 10251
rect 5767 10248 5779 10251
rect 6914 10248 6920 10260
rect 5767 10220 6920 10248
rect 5767 10217 5779 10220
rect 5721 10211 5779 10217
rect 6914 10208 6920 10220
rect 6972 10208 6978 10260
rect 9674 10208 9680 10260
rect 9732 10248 9738 10260
rect 10321 10251 10379 10257
rect 9732 10220 9777 10248
rect 9732 10208 9738 10220
rect 10321 10217 10333 10251
rect 10367 10248 10379 10251
rect 11882 10248 11888 10260
rect 10367 10220 11888 10248
rect 10367 10217 10379 10220
rect 10321 10211 10379 10217
rect 11882 10208 11888 10220
rect 11940 10208 11946 10260
rect 12158 10208 12164 10260
rect 12216 10248 12222 10260
rect 12216 10220 12756 10248
rect 12216 10208 12222 10220
rect 2041 10183 2099 10189
rect 2041 10149 2053 10183
rect 2087 10180 2099 10183
rect 2866 10180 2872 10192
rect 2087 10152 2872 10180
rect 2087 10149 2099 10152
rect 2041 10143 2099 10149
rect 2866 10140 2872 10152
rect 2924 10140 2930 10192
rect 6086 10180 6092 10192
rect 5276 10152 6092 10180
rect 4249 10115 4307 10121
rect 1964 10084 3832 10112
rect 566 10004 572 10056
rect 624 10044 630 10056
rect 1964 10053 1992 10084
rect 1949 10047 2007 10053
rect 1949 10044 1961 10047
rect 624 10016 1961 10044
rect 624 10004 630 10016
rect 1949 10013 1961 10016
rect 1995 10013 2007 10047
rect 1949 10007 2007 10013
rect 2777 10047 2835 10053
rect 2777 10013 2789 10047
rect 2823 10044 2835 10047
rect 3142 10044 3148 10056
rect 2823 10016 3148 10044
rect 2823 10013 2835 10016
rect 2777 10007 2835 10013
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10044 3295 10047
rect 3694 10044 3700 10056
rect 3283 10016 3700 10044
rect 3283 10013 3295 10016
rect 3237 10007 3295 10013
rect 3694 10004 3700 10016
rect 3752 10004 3758 10056
rect 3804 9976 3832 10084
rect 4249 10081 4261 10115
rect 4295 10112 4307 10115
rect 5276 10112 5304 10152
rect 6086 10140 6092 10152
rect 6144 10140 6150 10192
rect 12728 10180 12756 10220
rect 14366 10208 14372 10260
rect 14424 10248 14430 10260
rect 22646 10248 22652 10260
rect 14424 10220 22652 10248
rect 14424 10208 14430 10220
rect 22646 10208 22652 10220
rect 22704 10208 22710 10260
rect 14182 10180 14188 10192
rect 12728 10152 14188 10180
rect 14182 10140 14188 10152
rect 14240 10140 14246 10192
rect 15562 10140 15568 10192
rect 15620 10180 15626 10192
rect 18966 10180 18972 10192
rect 15620 10152 18972 10180
rect 15620 10140 15626 10152
rect 18966 10140 18972 10152
rect 19024 10140 19030 10192
rect 19150 10140 19156 10192
rect 19208 10180 19214 10192
rect 21450 10180 21456 10192
rect 19208 10152 21456 10180
rect 19208 10140 19214 10152
rect 8570 10112 8576 10124
rect 4295 10084 5304 10112
rect 5368 10084 8576 10112
rect 4295 10081 4307 10084
rect 4249 10075 4307 10081
rect 3970 10044 3976 10056
rect 3931 10016 3976 10044
rect 3970 10004 3976 10016
rect 4028 10004 4034 10056
rect 5368 10030 5396 10084
rect 8570 10072 8576 10084
rect 8628 10072 8634 10124
rect 10873 10115 10931 10121
rect 10873 10081 10885 10115
rect 10919 10112 10931 10115
rect 12452 10112 12572 10124
rect 13814 10112 13820 10124
rect 10919 10096 13820 10112
rect 10919 10084 12480 10096
rect 12544 10084 13820 10096
rect 10919 10081 10931 10084
rect 10873 10075 10931 10081
rect 13814 10072 13820 10084
rect 13872 10112 13878 10124
rect 14274 10112 14280 10124
rect 13872 10084 14280 10112
rect 13872 10072 13878 10084
rect 14274 10072 14280 10084
rect 14332 10112 14338 10124
rect 17313 10115 17371 10121
rect 17313 10112 17325 10115
rect 14332 10084 17325 10112
rect 14332 10072 14338 10084
rect 17313 10081 17325 10084
rect 17359 10081 17371 10115
rect 17313 10075 17371 10081
rect 17586 10072 17592 10124
rect 17644 10112 17650 10124
rect 19521 10115 19579 10121
rect 19521 10112 19533 10115
rect 17644 10084 19533 10112
rect 17644 10072 17650 10084
rect 19521 10081 19533 10084
rect 19567 10112 19579 10115
rect 20070 10112 20076 10124
rect 19567 10084 20076 10112
rect 19567 10081 19579 10084
rect 19521 10075 19579 10081
rect 20070 10072 20076 10084
rect 20128 10072 20134 10124
rect 20548 10121 20576 10152
rect 21450 10140 21456 10152
rect 21508 10140 21514 10192
rect 21542 10140 21548 10192
rect 21600 10180 21606 10192
rect 21637 10183 21695 10189
rect 21637 10180 21649 10183
rect 21600 10152 21649 10180
rect 21600 10140 21606 10152
rect 21637 10149 21649 10152
rect 21683 10149 21695 10183
rect 29825 10183 29883 10189
rect 29825 10180 29837 10183
rect 21637 10143 21695 10149
rect 22066 10152 29837 10180
rect 20533 10115 20591 10121
rect 20533 10081 20545 10115
rect 20579 10081 20591 10115
rect 20533 10075 20591 10081
rect 20622 10072 20628 10124
rect 20680 10112 20686 10124
rect 22066 10112 22094 10152
rect 29825 10149 29837 10152
rect 29871 10149 29883 10183
rect 29825 10143 29883 10149
rect 20680 10084 22094 10112
rect 22465 10115 22523 10121
rect 20680 10072 20686 10084
rect 22465 10081 22477 10115
rect 22511 10112 22523 10115
rect 23477 10115 23535 10121
rect 23477 10112 23489 10115
rect 22511 10084 23489 10112
rect 22511 10081 22523 10084
rect 22465 10075 22523 10081
rect 23477 10081 23489 10084
rect 23523 10081 23535 10115
rect 23477 10075 23535 10081
rect 6457 10047 6515 10053
rect 6457 10013 6469 10047
rect 6503 10013 6515 10047
rect 6457 10007 6515 10013
rect 9585 10047 9643 10053
rect 9585 10013 9597 10047
rect 9631 10044 9643 10047
rect 9858 10044 9864 10056
rect 9631 10016 9864 10044
rect 9631 10013 9643 10016
rect 9585 10007 9643 10013
rect 4522 9976 4528 9988
rect 3804 9948 4528 9976
rect 4522 9936 4528 9948
rect 4580 9936 4586 9988
rect 6472 9976 6500 10007
rect 9858 10004 9864 10016
rect 9916 10004 9922 10056
rect 10229 10047 10287 10053
rect 10229 10013 10241 10047
rect 10275 10044 10287 10047
rect 10778 10044 10784 10056
rect 10275 10016 10784 10044
rect 10275 10013 10287 10016
rect 10229 10007 10287 10013
rect 6472 9948 6592 9976
rect 4154 9868 4160 9920
rect 4212 9908 4218 9920
rect 6178 9908 6184 9920
rect 4212 9880 6184 9908
rect 4212 9868 4218 9880
rect 6178 9868 6184 9880
rect 6236 9868 6242 9920
rect 6564 9908 6592 9948
rect 6638 9936 6644 9988
rect 6696 9976 6702 9988
rect 6733 9979 6791 9985
rect 6733 9976 6745 9979
rect 6696 9948 6745 9976
rect 6696 9936 6702 9948
rect 6733 9945 6745 9948
rect 6779 9945 6791 9979
rect 6733 9939 6791 9945
rect 7190 9936 7196 9988
rect 7248 9936 7254 9988
rect 9674 9936 9680 9988
rect 9732 9976 9738 9988
rect 10244 9976 10272 10007
rect 10778 10004 10784 10016
rect 10836 10004 10842 10056
rect 12894 10044 12900 10056
rect 12855 10016 12900 10044
rect 12894 10004 12900 10016
rect 12952 10004 12958 10056
rect 13541 10047 13599 10053
rect 13541 10013 13553 10047
rect 13587 10044 13599 10047
rect 13998 10044 14004 10056
rect 13587 10016 14004 10044
rect 13587 10013 13599 10016
rect 13541 10007 13599 10013
rect 13998 10004 14004 10016
rect 14056 10004 14062 10056
rect 16577 10047 16635 10053
rect 16577 10013 16589 10047
rect 16623 10044 16635 10047
rect 16666 10044 16672 10056
rect 16623 10016 16672 10044
rect 16623 10013 16635 10016
rect 16577 10007 16635 10013
rect 16666 10004 16672 10016
rect 16724 10004 16730 10056
rect 17957 10047 18015 10053
rect 17957 10013 17969 10047
rect 18003 10044 18015 10047
rect 18046 10044 18052 10056
rect 18003 10016 18052 10044
rect 18003 10013 18015 10016
rect 17957 10007 18015 10013
rect 18046 10004 18052 10016
rect 18104 10004 18110 10056
rect 22278 10044 22284 10056
rect 18156 10016 19380 10044
rect 22239 10016 22284 10044
rect 11146 9976 11152 9988
rect 9732 9948 10272 9976
rect 11107 9948 11152 9976
rect 9732 9936 9738 9948
rect 11146 9936 11152 9948
rect 11204 9936 11210 9988
rect 12618 9976 12624 9988
rect 12374 9948 12624 9976
rect 12618 9936 12624 9948
rect 12676 9936 12682 9988
rect 14553 9979 14611 9985
rect 14553 9976 14565 9979
rect 14384 9948 14565 9976
rect 14384 9920 14412 9948
rect 14553 9945 14565 9948
rect 14599 9945 14611 9979
rect 14553 9939 14611 9945
rect 15286 9936 15292 9988
rect 15344 9936 15350 9988
rect 15838 9936 15844 9988
rect 15896 9976 15902 9988
rect 18156 9976 18184 10016
rect 15896 9948 18184 9976
rect 18233 9979 18291 9985
rect 15896 9936 15902 9948
rect 18233 9945 18245 9979
rect 18279 9976 18291 9979
rect 18414 9976 18420 9988
rect 18279 9948 18420 9976
rect 18279 9945 18291 9948
rect 18233 9939 18291 9945
rect 18414 9936 18420 9948
rect 18472 9976 18478 9988
rect 19242 9976 19248 9988
rect 18472 9948 19248 9976
rect 18472 9936 18478 9948
rect 19242 9936 19248 9948
rect 19300 9936 19306 9988
rect 19352 9976 19380 10016
rect 22278 10004 22284 10016
rect 22336 10004 22342 10056
rect 23198 10004 23204 10056
rect 23256 10044 23262 10056
rect 23385 10047 23443 10053
rect 23385 10044 23397 10047
rect 23256 10016 23397 10044
rect 23256 10004 23262 10016
rect 23385 10013 23397 10016
rect 23431 10013 23443 10047
rect 23385 10007 23443 10013
rect 29733 10047 29791 10053
rect 29733 10013 29745 10047
rect 29779 10044 29791 10047
rect 29779 10016 35894 10044
rect 29779 10013 29791 10016
rect 29733 10007 29791 10013
rect 19518 9976 19524 9988
rect 19352 9948 19524 9976
rect 19518 9936 19524 9948
rect 19576 9936 19582 9988
rect 19613 9979 19671 9985
rect 19613 9945 19625 9979
rect 19659 9976 19671 9979
rect 20346 9976 20352 9988
rect 19659 9948 20352 9976
rect 19659 9945 19671 9948
rect 19613 9939 19671 9945
rect 20346 9936 20352 9948
rect 20404 9936 20410 9988
rect 21082 9976 21088 9988
rect 21043 9948 21088 9976
rect 21082 9936 21088 9948
rect 21140 9936 21146 9988
rect 21177 9979 21235 9985
rect 21177 9945 21189 9979
rect 21223 9976 21235 9979
rect 21726 9976 21732 9988
rect 21223 9948 21732 9976
rect 21223 9945 21235 9948
rect 21177 9939 21235 9945
rect 21726 9936 21732 9948
rect 21784 9936 21790 9988
rect 21910 9936 21916 9988
rect 21968 9976 21974 9988
rect 22925 9979 22983 9985
rect 22925 9976 22937 9979
rect 21968 9948 22937 9976
rect 21968 9936 21974 9948
rect 22925 9945 22937 9948
rect 22971 9976 22983 9979
rect 23014 9976 23020 9988
rect 22971 9948 23020 9976
rect 22971 9945 22983 9948
rect 22925 9939 22983 9945
rect 23014 9936 23020 9948
rect 23072 9936 23078 9988
rect 35866 9976 35894 10016
rect 36906 10004 36912 10056
rect 36964 10044 36970 10056
rect 38013 10047 38071 10053
rect 38013 10044 38025 10047
rect 36964 10016 38025 10044
rect 36964 10004 36970 10016
rect 38013 10013 38025 10016
rect 38059 10013 38071 10047
rect 38013 10007 38071 10013
rect 37734 9976 37740 9988
rect 35866 9948 37740 9976
rect 37734 9936 37740 9948
rect 37792 9936 37798 9988
rect 6914 9908 6920 9920
rect 6564 9880 6920 9908
rect 6914 9868 6920 9880
rect 6972 9868 6978 9920
rect 7466 9868 7472 9920
rect 7524 9908 7530 9920
rect 7650 9908 7656 9920
rect 7524 9880 7656 9908
rect 7524 9868 7530 9880
rect 7650 9868 7656 9880
rect 7708 9868 7714 9920
rect 8110 9868 8116 9920
rect 8168 9908 8174 9920
rect 8205 9911 8263 9917
rect 8205 9908 8217 9911
rect 8168 9880 8217 9908
rect 8168 9868 8174 9880
rect 8205 9877 8217 9880
rect 8251 9877 8263 9911
rect 8205 9871 8263 9877
rect 13633 9911 13691 9917
rect 13633 9877 13645 9911
rect 13679 9908 13691 9911
rect 13722 9908 13728 9920
rect 13679 9880 13728 9908
rect 13679 9877 13691 9880
rect 13633 9871 13691 9877
rect 13722 9868 13728 9880
rect 13780 9868 13786 9920
rect 14366 9868 14372 9920
rect 14424 9868 14430 9920
rect 14458 9868 14464 9920
rect 14516 9908 14522 9920
rect 16025 9911 16083 9917
rect 16025 9908 16037 9911
rect 14516 9880 16037 9908
rect 14516 9868 14522 9880
rect 16025 9877 16037 9880
rect 16071 9877 16083 9911
rect 16025 9871 16083 9877
rect 17218 9868 17224 9920
rect 17276 9908 17282 9920
rect 22002 9908 22008 9920
rect 17276 9880 22008 9908
rect 17276 9868 17282 9880
rect 22002 9868 22008 9880
rect 22060 9868 22066 9920
rect 24946 9868 24952 9920
rect 25004 9908 25010 9920
rect 25041 9911 25099 9917
rect 25041 9908 25053 9911
rect 25004 9880 25053 9908
rect 25004 9868 25010 9880
rect 25041 9877 25053 9880
rect 25087 9877 25099 9911
rect 38194 9908 38200 9920
rect 38155 9880 38200 9908
rect 25041 9871 25099 9877
rect 38194 9868 38200 9880
rect 38252 9868 38258 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 3786 9664 3792 9716
rect 3844 9704 3850 9716
rect 5350 9704 5356 9716
rect 3844 9676 5356 9704
rect 3844 9664 3850 9676
rect 5350 9664 5356 9676
rect 5408 9664 5414 9716
rect 5534 9664 5540 9716
rect 5592 9704 5598 9716
rect 5997 9707 6055 9713
rect 5592 9676 5856 9704
rect 5592 9664 5598 9676
rect 3878 9636 3884 9648
rect 3082 9608 3884 9636
rect 3878 9596 3884 9608
rect 3936 9596 3942 9648
rect 4982 9596 4988 9648
rect 5040 9596 5046 9648
rect 5828 9636 5856 9676
rect 5997 9673 6009 9707
rect 6043 9704 6055 9707
rect 6546 9704 6552 9716
rect 6043 9676 6552 9704
rect 6043 9673 6055 9676
rect 5997 9667 6055 9673
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 6638 9664 6644 9716
rect 6696 9704 6702 9716
rect 13354 9704 13360 9716
rect 6696 9676 13360 9704
rect 6696 9664 6702 9676
rect 13354 9664 13360 9676
rect 13412 9664 13418 9716
rect 14182 9664 14188 9716
rect 14240 9704 14246 9716
rect 17218 9704 17224 9716
rect 14240 9676 17224 9704
rect 14240 9664 14246 9676
rect 17218 9664 17224 9676
rect 17276 9664 17282 9716
rect 18325 9707 18383 9713
rect 18325 9673 18337 9707
rect 18371 9704 18383 9707
rect 21910 9704 21916 9716
rect 18371 9676 21916 9704
rect 18371 9673 18383 9676
rect 18325 9667 18383 9673
rect 21910 9664 21916 9676
rect 21968 9664 21974 9716
rect 22278 9664 22284 9716
rect 22336 9704 22342 9716
rect 22649 9707 22707 9713
rect 22649 9704 22661 9707
rect 22336 9676 22661 9704
rect 22336 9664 22342 9676
rect 22649 9673 22661 9676
rect 22695 9673 22707 9707
rect 22649 9667 22707 9673
rect 6656 9636 6684 9664
rect 5828 9608 6684 9636
rect 7098 9596 7104 9648
rect 7156 9636 7162 9648
rect 7653 9639 7711 9645
rect 7653 9636 7665 9639
rect 7156 9608 7665 9636
rect 7156 9596 7162 9608
rect 7653 9605 7665 9608
rect 7699 9605 7711 9639
rect 7653 9599 7711 9605
rect 8481 9639 8539 9645
rect 8481 9605 8493 9639
rect 8527 9636 8539 9639
rect 8570 9636 8576 9648
rect 8527 9608 8576 9636
rect 8527 9605 8539 9608
rect 8481 9599 8539 9605
rect 8570 9596 8576 9608
rect 8628 9596 8634 9648
rect 10778 9636 10784 9648
rect 10534 9608 10784 9636
rect 10778 9596 10784 9608
rect 10836 9596 10842 9648
rect 11054 9596 11060 9648
rect 11112 9636 11118 9648
rect 11698 9636 11704 9648
rect 11112 9608 11704 9636
rect 11112 9596 11118 9608
rect 11698 9596 11704 9608
rect 11756 9596 11762 9648
rect 11974 9596 11980 9648
rect 12032 9636 12038 9648
rect 12437 9639 12495 9645
rect 12437 9636 12449 9639
rect 12032 9608 12449 9636
rect 12032 9596 12038 9608
rect 12437 9605 12449 9608
rect 12483 9605 12495 9639
rect 13262 9636 13268 9648
rect 13223 9608 13268 9636
rect 12437 9599 12495 9605
rect 13262 9596 13268 9608
rect 13320 9596 13326 9648
rect 15470 9596 15476 9648
rect 15528 9636 15534 9648
rect 15838 9636 15844 9648
rect 15528 9608 15844 9636
rect 15528 9596 15534 9608
rect 15838 9596 15844 9608
rect 15896 9596 15902 9648
rect 16132 9608 16988 9636
rect 4154 9568 4160 9580
rect 3896 9540 4160 9568
rect 1578 9500 1584 9512
rect 1539 9472 1584 9500
rect 1578 9460 1584 9472
rect 1636 9460 1642 9512
rect 1857 9503 1915 9509
rect 1857 9469 1869 9503
rect 1903 9500 1915 9503
rect 3896 9500 3924 9540
rect 4154 9528 4160 9540
rect 4212 9528 4218 9580
rect 6917 9571 6975 9577
rect 6917 9537 6929 9571
rect 6963 9568 6975 9571
rect 7006 9568 7012 9580
rect 6963 9540 7012 9568
rect 6963 9537 6975 9540
rect 6917 9531 6975 9537
rect 7006 9528 7012 9540
rect 7064 9528 7070 9580
rect 8381 9571 8439 9577
rect 8381 9537 8393 9571
rect 8427 9568 8439 9571
rect 8938 9568 8944 9580
rect 8427 9540 8944 9568
rect 8427 9537 8439 9540
rect 8381 9531 8439 9537
rect 8938 9528 8944 9540
rect 8996 9528 9002 9580
rect 12250 9528 12256 9580
rect 12308 9568 12314 9580
rect 13173 9571 13231 9577
rect 13173 9568 13185 9571
rect 12308 9566 12388 9568
rect 12452 9566 13185 9568
rect 12308 9540 13185 9566
rect 12308 9528 12314 9540
rect 12360 9538 12480 9540
rect 13173 9537 13185 9540
rect 13219 9537 13231 9571
rect 13814 9568 13820 9580
rect 13775 9540 13820 9568
rect 13173 9531 13231 9537
rect 13814 9528 13820 9540
rect 13872 9528 13878 9580
rect 16022 9568 16028 9580
rect 15226 9540 16028 9568
rect 16022 9528 16028 9540
rect 16080 9528 16086 9580
rect 1903 9472 3924 9500
rect 1903 9469 1915 9472
rect 1857 9463 1915 9469
rect 3970 9460 3976 9512
rect 4028 9500 4034 9512
rect 4249 9503 4307 9509
rect 4249 9500 4261 9503
rect 4028 9472 4261 9500
rect 4028 9460 4034 9472
rect 4249 9469 4261 9472
rect 4295 9500 4307 9503
rect 4525 9503 4583 9509
rect 4295 9472 4384 9500
rect 4295 9469 4307 9472
rect 4249 9463 4307 9469
rect 3988 9432 4016 9460
rect 3252 9404 4016 9432
rect 1578 9324 1584 9376
rect 1636 9364 1642 9376
rect 3252 9364 3280 9404
rect 1636 9336 3280 9364
rect 3329 9367 3387 9373
rect 1636 9324 1642 9336
rect 3329 9333 3341 9367
rect 3375 9364 3387 9367
rect 3418 9364 3424 9376
rect 3375 9336 3424 9364
rect 3375 9333 3387 9336
rect 3329 9327 3387 9333
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 4356 9364 4384 9472
rect 4525 9469 4537 9503
rect 4571 9500 4583 9503
rect 5166 9500 5172 9512
rect 4571 9472 5172 9500
rect 4571 9469 4583 9472
rect 4525 9463 4583 9469
rect 5166 9460 5172 9472
rect 5224 9460 5230 9512
rect 8202 9460 8208 9512
rect 8260 9500 8266 9512
rect 9033 9503 9091 9509
rect 9033 9500 9045 9503
rect 8260 9472 9045 9500
rect 8260 9460 8266 9472
rect 9033 9469 9045 9472
rect 9079 9469 9091 9503
rect 9309 9503 9367 9509
rect 9309 9500 9321 9503
rect 9033 9463 9091 9469
rect 9140 9472 9321 9500
rect 8018 9392 8024 9444
rect 8076 9432 8082 9444
rect 9140 9432 9168 9472
rect 9309 9469 9321 9472
rect 9355 9469 9367 9503
rect 9309 9463 9367 9469
rect 9674 9460 9680 9512
rect 9732 9500 9738 9512
rect 9732 9472 11836 9500
rect 9732 9460 9738 9472
rect 8076 9404 9168 9432
rect 10781 9435 10839 9441
rect 8076 9392 8082 9404
rect 10781 9401 10793 9435
rect 10827 9432 10839 9435
rect 10962 9432 10968 9444
rect 10827 9404 10968 9432
rect 10827 9401 10839 9404
rect 10781 9395 10839 9401
rect 10962 9392 10968 9404
rect 11020 9392 11026 9444
rect 11808 9432 11836 9472
rect 11882 9460 11888 9512
rect 11940 9500 11946 9512
rect 14093 9503 14151 9509
rect 14093 9500 14105 9503
rect 11940 9472 14105 9500
rect 11940 9460 11946 9472
rect 14093 9469 14105 9472
rect 14139 9500 14151 9503
rect 14182 9500 14188 9512
rect 14139 9472 14188 9500
rect 14139 9469 14151 9472
rect 14093 9463 14151 9469
rect 14182 9460 14188 9472
rect 14240 9460 14246 9512
rect 14458 9460 14464 9512
rect 14516 9500 14522 9512
rect 16132 9500 16160 9608
rect 16298 9568 16304 9580
rect 16259 9540 16304 9568
rect 16298 9528 16304 9540
rect 16356 9528 16362 9580
rect 16853 9571 16911 9577
rect 16853 9537 16865 9571
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 14516 9472 16160 9500
rect 14516 9460 14522 9472
rect 16868 9432 16896 9531
rect 16960 9500 16988 9608
rect 18138 9596 18144 9648
rect 18196 9636 18202 9648
rect 19245 9639 19303 9645
rect 19245 9636 19257 9639
rect 18196 9608 19257 9636
rect 18196 9596 18202 9608
rect 19245 9605 19257 9608
rect 19291 9605 19303 9639
rect 19245 9599 19303 9605
rect 19889 9639 19947 9645
rect 19889 9605 19901 9639
rect 19935 9636 19947 9639
rect 20530 9636 20536 9648
rect 19935 9608 20536 9636
rect 19935 9605 19947 9608
rect 19889 9599 19947 9605
rect 20530 9596 20536 9608
rect 20588 9596 20594 9648
rect 20901 9639 20959 9645
rect 20901 9605 20913 9639
rect 20947 9636 20959 9639
rect 23477 9639 23535 9645
rect 23477 9636 23489 9639
rect 20947 9608 23489 9636
rect 20947 9605 20959 9608
rect 20901 9599 20959 9605
rect 23477 9605 23489 9608
rect 23523 9605 23535 9639
rect 24946 9636 24952 9648
rect 24907 9608 24952 9636
rect 23477 9599 23535 9605
rect 24946 9596 24952 9608
rect 25004 9596 25010 9648
rect 25038 9596 25044 9648
rect 25096 9636 25102 9648
rect 25096 9608 25141 9636
rect 25096 9596 25102 9608
rect 17402 9528 17408 9580
rect 17460 9568 17466 9580
rect 17681 9571 17739 9577
rect 17681 9568 17693 9571
rect 17460 9540 17693 9568
rect 17460 9528 17466 9540
rect 17681 9537 17693 9540
rect 17727 9537 17739 9571
rect 17681 9531 17739 9537
rect 17865 9571 17923 9577
rect 17865 9537 17877 9571
rect 17911 9568 17923 9571
rect 19058 9568 19064 9580
rect 17911 9540 19064 9568
rect 17911 9537 17923 9540
rect 17865 9531 17923 9537
rect 19058 9528 19064 9540
rect 19116 9528 19122 9580
rect 19150 9528 19156 9580
rect 19208 9568 19214 9580
rect 19797 9571 19855 9577
rect 19208 9540 19253 9568
rect 19208 9528 19214 9540
rect 19797 9537 19809 9571
rect 19843 9537 19855 9571
rect 19797 9531 19855 9537
rect 19812 9500 19840 9531
rect 19978 9528 19984 9580
rect 20036 9568 20042 9580
rect 20622 9568 20628 9580
rect 20036 9540 20628 9568
rect 20036 9528 20042 9540
rect 20622 9528 20628 9540
rect 20680 9528 20686 9580
rect 21453 9571 21511 9577
rect 21453 9537 21465 9571
rect 21499 9568 21511 9571
rect 21542 9568 21548 9580
rect 21499 9540 21548 9568
rect 21499 9537 21511 9540
rect 21453 9531 21511 9537
rect 21542 9528 21548 9540
rect 21600 9528 21606 9580
rect 22002 9568 22008 9580
rect 21963 9540 22008 9568
rect 22002 9528 22008 9540
rect 22060 9528 22066 9580
rect 22094 9528 22100 9580
rect 22152 9568 22158 9580
rect 22152 9540 22197 9568
rect 22152 9528 22158 9540
rect 22278 9528 22284 9580
rect 22336 9568 22342 9580
rect 22830 9568 22836 9580
rect 22336 9540 22836 9568
rect 22336 9528 22342 9540
rect 22830 9528 22836 9540
rect 22888 9528 22894 9580
rect 23382 9568 23388 9580
rect 23343 9540 23388 9568
rect 23382 9528 23388 9540
rect 23440 9528 23446 9580
rect 23934 9528 23940 9580
rect 23992 9568 23998 9580
rect 24029 9571 24087 9577
rect 24029 9568 24041 9571
rect 23992 9540 24041 9568
rect 23992 9528 23998 9540
rect 24029 9537 24041 9540
rect 24075 9537 24087 9571
rect 24029 9531 24087 9537
rect 29917 9571 29975 9577
rect 29917 9537 29929 9571
rect 29963 9568 29975 9571
rect 31386 9568 31392 9580
rect 29963 9540 31392 9568
rect 29963 9537 29975 9540
rect 29917 9531 29975 9537
rect 31386 9528 31392 9540
rect 31444 9528 31450 9580
rect 16960 9472 19840 9500
rect 20809 9503 20867 9509
rect 20809 9469 20821 9503
rect 20855 9500 20867 9503
rect 20990 9500 20996 9512
rect 20855 9472 20996 9500
rect 20855 9469 20867 9472
rect 20809 9463 20867 9469
rect 20990 9460 20996 9472
rect 21048 9460 21054 9512
rect 21082 9460 21088 9512
rect 21140 9500 21146 9512
rect 25225 9503 25283 9509
rect 25225 9500 25237 9503
rect 21140 9472 25237 9500
rect 21140 9460 21146 9472
rect 24872 9444 24900 9472
rect 25225 9469 25237 9472
rect 25271 9469 25283 9503
rect 25225 9463 25283 9469
rect 18046 9432 18052 9444
rect 11808 9404 13952 9432
rect 4706 9364 4712 9376
rect 4356 9336 4712 9364
rect 4706 9324 4712 9336
rect 4764 9324 4770 9376
rect 8110 9324 8116 9376
rect 8168 9364 8174 9376
rect 12250 9364 12256 9376
rect 8168 9336 12256 9364
rect 8168 9324 8174 9336
rect 12250 9324 12256 9336
rect 12308 9324 12314 9376
rect 13924 9364 13952 9404
rect 15488 9404 18052 9432
rect 15488 9364 15516 9404
rect 18046 9392 18052 9404
rect 18104 9392 18110 9444
rect 18598 9392 18604 9444
rect 18656 9432 18662 9444
rect 21726 9432 21732 9444
rect 18656 9404 21732 9432
rect 18656 9392 18662 9404
rect 21726 9392 21732 9404
rect 21784 9392 21790 9444
rect 22002 9392 22008 9444
rect 22060 9432 22066 9444
rect 24026 9432 24032 9444
rect 22060 9404 24032 9432
rect 22060 9392 22094 9404
rect 24026 9392 24032 9404
rect 24084 9392 24090 9444
rect 24854 9392 24860 9444
rect 24912 9392 24918 9444
rect 13924 9336 15516 9364
rect 15562 9324 15568 9376
rect 15620 9364 15626 9376
rect 16117 9367 16175 9373
rect 15620 9336 15665 9364
rect 15620 9324 15626 9336
rect 16117 9333 16129 9367
rect 16163 9364 16175 9367
rect 16942 9364 16948 9376
rect 16163 9336 16948 9364
rect 16163 9333 16175 9336
rect 16117 9327 16175 9333
rect 16942 9324 16948 9336
rect 17000 9324 17006 9376
rect 17037 9367 17095 9373
rect 17037 9333 17049 9367
rect 17083 9364 17095 9367
rect 19334 9364 19340 9376
rect 17083 9336 19340 9364
rect 17083 9333 17095 9336
rect 17037 9327 17095 9333
rect 19334 9324 19340 9336
rect 19392 9364 19398 9376
rect 20070 9364 20076 9376
rect 19392 9336 20076 9364
rect 19392 9324 19398 9336
rect 20070 9324 20076 9336
rect 20128 9324 20134 9376
rect 20162 9324 20168 9376
rect 20220 9364 20226 9376
rect 22066 9364 22094 9392
rect 20220 9336 22094 9364
rect 20220 9324 20226 9336
rect 22186 9324 22192 9376
rect 22244 9364 22250 9376
rect 24121 9367 24179 9373
rect 24121 9364 24133 9367
rect 22244 9336 24133 9364
rect 22244 9324 22250 9336
rect 24121 9333 24133 9336
rect 24167 9333 24179 9367
rect 30006 9364 30012 9376
rect 29967 9336 30012 9364
rect 24121 9327 24179 9333
rect 30006 9324 30012 9336
rect 30064 9324 30070 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 2038 9160 2044 9172
rect 1999 9132 2044 9160
rect 2038 9120 2044 9132
rect 2096 9120 2102 9172
rect 2498 9120 2504 9172
rect 2556 9160 2562 9172
rect 2593 9163 2651 9169
rect 2593 9160 2605 9163
rect 2556 9132 2605 9160
rect 2556 9120 2562 9132
rect 2593 9129 2605 9132
rect 2639 9129 2651 9163
rect 3326 9160 3332 9172
rect 3287 9132 3332 9160
rect 2593 9123 2651 9129
rect 3326 9120 3332 9132
rect 3384 9120 3390 9172
rect 6641 9163 6699 9169
rect 6641 9129 6653 9163
rect 6687 9160 6699 9163
rect 7742 9160 7748 9172
rect 6687 9132 7748 9160
rect 6687 9129 6699 9132
rect 6641 9123 6699 9129
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 8938 9120 8944 9172
rect 8996 9160 9002 9172
rect 9858 9160 9864 9172
rect 8996 9132 9864 9160
rect 8996 9120 9002 9132
rect 9858 9120 9864 9132
rect 9916 9160 9922 9172
rect 12250 9160 12256 9172
rect 9916 9132 12256 9160
rect 9916 9120 9922 9132
rect 12250 9120 12256 9132
rect 12308 9120 12314 9172
rect 12618 9160 12624 9172
rect 12579 9132 12624 9160
rect 12618 9120 12624 9132
rect 12676 9120 12682 9172
rect 13265 9163 13323 9169
rect 13265 9129 13277 9163
rect 13311 9160 13323 9163
rect 15286 9160 15292 9172
rect 13311 9132 15292 9160
rect 13311 9129 13323 9132
rect 13265 9123 13323 9129
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 16022 9120 16028 9172
rect 16080 9160 16086 9172
rect 21542 9160 21548 9172
rect 16080 9132 21548 9160
rect 16080 9120 16086 9132
rect 21542 9120 21548 9132
rect 21600 9120 21606 9172
rect 21726 9120 21732 9172
rect 21784 9160 21790 9172
rect 23474 9160 23480 9172
rect 21784 9132 23336 9160
rect 23435 9132 23480 9160
rect 21784 9120 21790 9132
rect 5445 9095 5503 9101
rect 5445 9061 5457 9095
rect 5491 9092 5503 9095
rect 7466 9092 7472 9104
rect 5491 9064 7472 9092
rect 5491 9061 5503 9064
rect 5445 9055 5503 9061
rect 7466 9052 7472 9064
rect 7524 9052 7530 9104
rect 8386 9052 8392 9104
rect 8444 9092 8450 9104
rect 11701 9095 11759 9101
rect 11701 9092 11713 9095
rect 8444 9064 10088 9092
rect 8444 9052 8450 9064
rect 4706 9024 4712 9036
rect 4667 8996 4712 9024
rect 4706 8984 4712 8996
rect 4764 8984 4770 9036
rect 7006 9024 7012 9036
rect 5276 8996 7012 9024
rect 1946 8956 1952 8968
rect 1907 8928 1952 8956
rect 1946 8916 1952 8928
rect 2004 8916 2010 8968
rect 2774 8916 2780 8968
rect 2832 8956 2838 8968
rect 3237 8959 3295 8965
rect 2832 8928 2877 8956
rect 2832 8916 2838 8928
rect 3237 8925 3249 8959
rect 3283 8956 3295 8959
rect 3510 8956 3516 8968
rect 3283 8928 3516 8956
rect 3283 8925 3295 8928
rect 3237 8919 3295 8925
rect 3510 8916 3516 8928
rect 3568 8916 3574 8968
rect 3973 8959 4031 8965
rect 3973 8925 3985 8959
rect 4019 8956 4031 8959
rect 4062 8956 4068 8968
rect 4019 8928 4068 8956
rect 4019 8925 4031 8928
rect 3973 8919 4031 8925
rect 4062 8916 4068 8928
rect 4120 8956 4126 8968
rect 5276 8956 5304 8996
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 9766 8984 9772 9036
rect 9824 9024 9830 9036
rect 9953 9027 10011 9033
rect 9953 9024 9965 9027
rect 9824 8996 9965 9024
rect 9824 8984 9830 8996
rect 9953 8993 9965 8996
rect 9999 8993 10011 9027
rect 10060 9024 10088 9064
rect 11256 9064 11713 9092
rect 11256 9024 11284 9064
rect 11701 9061 11713 9064
rect 11747 9092 11759 9095
rect 11882 9092 11888 9104
rect 11747 9064 11888 9092
rect 11747 9061 11759 9064
rect 11701 9055 11759 9061
rect 11882 9052 11888 9064
rect 11940 9052 11946 9104
rect 12526 9052 12532 9104
rect 12584 9092 12590 9104
rect 12584 9064 14412 9092
rect 12584 9052 12590 9064
rect 13722 9024 13728 9036
rect 10060 8996 11284 9024
rect 11348 8996 13728 9024
rect 9953 8987 10011 8993
rect 4120 8928 5304 8956
rect 5353 8959 5411 8965
rect 4120 8916 4126 8928
rect 5353 8925 5365 8959
rect 5399 8925 5411 8959
rect 5353 8919 5411 8925
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8956 6607 8959
rect 6638 8956 6644 8968
rect 6595 8928 6644 8956
rect 6595 8925 6607 8928
rect 6549 8919 6607 8925
rect 3694 8848 3700 8900
rect 3752 8888 3758 8900
rect 5368 8888 5396 8919
rect 6638 8916 6644 8928
rect 6696 8916 6702 8968
rect 6914 8916 6920 8968
rect 6972 8956 6978 8968
rect 8202 8956 8208 8968
rect 6972 8928 8208 8956
rect 6972 8916 6978 8928
rect 8202 8916 8208 8928
rect 8260 8956 8266 8968
rect 8389 8959 8447 8965
rect 8389 8956 8401 8959
rect 8260 8928 8401 8956
rect 8260 8916 8266 8928
rect 8389 8925 8401 8928
rect 8435 8925 8447 8959
rect 8389 8919 8447 8925
rect 9309 8959 9367 8965
rect 9309 8925 9321 8959
rect 9355 8956 9367 8959
rect 9858 8956 9864 8968
rect 9355 8928 9864 8956
rect 9355 8925 9367 8928
rect 9309 8919 9367 8925
rect 9858 8916 9864 8928
rect 9916 8916 9922 8968
rect 11348 8942 11376 8996
rect 13722 8984 13728 8996
rect 13780 8984 13786 9036
rect 13814 8984 13820 9036
rect 13872 9024 13878 9036
rect 14277 9027 14335 9033
rect 14277 9024 14289 9027
rect 13872 8996 14289 9024
rect 13872 8984 13878 8996
rect 14277 8993 14289 8996
rect 14323 8993 14335 9027
rect 14384 9024 14412 9064
rect 15838 9052 15844 9104
rect 15896 9092 15902 9104
rect 15896 9064 16988 9092
rect 15896 9052 15902 9064
rect 15562 9024 15568 9036
rect 14384 8996 15568 9024
rect 14277 8987 14335 8993
rect 15562 8984 15568 8996
rect 15620 8984 15626 9036
rect 16040 9033 16068 9064
rect 16025 9027 16083 9033
rect 16025 8993 16037 9027
rect 16071 8993 16083 9027
rect 16025 8987 16083 8993
rect 16577 9027 16635 9033
rect 16577 8993 16589 9027
rect 16623 9024 16635 9027
rect 16850 9024 16856 9036
rect 16623 8996 16856 9024
rect 16623 8993 16635 8996
rect 16577 8987 16635 8993
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 16960 9024 16988 9064
rect 17218 9052 17224 9104
rect 17276 9092 17282 9104
rect 23308 9092 23336 9132
rect 23474 9120 23480 9132
rect 23532 9120 23538 9172
rect 25038 9092 25044 9104
rect 17276 9064 23244 9092
rect 23308 9064 25044 9092
rect 17276 9052 17282 9064
rect 17402 9024 17408 9036
rect 16960 8996 17408 9024
rect 17402 8984 17408 8996
rect 17460 8984 17466 9036
rect 17512 8996 23152 9024
rect 12342 8916 12348 8968
rect 12400 8956 12406 8968
rect 12529 8959 12587 8965
rect 12529 8956 12541 8959
rect 12400 8928 12541 8956
rect 12400 8916 12406 8928
rect 12529 8925 12541 8928
rect 12575 8925 12587 8959
rect 12529 8919 12587 8925
rect 13173 8959 13231 8965
rect 13173 8925 13185 8959
rect 13219 8956 13231 8959
rect 13906 8956 13912 8968
rect 13219 8928 13912 8956
rect 13219 8925 13231 8928
rect 13173 8919 13231 8925
rect 13906 8916 13912 8928
rect 13964 8916 13970 8968
rect 6730 8888 6736 8900
rect 3752 8860 6736 8888
rect 3752 8848 3758 8860
rect 6730 8848 6736 8860
rect 6788 8848 6794 8900
rect 7006 8848 7012 8900
rect 7064 8888 7070 8900
rect 7653 8891 7711 8897
rect 7653 8888 7665 8891
rect 7064 8860 7665 8888
rect 7064 8848 7070 8860
rect 7653 8857 7665 8860
rect 7699 8857 7711 8891
rect 9674 8888 9680 8900
rect 7653 8851 7711 8857
rect 7760 8860 9680 8888
rect 2774 8780 2780 8832
rect 2832 8820 2838 8832
rect 3234 8820 3240 8832
rect 2832 8792 3240 8820
rect 2832 8780 2838 8792
rect 3234 8780 3240 8792
rect 3292 8780 3298 8832
rect 6086 8780 6092 8832
rect 6144 8820 6150 8832
rect 7760 8820 7788 8860
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 9950 8848 9956 8900
rect 10008 8888 10014 8900
rect 10229 8891 10287 8897
rect 10229 8888 10241 8891
rect 10008 8860 10241 8888
rect 10008 8848 10014 8860
rect 10229 8857 10241 8860
rect 10275 8857 10287 8891
rect 10229 8851 10287 8857
rect 12158 8848 12164 8900
rect 12216 8888 12222 8900
rect 14458 8888 14464 8900
rect 12216 8860 14464 8888
rect 12216 8848 12222 8860
rect 14458 8848 14464 8860
rect 14516 8848 14522 8900
rect 14553 8891 14611 8897
rect 14553 8857 14565 8891
rect 14599 8888 14611 8891
rect 14826 8888 14832 8900
rect 14599 8860 14832 8888
rect 14599 8857 14611 8860
rect 14553 8851 14611 8857
rect 14826 8848 14832 8860
rect 14884 8848 14890 8900
rect 15838 8888 15844 8900
rect 15778 8860 15844 8888
rect 15838 8848 15844 8860
rect 15896 8848 15902 8900
rect 16669 8891 16727 8897
rect 16669 8857 16681 8891
rect 16715 8888 16727 8891
rect 17512 8888 17540 8996
rect 19705 8959 19763 8965
rect 19705 8925 19717 8959
rect 19751 8956 19763 8959
rect 20530 8956 20536 8968
rect 19751 8928 20536 8956
rect 19751 8925 19763 8928
rect 19705 8919 19763 8925
rect 20530 8916 20536 8928
rect 20588 8916 20594 8968
rect 21634 8916 21640 8968
rect 21692 8956 21698 8968
rect 21692 8928 21737 8956
rect 21692 8916 21698 8928
rect 22094 8916 22100 8968
rect 22152 8956 22158 8968
rect 22738 8956 22744 8968
rect 22152 8928 22197 8956
rect 22699 8928 22744 8956
rect 22152 8916 22158 8928
rect 22738 8916 22744 8928
rect 22796 8916 22802 8968
rect 16715 8860 17540 8888
rect 17589 8891 17647 8897
rect 16715 8857 16727 8860
rect 16669 8851 16727 8857
rect 17589 8857 17601 8891
rect 17635 8888 17647 8891
rect 17678 8888 17684 8900
rect 17635 8860 17684 8888
rect 17635 8857 17647 8860
rect 17589 8851 17647 8857
rect 17678 8848 17684 8860
rect 17736 8848 17742 8900
rect 18138 8888 18144 8900
rect 18099 8860 18144 8888
rect 18138 8848 18144 8860
rect 18196 8848 18202 8900
rect 18233 8891 18291 8897
rect 18233 8857 18245 8891
rect 18279 8857 18291 8891
rect 18233 8851 18291 8857
rect 6144 8792 7788 8820
rect 9401 8823 9459 8829
rect 6144 8780 6150 8792
rect 9401 8789 9413 8823
rect 9447 8820 9459 8823
rect 10318 8820 10324 8832
rect 9447 8792 10324 8820
rect 9447 8789 9459 8792
rect 9401 8783 9459 8789
rect 10318 8780 10324 8792
rect 10376 8780 10382 8832
rect 11054 8780 11060 8832
rect 11112 8820 11118 8832
rect 12434 8820 12440 8832
rect 11112 8792 12440 8820
rect 11112 8780 11118 8792
rect 12434 8780 12440 8792
rect 12492 8780 12498 8832
rect 12526 8780 12532 8832
rect 12584 8820 12590 8832
rect 17862 8820 17868 8832
rect 12584 8792 17868 8820
rect 12584 8780 12590 8792
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 18248 8820 18276 8851
rect 18506 8848 18512 8900
rect 18564 8888 18570 8900
rect 18785 8891 18843 8897
rect 18785 8888 18797 8891
rect 18564 8860 18797 8888
rect 18564 8848 18570 8860
rect 18785 8857 18797 8860
rect 18831 8857 18843 8891
rect 18785 8851 18843 8857
rect 19150 8848 19156 8900
rect 19208 8888 19214 8900
rect 20990 8888 20996 8900
rect 19208 8860 19932 8888
rect 20951 8860 20996 8888
rect 19208 8848 19214 8860
rect 19797 8823 19855 8829
rect 19797 8820 19809 8823
rect 18248 8792 19809 8820
rect 19797 8789 19809 8792
rect 19843 8789 19855 8823
rect 19904 8820 19932 8860
rect 20990 8848 20996 8860
rect 21048 8848 21054 8900
rect 21085 8891 21143 8897
rect 21085 8857 21097 8891
rect 21131 8857 21143 8891
rect 21085 8851 21143 8857
rect 20898 8820 20904 8832
rect 19904 8792 20904 8820
rect 19797 8783 19855 8789
rect 20898 8780 20904 8792
rect 20956 8780 20962 8832
rect 21100 8820 21128 8851
rect 22189 8823 22247 8829
rect 22189 8820 22201 8823
rect 21100 8792 22201 8820
rect 22189 8789 22201 8792
rect 22235 8789 22247 8823
rect 22830 8820 22836 8832
rect 22791 8792 22836 8820
rect 22189 8783 22247 8789
rect 22830 8780 22836 8792
rect 22888 8780 22894 8832
rect 23124 8820 23152 8996
rect 23216 8956 23244 9064
rect 25038 9052 25044 9064
rect 25096 9052 25102 9104
rect 23385 8959 23443 8965
rect 23385 8956 23397 8959
rect 23216 8928 23397 8956
rect 23385 8925 23397 8928
rect 23431 8925 23443 8959
rect 24578 8956 24584 8968
rect 24539 8928 24584 8956
rect 23385 8919 23443 8925
rect 23400 8888 23428 8919
rect 24578 8916 24584 8928
rect 24636 8916 24642 8968
rect 25222 8888 25228 8900
rect 23400 8860 25228 8888
rect 25222 8848 25228 8860
rect 25280 8848 25286 8900
rect 24673 8823 24731 8829
rect 24673 8820 24685 8823
rect 23124 8792 24685 8820
rect 24673 8789 24685 8792
rect 24719 8789 24731 8823
rect 24673 8783 24731 8789
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 1946 8576 1952 8628
rect 2004 8616 2010 8628
rect 5077 8619 5135 8625
rect 5077 8616 5089 8619
rect 2004 8588 5089 8616
rect 2004 8576 2010 8588
rect 5077 8585 5089 8588
rect 5123 8585 5135 8619
rect 5077 8579 5135 8585
rect 7098 8576 7104 8628
rect 7156 8616 7162 8628
rect 7193 8619 7251 8625
rect 7193 8616 7205 8619
rect 7156 8588 7205 8616
rect 7156 8576 7162 8588
rect 7193 8585 7205 8588
rect 7239 8585 7251 8619
rect 11054 8616 11060 8628
rect 7193 8579 7251 8585
rect 9692 8588 11060 8616
rect 2774 8548 2780 8560
rect 2240 8520 2780 8548
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8480 1823 8483
rect 2240 8480 2268 8520
rect 2774 8508 2780 8520
rect 2832 8508 2838 8560
rect 3510 8508 3516 8560
rect 3568 8508 3574 8560
rect 3970 8508 3976 8560
rect 4028 8548 4034 8560
rect 4028 8520 5304 8548
rect 4028 8508 4034 8520
rect 1811 8452 2268 8480
rect 4433 8483 4491 8489
rect 1811 8449 1823 8452
rect 1765 8443 1823 8449
rect 4433 8449 4445 8483
rect 4479 8449 4491 8483
rect 4433 8443 4491 8449
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8480 4583 8483
rect 4798 8480 4804 8492
rect 4571 8452 4804 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 1670 8372 1676 8424
rect 1728 8412 1734 8424
rect 2225 8415 2283 8421
rect 2225 8412 2237 8415
rect 1728 8384 2237 8412
rect 1728 8372 1734 8384
rect 2225 8381 2237 8384
rect 2271 8381 2283 8415
rect 2225 8375 2283 8381
rect 2501 8415 2559 8421
rect 2501 8381 2513 8415
rect 2547 8412 2559 8415
rect 4448 8412 4476 8443
rect 4798 8440 4804 8452
rect 4856 8440 4862 8492
rect 5276 8489 5304 8520
rect 5350 8508 5356 8560
rect 5408 8548 5414 8560
rect 9692 8557 9720 8588
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 11624 8588 12434 8616
rect 9677 8551 9735 8557
rect 5408 8520 7420 8548
rect 5408 8508 5414 8520
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8449 5319 8483
rect 5261 8443 5319 8449
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8480 6607 8483
rect 6730 8480 6736 8492
rect 6595 8452 6736 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 7392 8489 7420 8520
rect 9677 8517 9689 8551
rect 9723 8517 9735 8551
rect 9677 8511 9735 8517
rect 10686 8508 10692 8560
rect 10744 8508 10750 8560
rect 7377 8483 7435 8489
rect 7377 8449 7389 8483
rect 7423 8449 7435 8483
rect 8757 8483 8815 8489
rect 8757 8480 8769 8483
rect 7377 8443 7435 8449
rect 8036 8452 8769 8480
rect 4706 8412 4712 8424
rect 2547 8384 4200 8412
rect 4448 8384 4712 8412
rect 2547 8381 2559 8384
rect 2501 8375 2559 8381
rect 750 8304 756 8356
rect 808 8344 814 8356
rect 4172 8344 4200 8384
rect 4706 8372 4712 8384
rect 4764 8372 4770 8424
rect 4890 8372 4896 8424
rect 4948 8412 4954 8424
rect 6641 8415 6699 8421
rect 6641 8412 6653 8415
rect 4948 8384 6653 8412
rect 4948 8372 4954 8384
rect 6641 8381 6653 8384
rect 6687 8381 6699 8415
rect 6641 8375 6699 8381
rect 5442 8344 5448 8356
rect 808 8316 1072 8344
rect 4172 8316 5448 8344
rect 808 8304 814 8316
rect 1044 8072 1072 8316
rect 5442 8304 5448 8316
rect 5500 8304 5506 8356
rect 7834 8344 7840 8356
rect 5552 8316 7840 8344
rect 3970 8276 3976 8288
rect 3931 8248 3976 8276
rect 3970 8236 3976 8248
rect 4028 8236 4034 8288
rect 4706 8236 4712 8288
rect 4764 8276 4770 8288
rect 5552 8276 5580 8316
rect 7834 8304 7840 8316
rect 7892 8344 7898 8356
rect 8036 8344 8064 8452
rect 8757 8449 8769 8452
rect 8803 8449 8815 8483
rect 11624 8480 11652 8588
rect 11974 8548 11980 8560
rect 11716 8520 11980 8548
rect 11716 8489 11744 8520
rect 11974 8508 11980 8520
rect 12032 8508 12038 8560
rect 12406 8548 12434 8588
rect 12618 8576 12624 8628
rect 12676 8616 12682 8628
rect 13630 8616 13636 8628
rect 12676 8588 13636 8616
rect 12676 8576 12682 8588
rect 13630 8576 13636 8588
rect 13688 8576 13694 8628
rect 17218 8616 17224 8628
rect 13740 8588 17224 8616
rect 12406 8520 12466 8548
rect 8757 8443 8815 8449
rect 10888 8452 11652 8480
rect 11701 8483 11759 8489
rect 8202 8372 8208 8424
rect 8260 8412 8266 8424
rect 9401 8415 9459 8421
rect 9401 8412 9413 8415
rect 8260 8384 9413 8412
rect 8260 8372 8266 8384
rect 9401 8381 9413 8384
rect 9447 8381 9459 8415
rect 10134 8412 10140 8424
rect 9401 8375 9459 8381
rect 9508 8384 10140 8412
rect 7892 8316 8064 8344
rect 8849 8347 8907 8353
rect 7892 8304 7898 8316
rect 8849 8313 8861 8347
rect 8895 8344 8907 8347
rect 9508 8344 9536 8384
rect 10134 8372 10140 8384
rect 10192 8372 10198 8424
rect 10226 8372 10232 8424
rect 10284 8412 10290 8424
rect 10888 8412 10916 8452
rect 11701 8449 11713 8483
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 10284 8384 10916 8412
rect 11149 8415 11207 8421
rect 10284 8372 10290 8384
rect 11149 8381 11161 8415
rect 11195 8412 11207 8415
rect 11977 8415 12035 8421
rect 11977 8412 11989 8415
rect 11195 8384 11989 8412
rect 11195 8381 11207 8384
rect 11149 8375 11207 8381
rect 11977 8381 11989 8384
rect 12023 8412 12035 8415
rect 13740 8412 13768 8588
rect 17218 8576 17224 8588
rect 17276 8576 17282 8628
rect 17402 8576 17408 8628
rect 17460 8616 17466 8628
rect 17460 8588 17724 8616
rect 17460 8576 17466 8588
rect 15562 8548 15568 8560
rect 15410 8520 15568 8548
rect 15562 8508 15568 8520
rect 15620 8508 15626 8560
rect 16298 8508 16304 8560
rect 16356 8548 16362 8560
rect 17037 8551 17095 8557
rect 17037 8548 17049 8551
rect 16356 8520 17049 8548
rect 16356 8508 16362 8520
rect 17037 8517 17049 8520
rect 17083 8517 17095 8551
rect 17586 8548 17592 8560
rect 17547 8520 17592 8548
rect 17037 8511 17095 8517
rect 17586 8508 17592 8520
rect 17644 8508 17650 8560
rect 13814 8440 13820 8492
rect 13872 8480 13878 8492
rect 13909 8483 13967 8489
rect 13909 8480 13921 8483
rect 13872 8452 13921 8480
rect 13872 8440 13878 8452
rect 13909 8449 13921 8452
rect 13955 8449 13967 8483
rect 13909 8443 13967 8449
rect 15470 8440 15476 8492
rect 15528 8480 15534 8492
rect 16117 8483 16175 8489
rect 16117 8480 16129 8483
rect 15528 8452 16129 8480
rect 15528 8440 15534 8452
rect 16117 8449 16129 8452
rect 16163 8449 16175 8483
rect 16117 8443 16175 8449
rect 12023 8384 13768 8412
rect 14185 8415 14243 8421
rect 12023 8381 12035 8384
rect 11977 8375 12035 8381
rect 14185 8381 14197 8415
rect 14231 8412 14243 8415
rect 16209 8415 16267 8421
rect 14231 8384 16160 8412
rect 14231 8381 14243 8384
rect 14185 8375 14243 8381
rect 16132 8356 16160 8384
rect 16209 8381 16221 8415
rect 16255 8412 16267 8415
rect 16390 8412 16396 8424
rect 16255 8384 16396 8412
rect 16255 8381 16267 8384
rect 16209 8375 16267 8381
rect 16390 8372 16396 8384
rect 16448 8372 16454 8424
rect 16945 8415 17003 8421
rect 16945 8381 16957 8415
rect 16991 8381 17003 8415
rect 17696 8412 17724 8588
rect 18138 8576 18144 8628
rect 18196 8616 18202 8628
rect 20438 8616 20444 8628
rect 18196 8588 20444 8616
rect 18196 8576 18202 8588
rect 20438 8576 20444 8588
rect 20496 8576 20502 8628
rect 20990 8576 20996 8628
rect 21048 8616 21054 8628
rect 30006 8616 30012 8628
rect 21048 8588 30012 8616
rect 21048 8576 21054 8588
rect 30006 8576 30012 8588
rect 30064 8576 30070 8628
rect 17862 8508 17868 8560
rect 17920 8548 17926 8560
rect 18325 8551 18383 8557
rect 18325 8548 18337 8551
rect 17920 8520 18337 8548
rect 17920 8508 17926 8520
rect 18325 8517 18337 8520
rect 18371 8548 18383 8551
rect 19334 8548 19340 8560
rect 18371 8520 19340 8548
rect 18371 8517 18383 8520
rect 18325 8511 18383 8517
rect 19334 8508 19340 8520
rect 19392 8508 19398 8560
rect 19429 8551 19487 8557
rect 19429 8517 19441 8551
rect 19475 8548 19487 8551
rect 22830 8548 22836 8560
rect 19475 8520 22836 8548
rect 19475 8517 19487 8520
rect 19429 8511 19487 8517
rect 22830 8508 22836 8520
rect 22888 8508 22894 8560
rect 38289 8551 38347 8557
rect 38289 8517 38301 8551
rect 38335 8548 38347 8551
rect 38378 8548 38384 8560
rect 38335 8520 38384 8548
rect 38335 8517 38347 8520
rect 38289 8511 38347 8517
rect 38378 8508 38384 8520
rect 38436 8508 38442 8560
rect 18046 8480 18052 8492
rect 18007 8452 18052 8480
rect 18046 8440 18052 8452
rect 18104 8440 18110 8492
rect 18690 8440 18696 8492
rect 18748 8480 18754 8492
rect 18966 8480 18972 8492
rect 18748 8452 18972 8480
rect 18748 8440 18754 8452
rect 18966 8440 18972 8452
rect 19024 8440 19030 8492
rect 22370 8480 22376 8492
rect 20364 8452 22376 8480
rect 19334 8412 19340 8424
rect 17696 8384 18552 8412
rect 19295 8384 19340 8412
rect 16945 8375 17003 8381
rect 13449 8347 13507 8353
rect 8895 8316 9536 8344
rect 10704 8316 11836 8344
rect 8895 8313 8907 8316
rect 8849 8307 8907 8313
rect 4764 8248 5580 8276
rect 4764 8236 4770 8248
rect 10134 8236 10140 8288
rect 10192 8276 10198 8288
rect 10704 8276 10732 8316
rect 10192 8248 10732 8276
rect 11808 8276 11836 8316
rect 13449 8313 13461 8347
rect 13495 8344 13507 8347
rect 13495 8316 14044 8344
rect 13495 8313 13507 8316
rect 13449 8307 13507 8313
rect 12526 8276 12532 8288
rect 11808 8248 12532 8276
rect 10192 8236 10198 8248
rect 12526 8236 12532 8248
rect 12584 8236 12590 8288
rect 14016 8276 14044 8316
rect 16114 8304 16120 8356
rect 16172 8304 16178 8356
rect 14274 8276 14280 8288
rect 14016 8248 14280 8276
rect 14274 8236 14280 8248
rect 14332 8276 14338 8288
rect 14918 8276 14924 8288
rect 14332 8248 14924 8276
rect 14332 8236 14338 8248
rect 14918 8236 14924 8248
rect 14976 8236 14982 8288
rect 15194 8236 15200 8288
rect 15252 8276 15258 8288
rect 15657 8279 15715 8285
rect 15657 8276 15669 8279
rect 15252 8248 15669 8276
rect 15252 8236 15258 8248
rect 15657 8245 15669 8248
rect 15703 8276 15715 8279
rect 16022 8276 16028 8288
rect 15703 8248 16028 8276
rect 15703 8245 15715 8248
rect 15657 8239 15715 8245
rect 16022 8236 16028 8248
rect 16080 8236 16086 8288
rect 16960 8276 16988 8375
rect 18524 8344 18552 8384
rect 19334 8372 19340 8384
rect 19392 8372 19398 8424
rect 20364 8421 20392 8452
rect 22370 8440 22376 8452
rect 22428 8440 22434 8492
rect 22646 8480 22652 8492
rect 22607 8452 22652 8480
rect 22646 8440 22652 8452
rect 22704 8440 22710 8492
rect 23290 8480 23296 8492
rect 23251 8452 23296 8480
rect 23290 8440 23296 8452
rect 23348 8440 23354 8492
rect 23382 8440 23388 8492
rect 23440 8480 23446 8492
rect 23937 8483 23995 8489
rect 23937 8480 23949 8483
rect 23440 8452 23949 8480
rect 23440 8440 23446 8452
rect 23937 8449 23949 8452
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 24026 8440 24032 8492
rect 24084 8480 24090 8492
rect 24581 8483 24639 8489
rect 24581 8480 24593 8483
rect 24084 8452 24593 8480
rect 24084 8440 24090 8452
rect 24581 8449 24593 8452
rect 24627 8449 24639 8483
rect 25222 8480 25228 8492
rect 25183 8452 25228 8480
rect 24581 8443 24639 8449
rect 25222 8440 25228 8452
rect 25280 8440 25286 8492
rect 38102 8480 38108 8492
rect 38063 8452 38108 8480
rect 38102 8440 38108 8452
rect 38160 8440 38166 8492
rect 20349 8415 20407 8421
rect 20349 8381 20361 8415
rect 20395 8381 20407 8415
rect 20349 8375 20407 8381
rect 20806 8372 20812 8424
rect 20864 8412 20870 8424
rect 20993 8415 21051 8421
rect 20993 8412 21005 8415
rect 20864 8384 21005 8412
rect 20864 8372 20870 8384
rect 20993 8381 21005 8384
rect 21039 8381 21051 8415
rect 22002 8412 22008 8424
rect 21963 8384 22008 8412
rect 20993 8375 21051 8381
rect 22002 8372 22008 8384
rect 22060 8372 22066 8424
rect 22738 8412 22744 8424
rect 22699 8384 22744 8412
rect 22738 8372 22744 8384
rect 22796 8372 22802 8424
rect 20622 8344 20628 8356
rect 18524 8316 20628 8344
rect 20622 8304 20628 8316
rect 20680 8304 20686 8356
rect 20714 8304 20720 8356
rect 20772 8344 20778 8356
rect 24029 8347 24087 8353
rect 24029 8344 24041 8347
rect 20772 8316 24041 8344
rect 20772 8304 20778 8316
rect 24029 8313 24041 8316
rect 24075 8313 24087 8347
rect 25314 8344 25320 8356
rect 25275 8316 25320 8344
rect 24029 8307 24087 8313
rect 25314 8304 25320 8316
rect 25372 8304 25378 8356
rect 18230 8276 18236 8288
rect 16960 8248 18236 8276
rect 18230 8236 18236 8248
rect 18288 8236 18294 8288
rect 18690 8236 18696 8288
rect 18748 8276 18754 8288
rect 21082 8276 21088 8288
rect 18748 8248 21088 8276
rect 18748 8236 18754 8248
rect 21082 8236 21088 8248
rect 21140 8236 21146 8288
rect 21174 8236 21180 8288
rect 21232 8276 21238 8288
rect 21910 8276 21916 8288
rect 21232 8248 21916 8276
rect 21232 8236 21238 8248
rect 21910 8236 21916 8248
rect 21968 8236 21974 8288
rect 22830 8236 22836 8288
rect 22888 8276 22894 8288
rect 23385 8279 23443 8285
rect 23385 8276 23397 8279
rect 22888 8248 23397 8276
rect 22888 8236 22894 8248
rect 23385 8245 23397 8248
rect 23431 8245 23443 8279
rect 24670 8276 24676 8288
rect 24631 8248 24676 8276
rect 23385 8239 23443 8245
rect 24670 8236 24676 8248
rect 24728 8236 24734 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 3418 8072 3424 8084
rect 1044 8044 1808 8072
rect 3379 8044 3424 8072
rect 1670 7936 1676 7948
rect 1631 7908 1676 7936
rect 1670 7896 1676 7908
rect 1728 7896 1734 7948
rect 1780 7936 1808 8044
rect 3418 8032 3424 8044
rect 3476 8032 3482 8084
rect 5994 8072 6000 8084
rect 5955 8044 6000 8072
rect 5994 8032 6000 8044
rect 6052 8032 6058 8084
rect 6825 8075 6883 8081
rect 6825 8041 6837 8075
rect 6871 8072 6883 8075
rect 7190 8072 7196 8084
rect 6871 8044 7196 8072
rect 6871 8041 6883 8044
rect 6825 8035 6883 8041
rect 7190 8032 7196 8044
rect 7248 8032 7254 8084
rect 11333 8075 11391 8081
rect 11333 8041 11345 8075
rect 11379 8072 11391 8075
rect 12066 8072 12072 8084
rect 11379 8044 12072 8072
rect 11379 8041 11391 8044
rect 11333 8035 11391 8041
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 12710 8032 12716 8084
rect 12768 8072 12774 8084
rect 16025 8075 16083 8081
rect 12768 8044 15608 8072
rect 12768 8032 12774 8044
rect 11606 7964 11612 8016
rect 11664 8004 11670 8016
rect 11701 8007 11759 8013
rect 11701 8004 11713 8007
rect 11664 7976 11713 8004
rect 11664 7964 11670 7976
rect 11701 7973 11713 7976
rect 11747 8004 11759 8007
rect 15580 8004 15608 8044
rect 16025 8041 16037 8075
rect 16071 8072 16083 8075
rect 16114 8072 16120 8084
rect 16071 8044 16120 8072
rect 16071 8041 16083 8044
rect 16025 8035 16083 8041
rect 16114 8032 16120 8044
rect 16172 8032 16178 8084
rect 16224 8044 19840 8072
rect 16224 8004 16252 8044
rect 18322 8004 18328 8016
rect 11747 7976 12112 8004
rect 15580 7976 16252 8004
rect 17604 7976 18328 8004
rect 11747 7973 11759 7976
rect 11701 7967 11759 7973
rect 1949 7939 2007 7945
rect 1949 7936 1961 7939
rect 1780 7908 1961 7936
rect 1949 7905 1961 7908
rect 1995 7936 2007 7939
rect 3970 7936 3976 7948
rect 1995 7908 3976 7936
rect 1995 7905 2007 7908
rect 1949 7899 2007 7905
rect 3970 7896 3976 7908
rect 4028 7896 4034 7948
rect 9861 7939 9919 7945
rect 9861 7905 9873 7939
rect 9907 7936 9919 7939
rect 11974 7936 11980 7948
rect 9907 7908 11836 7936
rect 11935 7908 11980 7936
rect 9907 7905 9919 7908
rect 9861 7899 9919 7905
rect 4065 7871 4123 7877
rect 4065 7837 4077 7871
rect 4111 7868 4123 7871
rect 4706 7868 4712 7880
rect 4111 7840 4712 7868
rect 4111 7837 4123 7840
rect 4065 7831 4123 7837
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 5905 7871 5963 7877
rect 5905 7837 5917 7871
rect 5951 7837 5963 7871
rect 5905 7831 5963 7837
rect 3970 7800 3976 7812
rect 3174 7772 3976 7800
rect 3970 7760 3976 7772
rect 4028 7760 4034 7812
rect 5534 7760 5540 7812
rect 5592 7800 5598 7812
rect 5920 7800 5948 7831
rect 6638 7828 6644 7880
rect 6696 7868 6702 7880
rect 6733 7871 6791 7877
rect 6733 7868 6745 7871
rect 6696 7840 6745 7868
rect 6696 7828 6702 7840
rect 6733 7837 6745 7840
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 9030 7828 9036 7880
rect 9088 7868 9094 7880
rect 9585 7871 9643 7877
rect 9585 7868 9597 7871
rect 9088 7840 9597 7868
rect 9088 7828 9094 7840
rect 9585 7837 9597 7840
rect 9631 7837 9643 7871
rect 9585 7831 9643 7837
rect 6454 7800 6460 7812
rect 5592 7772 6460 7800
rect 5592 7760 5598 7772
rect 6454 7760 6460 7772
rect 6512 7800 6518 7812
rect 9766 7800 9772 7812
rect 6512 7772 9772 7800
rect 6512 7760 6518 7772
rect 9766 7760 9772 7772
rect 9824 7760 9830 7812
rect 10318 7760 10324 7812
rect 10376 7760 10382 7812
rect 4154 7732 4160 7744
rect 4115 7704 4160 7732
rect 4154 7692 4160 7704
rect 4212 7692 4218 7744
rect 5442 7692 5448 7744
rect 5500 7732 5506 7744
rect 11606 7732 11612 7744
rect 5500 7704 11612 7732
rect 5500 7692 5506 7704
rect 11606 7692 11612 7704
rect 11664 7692 11670 7744
rect 11808 7732 11836 7908
rect 11974 7896 11980 7908
rect 12032 7896 12038 7948
rect 12084 7936 12112 7976
rect 12253 7939 12311 7945
rect 12253 7936 12265 7939
rect 12084 7908 12265 7936
rect 12253 7905 12265 7908
rect 12299 7936 12311 7939
rect 14090 7936 14096 7948
rect 12299 7908 14096 7936
rect 12299 7905 12311 7908
rect 12253 7899 12311 7905
rect 14090 7896 14096 7908
rect 14148 7896 14154 7948
rect 14553 7939 14611 7945
rect 14553 7905 14565 7939
rect 14599 7936 14611 7939
rect 16390 7936 16396 7948
rect 14599 7908 16396 7936
rect 14599 7905 14611 7908
rect 14553 7899 14611 7905
rect 16390 7896 16396 7908
rect 16448 7896 16454 7948
rect 17604 7945 17632 7976
rect 18322 7964 18328 7976
rect 18380 8004 18386 8016
rect 19242 8004 19248 8016
rect 18380 7976 19248 8004
rect 18380 7964 18386 7976
rect 19242 7964 19248 7976
rect 19300 7964 19306 8016
rect 19812 8004 19840 8044
rect 19886 8032 19892 8084
rect 19944 8072 19950 8084
rect 23934 8072 23940 8084
rect 19944 8044 23940 8072
rect 19944 8032 19950 8044
rect 23934 8032 23940 8044
rect 23992 8072 23998 8084
rect 23992 8044 24808 8072
rect 23992 8032 23998 8044
rect 23290 8004 23296 8016
rect 19812 7976 23296 8004
rect 23290 7964 23296 7976
rect 23348 7964 23354 8016
rect 16577 7939 16635 7945
rect 16577 7905 16589 7939
rect 16623 7936 16635 7939
rect 17589 7939 17647 7945
rect 16623 7908 17540 7936
rect 16623 7905 16635 7908
rect 16577 7899 16635 7905
rect 13722 7828 13728 7880
rect 13780 7868 13786 7880
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 13780 7840 14289 7868
rect 13780 7828 13786 7840
rect 14277 7837 14289 7840
rect 14323 7837 14335 7871
rect 17512 7868 17540 7908
rect 17589 7905 17601 7939
rect 17635 7905 17647 7939
rect 19518 7936 19524 7948
rect 17589 7899 17647 7905
rect 18064 7908 19334 7936
rect 19479 7908 19524 7936
rect 17862 7868 17868 7880
rect 17512 7840 17868 7868
rect 14277 7831 14335 7837
rect 17862 7828 17868 7840
rect 17920 7828 17926 7880
rect 14826 7800 14832 7812
rect 13478 7772 14832 7800
rect 14826 7760 14832 7772
rect 14884 7760 14890 7812
rect 16390 7800 16396 7812
rect 15778 7772 16396 7800
rect 16390 7760 16396 7772
rect 16448 7760 16454 7812
rect 16666 7760 16672 7812
rect 16724 7800 16730 7812
rect 16724 7772 16769 7800
rect 16724 7760 16730 7772
rect 12894 7732 12900 7744
rect 11808 7704 12900 7732
rect 12894 7692 12900 7704
rect 12952 7692 12958 7744
rect 13725 7735 13783 7741
rect 13725 7701 13737 7735
rect 13771 7732 13783 7735
rect 14550 7732 14556 7744
rect 13771 7704 14556 7732
rect 13771 7701 13783 7704
rect 13725 7695 13783 7701
rect 14550 7692 14556 7704
rect 14608 7732 14614 7744
rect 18064 7732 18092 7908
rect 18230 7800 18236 7812
rect 18191 7772 18236 7800
rect 18230 7760 18236 7772
rect 18288 7760 18294 7812
rect 18334 7803 18392 7809
rect 18334 7769 18346 7803
rect 18380 7800 18392 7803
rect 18877 7803 18935 7809
rect 18380 7772 18460 7800
rect 18380 7769 18392 7772
rect 18334 7763 18392 7769
rect 14608 7704 18092 7732
rect 18432 7732 18460 7772
rect 18877 7769 18889 7803
rect 18923 7800 18935 7803
rect 19058 7800 19064 7812
rect 18923 7772 19064 7800
rect 18923 7769 18935 7772
rect 18877 7763 18935 7769
rect 19058 7760 19064 7772
rect 19116 7760 19122 7812
rect 19306 7800 19334 7908
rect 19518 7896 19524 7908
rect 19576 7896 19582 7948
rect 20165 7939 20223 7945
rect 20165 7905 20177 7939
rect 20211 7936 20223 7939
rect 22002 7936 22008 7948
rect 20211 7908 22008 7936
rect 20211 7905 20223 7908
rect 20165 7899 20223 7905
rect 22002 7896 22008 7908
rect 22060 7896 22066 7948
rect 22094 7896 22100 7948
rect 22152 7936 22158 7948
rect 22152 7908 23244 7936
rect 22152 7896 22158 7908
rect 19426 7868 19432 7880
rect 19387 7840 19432 7868
rect 19426 7828 19432 7840
rect 19484 7828 19490 7880
rect 23216 7877 23244 7908
rect 23201 7871 23259 7877
rect 22756 7868 22968 7870
rect 22572 7842 23060 7868
rect 22572 7840 22784 7842
rect 22940 7840 23060 7842
rect 19886 7800 19892 7812
rect 19306 7772 19892 7800
rect 19886 7760 19892 7772
rect 19944 7760 19950 7812
rect 20254 7760 20260 7812
rect 20312 7800 20318 7812
rect 21174 7800 21180 7812
rect 20312 7772 20357 7800
rect 21135 7772 21180 7800
rect 20312 7760 20318 7772
rect 21174 7760 21180 7772
rect 21232 7760 21238 7812
rect 21266 7760 21272 7812
rect 21324 7800 21330 7812
rect 21729 7803 21787 7809
rect 21729 7800 21741 7803
rect 21324 7772 21741 7800
rect 21324 7760 21330 7772
rect 21729 7769 21741 7772
rect 21775 7769 21787 7803
rect 21729 7763 21787 7769
rect 21821 7803 21879 7809
rect 21821 7769 21833 7803
rect 21867 7800 21879 7803
rect 22572 7800 22600 7840
rect 21867 7772 22600 7800
rect 21867 7769 21879 7772
rect 21821 7763 21879 7769
rect 22646 7760 22652 7812
rect 22704 7800 22710 7812
rect 22741 7803 22799 7809
rect 22741 7800 22753 7803
rect 22704 7772 22753 7800
rect 22704 7760 22710 7772
rect 22741 7769 22753 7772
rect 22787 7769 22799 7803
rect 23032 7800 23060 7840
rect 23201 7837 23213 7871
rect 23247 7837 23259 7871
rect 23308 7868 23336 7964
rect 24780 7877 24808 8044
rect 26234 7896 26240 7948
rect 26292 7936 26298 7948
rect 29825 7939 29883 7945
rect 29825 7936 29837 7939
rect 26292 7908 29837 7936
rect 26292 7896 26298 7908
rect 29825 7905 29837 7908
rect 29871 7905 29883 7939
rect 37734 7936 37740 7948
rect 37695 7908 37740 7936
rect 29825 7899 29883 7905
rect 37734 7896 37740 7908
rect 37792 7896 37798 7948
rect 23845 7871 23903 7877
rect 23845 7868 23857 7871
rect 23308 7840 23857 7868
rect 23201 7831 23259 7837
rect 23845 7837 23857 7840
rect 23891 7837 23903 7871
rect 23845 7831 23903 7837
rect 24765 7871 24823 7877
rect 24765 7837 24777 7871
rect 24811 7837 24823 7871
rect 24765 7831 24823 7837
rect 29733 7871 29791 7877
rect 29733 7837 29745 7871
rect 29779 7868 29791 7871
rect 30742 7868 30748 7880
rect 29779 7840 30748 7868
rect 29779 7837 29791 7840
rect 29733 7831 29791 7837
rect 30742 7828 30748 7840
rect 30800 7828 30806 7880
rect 37458 7868 37464 7880
rect 37419 7840 37464 7868
rect 37458 7828 37464 7840
rect 37516 7828 37522 7880
rect 24670 7800 24676 7812
rect 23032 7772 24676 7800
rect 22741 7763 22799 7769
rect 24670 7760 24676 7772
rect 24728 7760 24734 7812
rect 22830 7732 22836 7744
rect 18432 7704 22836 7732
rect 14608 7692 14614 7704
rect 22830 7692 22836 7704
rect 22888 7692 22894 7744
rect 22922 7692 22928 7744
rect 22980 7732 22986 7744
rect 23293 7735 23351 7741
rect 23293 7732 23305 7735
rect 22980 7704 23305 7732
rect 22980 7692 22986 7704
rect 23293 7701 23305 7704
rect 23339 7701 23351 7735
rect 23293 7695 23351 7701
rect 23382 7692 23388 7744
rect 23440 7732 23446 7744
rect 23937 7735 23995 7741
rect 23937 7732 23949 7735
rect 23440 7704 23949 7732
rect 23440 7692 23446 7704
rect 23937 7701 23949 7704
rect 23983 7701 23995 7735
rect 24578 7732 24584 7744
rect 24539 7704 24584 7732
rect 23937 7695 23995 7701
rect 24578 7692 24584 7704
rect 24636 7692 24642 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 4525 7531 4583 7537
rect 4525 7497 4537 7531
rect 4571 7528 4583 7531
rect 5074 7528 5080 7540
rect 4571 7500 5080 7528
rect 4571 7497 4583 7500
rect 4525 7491 4583 7497
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 6638 7528 6644 7540
rect 5828 7500 6644 7528
rect 1394 7420 1400 7472
rect 1452 7460 1458 7472
rect 1673 7463 1731 7469
rect 1673 7460 1685 7463
rect 1452 7432 1685 7460
rect 1452 7420 1458 7432
rect 1673 7429 1685 7432
rect 1719 7429 1731 7463
rect 1673 7423 1731 7429
rect 1762 7352 1768 7404
rect 1820 7392 1826 7404
rect 2777 7395 2835 7401
rect 2777 7392 2789 7395
rect 1820 7364 2789 7392
rect 1820 7352 1826 7364
rect 2777 7361 2789 7364
rect 2823 7361 2835 7395
rect 2777 7355 2835 7361
rect 4154 7352 4160 7404
rect 4212 7352 4218 7404
rect 5828 7401 5856 7500
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 8389 7531 8447 7537
rect 8389 7497 8401 7531
rect 8435 7528 8447 7531
rect 9950 7528 9956 7540
rect 8435 7500 9956 7528
rect 8435 7497 8447 7500
rect 8389 7491 8447 7497
rect 9950 7488 9956 7500
rect 10008 7488 10014 7540
rect 17218 7528 17224 7540
rect 11072 7500 17224 7528
rect 5905 7463 5963 7469
rect 5905 7429 5917 7463
rect 5951 7460 5963 7463
rect 9122 7460 9128 7472
rect 5951 7432 7406 7460
rect 9083 7432 9128 7460
rect 5951 7429 5963 7432
rect 5905 7423 5963 7429
rect 9122 7420 9128 7432
rect 9180 7420 9186 7472
rect 10962 7460 10968 7472
rect 10350 7432 10968 7460
rect 10962 7420 10968 7432
rect 11020 7420 11026 7472
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7361 5871 7395
rect 11072 7392 11100 7500
rect 17218 7488 17224 7500
rect 17276 7488 17282 7540
rect 20714 7528 20720 7540
rect 17420 7500 20720 7528
rect 11974 7460 11980 7472
rect 11716 7432 11980 7460
rect 11716 7401 11744 7432
rect 11974 7420 11980 7432
rect 12032 7420 12038 7472
rect 13446 7460 13452 7472
rect 13202 7432 13452 7460
rect 13446 7420 13452 7432
rect 13504 7420 13510 7472
rect 13814 7420 13820 7472
rect 13872 7460 13878 7472
rect 17420 7469 17448 7500
rect 20714 7488 20720 7500
rect 20772 7488 20778 7540
rect 21266 7488 21272 7540
rect 21324 7528 21330 7540
rect 25501 7531 25559 7537
rect 25501 7528 25513 7531
rect 21324 7500 25513 7528
rect 21324 7488 21330 7500
rect 25501 7497 25513 7500
rect 25547 7497 25559 7531
rect 25501 7491 25559 7497
rect 25958 7488 25964 7540
rect 26016 7528 26022 7540
rect 27249 7531 27307 7537
rect 27249 7528 27261 7531
rect 26016 7500 27261 7528
rect 26016 7488 26022 7500
rect 27249 7497 27261 7500
rect 27295 7497 27307 7531
rect 27249 7491 27307 7497
rect 17405 7463 17463 7469
rect 13872 7432 14766 7460
rect 13872 7420 13878 7432
rect 17405 7429 17417 7463
rect 17451 7429 17463 7463
rect 17405 7423 17463 7429
rect 17678 7420 17684 7472
rect 17736 7460 17742 7472
rect 18138 7460 18144 7472
rect 17736 7432 18144 7460
rect 17736 7420 17742 7432
rect 18138 7420 18144 7432
rect 18196 7420 18202 7472
rect 18325 7463 18383 7469
rect 18325 7429 18337 7463
rect 18371 7460 18383 7463
rect 18690 7460 18696 7472
rect 18371 7432 18696 7460
rect 18371 7429 18383 7432
rect 18325 7423 18383 7429
rect 18690 7420 18696 7432
rect 18748 7420 18754 7472
rect 18874 7460 18880 7472
rect 18835 7432 18880 7460
rect 18874 7420 18880 7432
rect 18932 7420 18938 7472
rect 18969 7463 19027 7469
rect 18969 7429 18981 7463
rect 19015 7460 19027 7463
rect 23382 7460 23388 7472
rect 19015 7432 23388 7460
rect 19015 7429 19027 7432
rect 18969 7423 19027 7429
rect 23382 7420 23388 7432
rect 23440 7420 23446 7472
rect 5813 7355 5871 7361
rect 10612 7364 11100 7392
rect 11701 7395 11759 7401
rect 3053 7327 3111 7333
rect 3053 7293 3065 7327
rect 3099 7324 3111 7327
rect 3418 7324 3424 7336
rect 3099 7296 3424 7324
rect 3099 7293 3111 7296
rect 3053 7287 3111 7293
rect 3418 7284 3424 7296
rect 3476 7284 3482 7336
rect 6546 7284 6552 7336
rect 6604 7324 6610 7336
rect 6641 7327 6699 7333
rect 6641 7324 6653 7327
rect 6604 7296 6653 7324
rect 6604 7284 6610 7296
rect 6641 7293 6653 7296
rect 6687 7324 6699 7327
rect 8846 7324 8852 7336
rect 6687 7296 8852 7324
rect 6687 7293 6699 7296
rect 6641 7287 6699 7293
rect 8846 7284 8852 7296
rect 8904 7284 8910 7336
rect 1854 7256 1860 7268
rect 1815 7228 1860 7256
rect 1854 7216 1860 7228
rect 1912 7216 1918 7268
rect 6904 7191 6962 7197
rect 6904 7157 6916 7191
rect 6950 7188 6962 7191
rect 8110 7188 8116 7200
rect 6950 7160 8116 7188
rect 6950 7157 6962 7160
rect 6904 7151 6962 7157
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 8570 7148 8576 7200
rect 8628 7188 8634 7200
rect 10612 7197 10640 7364
rect 11701 7361 11713 7395
rect 11747 7361 11759 7395
rect 20162 7392 20168 7404
rect 11701 7355 11759 7361
rect 19904 7364 20168 7392
rect 11977 7327 12035 7333
rect 11977 7293 11989 7327
rect 12023 7324 12035 7327
rect 12710 7324 12716 7336
rect 12023 7296 12716 7324
rect 12023 7293 12035 7296
rect 11977 7287 12035 7293
rect 12710 7284 12716 7296
rect 12768 7284 12774 7336
rect 12986 7284 12992 7336
rect 13044 7324 13050 7336
rect 13449 7327 13507 7333
rect 13449 7324 13461 7327
rect 13044 7296 13461 7324
rect 13044 7284 13050 7296
rect 13449 7293 13461 7296
rect 13495 7324 13507 7327
rect 13630 7324 13636 7336
rect 13495 7296 13636 7324
rect 13495 7293 13507 7296
rect 13449 7287 13507 7293
rect 13630 7284 13636 7296
rect 13688 7284 13694 7336
rect 13722 7284 13728 7336
rect 13780 7324 13786 7336
rect 14001 7327 14059 7333
rect 14001 7324 14013 7327
rect 13780 7296 14013 7324
rect 13780 7284 13786 7296
rect 14001 7293 14013 7296
rect 14047 7293 14059 7327
rect 14274 7324 14280 7336
rect 14235 7296 14280 7324
rect 14001 7287 14059 7293
rect 14274 7284 14280 7296
rect 14332 7284 14338 7336
rect 15746 7324 15752 7336
rect 15707 7296 15752 7324
rect 15746 7284 15752 7296
rect 15804 7284 15810 7336
rect 17313 7327 17371 7333
rect 17313 7293 17325 7327
rect 17359 7324 17371 7327
rect 17586 7324 17592 7336
rect 17359 7296 17592 7324
rect 17359 7293 17371 7296
rect 17313 7287 17371 7293
rect 17586 7284 17592 7296
rect 17644 7324 17650 7336
rect 19904 7333 19932 7364
rect 20162 7352 20168 7364
rect 20220 7352 20226 7404
rect 20806 7392 20812 7404
rect 20767 7364 20812 7392
rect 20806 7352 20812 7364
rect 20864 7352 20870 7404
rect 20916 7364 21128 7392
rect 19889 7327 19947 7333
rect 19889 7324 19901 7327
rect 17644 7296 19901 7324
rect 17644 7284 17650 7296
rect 19889 7293 19901 7296
rect 19935 7293 19947 7327
rect 20916 7324 20944 7364
rect 19889 7287 19947 7293
rect 19996 7296 20944 7324
rect 20993 7327 21051 7333
rect 15562 7216 15568 7268
rect 15620 7256 15626 7268
rect 17678 7256 17684 7268
rect 15620 7228 17684 7256
rect 15620 7216 15626 7228
rect 17678 7216 17684 7228
rect 17736 7216 17742 7268
rect 19426 7216 19432 7268
rect 19484 7256 19490 7268
rect 19996 7256 20024 7296
rect 20993 7293 21005 7327
rect 21039 7293 21051 7327
rect 21100 7324 21128 7364
rect 21358 7352 21364 7404
rect 21416 7392 21422 7404
rect 22005 7395 22063 7401
rect 22005 7392 22017 7395
rect 21416 7364 22017 7392
rect 21416 7352 21422 7364
rect 22005 7361 22017 7364
rect 22051 7361 22063 7395
rect 22186 7392 22192 7404
rect 22147 7364 22192 7392
rect 22005 7355 22063 7361
rect 22186 7352 22192 7364
rect 22244 7352 22250 7404
rect 23109 7395 23167 7401
rect 23109 7392 23121 7395
rect 22388 7364 23121 7392
rect 22278 7324 22284 7336
rect 21100 7296 22284 7324
rect 20993 7287 21051 7293
rect 19484 7228 20024 7256
rect 19484 7216 19490 7228
rect 10597 7191 10655 7197
rect 10597 7188 10609 7191
rect 8628 7160 10609 7188
rect 8628 7148 8634 7160
rect 10597 7157 10609 7160
rect 10643 7157 10655 7191
rect 10597 7151 10655 7157
rect 16574 7148 16580 7200
rect 16632 7188 16638 7200
rect 18506 7188 18512 7200
rect 16632 7160 18512 7188
rect 16632 7148 16638 7160
rect 18506 7148 18512 7160
rect 18564 7148 18570 7200
rect 19150 7148 19156 7200
rect 19208 7188 19214 7200
rect 20898 7188 20904 7200
rect 19208 7160 20904 7188
rect 19208 7148 19214 7160
rect 20898 7148 20904 7160
rect 20956 7148 20962 7200
rect 21008 7188 21036 7287
rect 22278 7284 22284 7296
rect 22336 7284 22342 7336
rect 22388 7265 22416 7364
rect 23109 7361 23121 7364
rect 23155 7361 23167 7395
rect 23109 7355 23167 7361
rect 23937 7395 23995 7401
rect 23937 7361 23949 7395
rect 23983 7392 23995 7395
rect 24578 7392 24584 7404
rect 23983 7364 24584 7392
rect 23983 7361 23995 7364
rect 23937 7355 23995 7361
rect 24578 7352 24584 7364
rect 24636 7352 24642 7404
rect 25409 7395 25467 7401
rect 25409 7361 25421 7395
rect 25455 7361 25467 7395
rect 27154 7392 27160 7404
rect 27115 7364 27160 7392
rect 25409 7355 25467 7361
rect 22462 7284 22468 7336
rect 22520 7324 22526 7336
rect 23201 7327 23259 7333
rect 23201 7324 23213 7327
rect 22520 7296 23213 7324
rect 22520 7284 22526 7296
rect 23201 7293 23213 7296
rect 23247 7293 23259 7327
rect 25424 7324 25452 7355
rect 27154 7352 27160 7364
rect 27212 7352 27218 7404
rect 30098 7324 30104 7336
rect 25424 7296 30104 7324
rect 23201 7287 23259 7293
rect 30098 7284 30104 7296
rect 30156 7284 30162 7336
rect 21453 7259 21511 7265
rect 21453 7225 21465 7259
rect 21499 7256 21511 7259
rect 22373 7259 22431 7265
rect 22373 7256 22385 7259
rect 21499 7228 22385 7256
rect 21499 7225 21511 7228
rect 21453 7219 21511 7225
rect 22373 7225 22385 7228
rect 22419 7225 22431 7259
rect 23753 7259 23811 7265
rect 23753 7256 23765 7259
rect 22373 7219 22431 7225
rect 22572 7228 23765 7256
rect 22572 7188 22600 7228
rect 23753 7225 23765 7228
rect 23799 7225 23811 7259
rect 23753 7219 23811 7225
rect 21008 7160 22600 7188
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 5524 6987 5582 6993
rect 5524 6953 5536 6987
rect 5570 6984 5582 6987
rect 6822 6984 6828 6996
rect 5570 6956 6828 6984
rect 5570 6953 5582 6956
rect 5524 6947 5582 6953
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 9674 6984 9680 6996
rect 9646 6944 9680 6984
rect 9732 6944 9738 6996
rect 9766 6944 9772 6996
rect 9824 6944 9830 6996
rect 9953 6987 10011 6993
rect 9953 6953 9965 6987
rect 9999 6984 10011 6987
rect 9999 6956 12664 6984
rect 9999 6953 10011 6956
rect 9953 6947 10011 6953
rect 1762 6916 1768 6928
rect 1723 6888 1768 6916
rect 1762 6876 1768 6888
rect 1820 6876 1826 6928
rect 6656 6888 7144 6916
rect 3878 6808 3884 6860
rect 3936 6848 3942 6860
rect 4065 6851 4123 6857
rect 4065 6848 4077 6851
rect 3936 6820 4077 6848
rect 3936 6808 3942 6820
rect 4065 6817 4077 6820
rect 4111 6817 4123 6851
rect 4065 6811 4123 6817
rect 5261 6851 5319 6857
rect 5261 6817 5273 6851
rect 5307 6848 5319 6851
rect 6546 6848 6552 6860
rect 5307 6820 6552 6848
rect 5307 6817 5319 6820
rect 5261 6811 5319 6817
rect 6546 6808 6552 6820
rect 6604 6808 6610 6860
rect 1578 6780 1584 6792
rect 1539 6752 1584 6780
rect 1578 6740 1584 6752
rect 1636 6740 1642 6792
rect 1946 6740 1952 6792
rect 2004 6780 2010 6792
rect 2501 6783 2559 6789
rect 2501 6780 2513 6783
rect 2004 6752 2513 6780
rect 2004 6740 2010 6752
rect 2501 6749 2513 6752
rect 2547 6749 2559 6783
rect 2501 6743 2559 6749
rect 3145 6783 3203 6789
rect 3145 6749 3157 6783
rect 3191 6780 3203 6783
rect 3234 6780 3240 6792
rect 3191 6752 3240 6780
rect 3191 6749 3203 6752
rect 3145 6743 3203 6749
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 3602 6740 3608 6792
rect 3660 6780 3666 6792
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3660 6752 3985 6780
rect 3660 6740 3666 6752
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 6656 6766 6684 6888
rect 6730 6808 6736 6860
rect 6788 6848 6794 6860
rect 7009 6851 7067 6857
rect 7009 6848 7021 6851
rect 6788 6820 7021 6848
rect 6788 6808 6794 6820
rect 7009 6817 7021 6820
rect 7055 6817 7067 6851
rect 7116 6848 7144 6888
rect 8938 6848 8944 6860
rect 7116 6820 8944 6848
rect 7009 6811 7067 6817
rect 3973 6743 4031 6749
rect 7024 6712 7052 6811
rect 8938 6808 8944 6820
rect 8996 6808 9002 6860
rect 9030 6808 9036 6860
rect 9088 6848 9094 6860
rect 9646 6848 9674 6944
rect 9784 6916 9812 6944
rect 12636 6916 12664 6956
rect 12710 6944 12716 6996
rect 12768 6984 12774 6996
rect 12897 6987 12955 6993
rect 12897 6984 12909 6987
rect 12768 6956 12909 6984
rect 12768 6944 12774 6956
rect 12897 6953 12909 6956
rect 12943 6953 12955 6987
rect 13814 6984 13820 6996
rect 12897 6947 12955 6953
rect 13004 6956 13820 6984
rect 13004 6916 13032 6956
rect 13814 6944 13820 6956
rect 13872 6944 13878 6996
rect 14540 6987 14598 6993
rect 14540 6953 14552 6987
rect 14586 6984 14598 6987
rect 15930 6984 15936 6996
rect 14586 6956 15936 6984
rect 14586 6953 14598 6956
rect 14540 6947 14598 6953
rect 15930 6944 15936 6956
rect 15988 6944 15994 6996
rect 16390 6944 16396 6996
rect 16448 6984 16454 6996
rect 22649 6987 22707 6993
rect 22649 6984 22661 6987
rect 16448 6956 22661 6984
rect 16448 6944 16454 6956
rect 22649 6953 22661 6956
rect 22695 6953 22707 6987
rect 22649 6947 22707 6953
rect 9784 6888 11284 6916
rect 12636 6888 13032 6916
rect 9088 6820 9674 6848
rect 9088 6808 9094 6820
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6780 7895 6783
rect 8202 6780 8208 6792
rect 7883 6752 8208 6780
rect 7883 6749 7895 6752
rect 7837 6743 7895 6749
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 9214 6780 9220 6792
rect 9175 6752 9220 6780
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 9306 6740 9312 6792
rect 9364 6780 9370 6792
rect 9674 6780 9680 6792
rect 9364 6752 9409 6780
rect 9364 6740 9370 6752
rect 9646 6740 9680 6780
rect 9732 6740 9738 6792
rect 9853 6777 9911 6783
rect 10060 6780 10088 6888
rect 11146 6848 11152 6860
rect 11107 6820 11152 6848
rect 11146 6808 11152 6820
rect 11204 6808 11210 6860
rect 11256 6848 11284 6888
rect 13262 6876 13268 6928
rect 13320 6916 13326 6928
rect 16025 6919 16083 6925
rect 13320 6888 14044 6916
rect 13320 6876 13326 6888
rect 13449 6851 13507 6857
rect 11256 6820 13400 6848
rect 10502 6780 10508 6792
rect 9853 6743 9865 6777
rect 9899 6774 9911 6777
rect 9955 6774 10088 6780
rect 9899 6752 10088 6774
rect 10463 6752 10508 6780
rect 9899 6746 9983 6752
rect 9899 6743 9911 6746
rect 9646 6712 9674 6740
rect 9853 6737 9911 6743
rect 10502 6740 10508 6752
rect 10560 6740 10566 6792
rect 13170 6780 13176 6792
rect 12558 6752 13176 6780
rect 13170 6740 13176 6752
rect 13228 6740 13234 6792
rect 13372 6789 13400 6820
rect 13449 6817 13461 6851
rect 13495 6848 13507 6851
rect 13538 6848 13544 6860
rect 13495 6820 13544 6848
rect 13495 6817 13507 6820
rect 13449 6811 13507 6817
rect 13538 6808 13544 6820
rect 13596 6808 13602 6860
rect 14016 6848 14044 6888
rect 16025 6885 16037 6919
rect 16071 6916 16083 6919
rect 16482 6916 16488 6928
rect 16071 6888 16488 6916
rect 16071 6885 16083 6888
rect 16025 6879 16083 6885
rect 16482 6876 16488 6888
rect 16540 6876 16546 6928
rect 17129 6919 17187 6925
rect 17129 6885 17141 6919
rect 17175 6916 17187 6919
rect 17175 6888 17908 6916
rect 17175 6885 17187 6888
rect 17129 6879 17187 6885
rect 15562 6848 15568 6860
rect 14016 6820 15568 6848
rect 15562 6808 15568 6820
rect 15620 6808 15626 6860
rect 17770 6848 17776 6860
rect 15672 6820 17264 6848
rect 17731 6820 17776 6848
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6749 13415 6783
rect 13357 6743 13415 6749
rect 13722 6740 13728 6792
rect 13780 6780 13786 6792
rect 14277 6783 14335 6789
rect 14277 6780 14289 6783
rect 13780 6752 14289 6780
rect 13780 6740 13786 6752
rect 14277 6749 14289 6752
rect 14323 6749 14335 6783
rect 15672 6766 15700 6820
rect 14277 6743 14335 6749
rect 7024 6684 9674 6712
rect 10870 6672 10876 6724
rect 10928 6712 10934 6724
rect 11422 6712 11428 6724
rect 10928 6684 11192 6712
rect 11383 6684 11428 6712
rect 10928 6672 10934 6684
rect 2222 6604 2228 6656
rect 2280 6644 2286 6656
rect 2317 6647 2375 6653
rect 2317 6644 2329 6647
rect 2280 6616 2329 6644
rect 2280 6604 2286 6616
rect 2317 6613 2329 6616
rect 2363 6613 2375 6647
rect 2317 6607 2375 6613
rect 2961 6647 3019 6653
rect 2961 6613 2973 6647
rect 3007 6644 3019 6647
rect 6822 6644 6828 6656
rect 3007 6616 6828 6644
rect 3007 6613 3019 6616
rect 2961 6607 3019 6613
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 7650 6644 7656 6656
rect 7611 6616 7656 6644
rect 7650 6604 7656 6616
rect 7708 6604 7714 6656
rect 9674 6604 9680 6656
rect 9732 6644 9738 6656
rect 10410 6644 10416 6656
rect 9732 6616 10416 6644
rect 9732 6604 9738 6616
rect 10410 6604 10416 6616
rect 10468 6604 10474 6656
rect 10597 6647 10655 6653
rect 10597 6613 10609 6647
rect 10643 6644 10655 6647
rect 11054 6644 11060 6656
rect 10643 6616 11060 6644
rect 10643 6613 10655 6616
rect 10597 6607 10655 6613
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 11164 6644 11192 6684
rect 11422 6672 11428 6684
rect 11480 6672 11486 6724
rect 16574 6712 16580 6724
rect 16535 6684 16580 6712
rect 16574 6672 16580 6684
rect 16632 6672 16638 6724
rect 16669 6715 16727 6721
rect 16669 6681 16681 6715
rect 16715 6681 16727 6715
rect 17236 6712 17264 6820
rect 17770 6808 17776 6820
rect 17828 6808 17834 6860
rect 17880 6848 17908 6888
rect 18230 6876 18236 6928
rect 18288 6916 18294 6928
rect 19058 6916 19064 6928
rect 18288 6888 19064 6916
rect 18288 6876 18294 6888
rect 19058 6876 19064 6888
rect 19116 6916 19122 6928
rect 20073 6919 20131 6925
rect 20073 6916 20085 6919
rect 19116 6888 20085 6916
rect 19116 6876 19122 6888
rect 20073 6885 20085 6888
rect 20119 6885 20131 6919
rect 20073 6879 20131 6885
rect 20898 6876 20904 6928
rect 20956 6916 20962 6928
rect 21726 6916 21732 6928
rect 20956 6888 21732 6916
rect 20956 6876 20962 6888
rect 21726 6876 21732 6888
rect 21784 6876 21790 6928
rect 22278 6876 22284 6928
rect 22336 6916 22342 6928
rect 23382 6916 23388 6928
rect 22336 6888 23388 6916
rect 22336 6876 22342 6888
rect 23382 6876 23388 6888
rect 23440 6876 23446 6928
rect 18049 6851 18107 6857
rect 18049 6848 18061 6851
rect 17880 6820 18061 6848
rect 18049 6817 18061 6820
rect 18095 6848 18107 6851
rect 18506 6848 18512 6860
rect 18095 6820 18512 6848
rect 18095 6817 18107 6820
rect 18049 6811 18107 6817
rect 18506 6808 18512 6820
rect 18564 6808 18570 6860
rect 19334 6808 19340 6860
rect 19392 6848 19398 6860
rect 20625 6851 20683 6857
rect 20625 6848 20637 6851
rect 19392 6820 20637 6848
rect 19392 6808 19398 6820
rect 20625 6817 20637 6820
rect 20671 6817 20683 6851
rect 21361 6851 21419 6857
rect 21361 6848 21373 6851
rect 20625 6811 20683 6817
rect 20732 6820 21373 6848
rect 17402 6740 17408 6792
rect 17460 6780 17466 6792
rect 17460 6752 17632 6780
rect 17460 6740 17466 6752
rect 17604 6712 17632 6752
rect 20438 6740 20444 6792
rect 20496 6780 20502 6792
rect 20732 6780 20760 6820
rect 21361 6817 21373 6820
rect 21407 6817 21419 6851
rect 21361 6811 21419 6817
rect 21542 6808 21548 6860
rect 21600 6848 21606 6860
rect 22005 6851 22063 6857
rect 22005 6848 22017 6851
rect 21600 6820 22017 6848
rect 21600 6808 21606 6820
rect 22005 6817 22017 6820
rect 22051 6817 22063 6851
rect 22005 6811 22063 6817
rect 22480 6820 23888 6848
rect 20496 6752 20760 6780
rect 21269 6783 21327 6789
rect 20496 6740 20502 6752
rect 21269 6749 21281 6783
rect 21315 6749 21327 6783
rect 21269 6743 21327 6749
rect 21913 6783 21971 6789
rect 21913 6749 21925 6783
rect 21959 6780 21971 6783
rect 22094 6780 22100 6792
rect 21959 6752 22100 6780
rect 21959 6749 21971 6752
rect 21913 6743 21971 6749
rect 17865 6715 17923 6721
rect 17865 6712 17877 6715
rect 17236 6684 17540 6712
rect 17604 6684 17877 6712
rect 16669 6675 16727 6681
rect 16684 6644 16712 6675
rect 11164 6616 16712 6644
rect 17512 6644 17540 6684
rect 17865 6681 17877 6684
rect 17911 6681 17923 6715
rect 17865 6675 17923 6681
rect 19521 6715 19579 6721
rect 19521 6681 19533 6715
rect 19567 6681 19579 6715
rect 19521 6675 19579 6681
rect 19613 6715 19671 6721
rect 19613 6681 19625 6715
rect 19659 6712 19671 6715
rect 20898 6712 20904 6724
rect 19659 6684 20904 6712
rect 19659 6681 19671 6684
rect 19613 6675 19671 6681
rect 19426 6644 19432 6656
rect 17512 6616 19432 6644
rect 19426 6604 19432 6616
rect 19484 6604 19490 6656
rect 19536 6644 19564 6675
rect 20898 6672 20904 6684
rect 20956 6672 20962 6724
rect 21284 6712 21312 6743
rect 22094 6740 22100 6752
rect 22152 6780 22158 6792
rect 22480 6780 22508 6820
rect 22152 6752 22508 6780
rect 22557 6783 22615 6789
rect 22152 6740 22158 6752
rect 22557 6749 22569 6783
rect 22603 6780 22615 6783
rect 22646 6780 22652 6792
rect 22603 6752 22652 6780
rect 22603 6749 22615 6752
rect 22557 6743 22615 6749
rect 22646 6740 22652 6752
rect 22704 6740 22710 6792
rect 23106 6740 23112 6792
rect 23164 6780 23170 6792
rect 23201 6783 23259 6789
rect 23201 6780 23213 6783
rect 23164 6752 23213 6780
rect 23164 6740 23170 6752
rect 23201 6749 23213 6752
rect 23247 6749 23259 6783
rect 23201 6743 23259 6749
rect 23290 6740 23296 6792
rect 23348 6780 23354 6792
rect 23860 6789 23888 6820
rect 23845 6783 23903 6789
rect 23348 6752 23393 6780
rect 23348 6740 23354 6752
rect 23845 6749 23857 6783
rect 23891 6749 23903 6783
rect 23845 6743 23903 6749
rect 22370 6712 22376 6724
rect 21284 6684 22376 6712
rect 22370 6672 22376 6684
rect 22428 6672 22434 6724
rect 23937 6715 23995 6721
rect 23937 6681 23949 6715
rect 23983 6681 23995 6715
rect 23937 6675 23995 6681
rect 21266 6644 21272 6656
rect 19536 6616 21272 6644
rect 21266 6604 21272 6616
rect 21324 6604 21330 6656
rect 21450 6604 21456 6656
rect 21508 6644 21514 6656
rect 23952 6644 23980 6675
rect 21508 6616 23980 6644
rect 21508 6604 21514 6616
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 1946 6440 1952 6452
rect 1907 6412 1952 6440
rect 1946 6400 1952 6412
rect 2004 6400 2010 6452
rect 4525 6443 4583 6449
rect 4525 6409 4537 6443
rect 4571 6440 4583 6443
rect 4982 6440 4988 6452
rect 4571 6412 4988 6440
rect 4571 6409 4583 6412
rect 4525 6403 4583 6409
rect 4982 6400 4988 6412
rect 5040 6400 5046 6452
rect 7006 6440 7012 6452
rect 5092 6412 7012 6440
rect 5092 6381 5120 6412
rect 7006 6400 7012 6412
rect 7064 6400 7070 6452
rect 8297 6443 8355 6449
rect 8297 6409 8309 6443
rect 8343 6440 8355 6443
rect 8343 6412 10640 6440
rect 8343 6409 8355 6412
rect 8297 6403 8355 6409
rect 5077 6375 5135 6381
rect 5077 6341 5089 6375
rect 5123 6341 5135 6375
rect 6914 6372 6920 6384
rect 5077 6335 5135 6341
rect 6564 6344 6920 6372
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6304 1915 6307
rect 2314 6304 2320 6316
rect 1903 6276 2320 6304
rect 1903 6273 1915 6276
rect 1857 6267 1915 6273
rect 2314 6264 2320 6276
rect 2372 6264 2378 6316
rect 2685 6307 2743 6313
rect 2685 6273 2697 6307
rect 2731 6304 2743 6307
rect 3418 6304 3424 6316
rect 2731 6276 3424 6304
rect 2731 6273 2743 6276
rect 2685 6267 2743 6273
rect 3418 6264 3424 6276
rect 3476 6264 3482 6316
rect 3513 6307 3571 6313
rect 3513 6273 3525 6307
rect 3559 6273 3571 6307
rect 3513 6267 3571 6273
rect 4433 6307 4491 6313
rect 4433 6273 4445 6307
rect 4479 6304 4491 6307
rect 5534 6304 5540 6316
rect 4479 6276 5540 6304
rect 4479 6273 4491 6276
rect 4433 6267 4491 6273
rect 3528 6236 3556 6267
rect 5534 6264 5540 6276
rect 5592 6264 5598 6316
rect 6564 6313 6592 6344
rect 6914 6332 6920 6344
rect 6972 6332 6978 6384
rect 8662 6372 8668 6384
rect 8050 6344 8668 6372
rect 8662 6332 8668 6344
rect 8720 6332 8726 6384
rect 10612 6372 10640 6412
rect 11054 6400 11060 6452
rect 11112 6440 11118 6452
rect 13262 6440 13268 6452
rect 11112 6412 13268 6440
rect 11112 6400 11118 6412
rect 13262 6400 13268 6412
rect 13320 6400 13326 6452
rect 15746 6440 15752 6452
rect 13372 6412 15752 6440
rect 11330 6372 11336 6384
rect 10612 6344 11336 6372
rect 11330 6332 11336 6344
rect 11388 6332 11394 6384
rect 11698 6372 11704 6384
rect 11659 6344 11704 6372
rect 11698 6332 11704 6344
rect 11756 6332 11762 6384
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 9030 6304 9036 6316
rect 8991 6276 9036 6304
rect 6549 6267 6607 6273
rect 9030 6264 9036 6276
rect 9088 6264 9094 6316
rect 4706 6236 4712 6248
rect 3528 6208 4712 6236
rect 4706 6196 4712 6208
rect 4764 6196 4770 6248
rect 5258 6196 5264 6248
rect 5316 6236 5322 6248
rect 5813 6239 5871 6245
rect 5813 6236 5825 6239
rect 5316 6208 5825 6236
rect 5316 6196 5322 6208
rect 5813 6205 5825 6208
rect 5859 6205 5871 6239
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 5813 6199 5871 6205
rect 5920 6208 6837 6236
rect 5534 6128 5540 6180
rect 5592 6168 5598 6180
rect 5920 6168 5948 6208
rect 6825 6205 6837 6208
rect 6871 6205 6883 6239
rect 6825 6199 6883 6205
rect 9309 6239 9367 6245
rect 9309 6205 9321 6239
rect 9355 6236 9367 6239
rect 9858 6236 9864 6248
rect 9355 6208 9864 6236
rect 9355 6205 9367 6208
rect 9309 6199 9367 6205
rect 9858 6196 9864 6208
rect 9916 6196 9922 6248
rect 10428 6236 10456 6290
rect 11146 6264 11152 6316
rect 11204 6304 11210 6316
rect 12437 6307 12495 6313
rect 12437 6304 12449 6307
rect 11204 6276 12449 6304
rect 11204 6264 11210 6276
rect 12437 6273 12449 6276
rect 12483 6273 12495 6307
rect 12437 6267 12495 6273
rect 13372 6236 13400 6412
rect 15746 6400 15752 6412
rect 15804 6400 15810 6452
rect 15856 6412 17908 6440
rect 13722 6372 13728 6384
rect 13464 6344 13728 6372
rect 13464 6248 13492 6344
rect 13722 6332 13728 6344
rect 13780 6332 13786 6384
rect 13814 6332 13820 6384
rect 13872 6372 13878 6384
rect 13872 6344 14214 6372
rect 13872 6332 13878 6344
rect 15856 6313 15884 6412
rect 17126 6372 17132 6384
rect 15948 6344 17132 6372
rect 15841 6307 15899 6313
rect 15304 6276 15792 6304
rect 10428 6208 13400 6236
rect 13446 6196 13452 6248
rect 13504 6236 13510 6248
rect 13725 6239 13783 6245
rect 13504 6208 13549 6236
rect 13504 6196 13510 6208
rect 13725 6205 13737 6239
rect 13771 6236 13783 6239
rect 15194 6236 15200 6248
rect 13771 6208 15200 6236
rect 13771 6205 13783 6208
rect 13725 6199 13783 6205
rect 15194 6196 15200 6208
rect 15252 6196 15258 6248
rect 5592 6140 5948 6168
rect 5592 6128 5598 6140
rect 10318 6128 10324 6180
rect 10376 6168 10382 6180
rect 12250 6168 12256 6180
rect 10376 6140 12256 6168
rect 10376 6128 10382 6140
rect 12250 6128 12256 6140
rect 12308 6128 12314 6180
rect 15304 6168 15332 6276
rect 15654 6236 15660 6248
rect 15615 6208 15660 6236
rect 15654 6196 15660 6208
rect 15712 6196 15718 6248
rect 15764 6236 15792 6276
rect 15841 6273 15853 6307
rect 15887 6273 15899 6307
rect 15841 6267 15899 6273
rect 15948 6236 15976 6344
rect 17126 6332 17132 6344
rect 17184 6332 17190 6384
rect 17770 6372 17776 6384
rect 17731 6344 17776 6372
rect 17770 6332 17776 6344
rect 17828 6332 17834 6384
rect 17880 6372 17908 6412
rect 18046 6400 18052 6452
rect 18104 6440 18110 6452
rect 19794 6440 19800 6452
rect 18104 6412 19800 6440
rect 18104 6400 18110 6412
rect 19794 6400 19800 6412
rect 19852 6400 19858 6452
rect 20346 6400 20352 6452
rect 20404 6440 20410 6452
rect 20404 6412 20449 6440
rect 20404 6400 20410 6412
rect 20898 6400 20904 6452
rect 20956 6440 20962 6452
rect 22738 6440 22744 6452
rect 20956 6412 22744 6440
rect 20956 6400 20962 6412
rect 22738 6400 22744 6412
rect 22796 6400 22802 6452
rect 38105 6443 38163 6449
rect 38105 6440 38117 6443
rect 35866 6412 38117 6440
rect 20993 6375 21051 6381
rect 20993 6372 21005 6375
rect 17880 6344 21005 6372
rect 20993 6341 21005 6344
rect 21039 6341 21051 6375
rect 20993 6335 21051 6341
rect 21082 6332 21088 6384
rect 21140 6372 21146 6384
rect 22649 6375 22707 6381
rect 22649 6372 22661 6375
rect 21140 6344 22661 6372
rect 21140 6332 21146 6344
rect 22649 6341 22661 6344
rect 22695 6341 22707 6375
rect 22649 6335 22707 6341
rect 16853 6307 16911 6313
rect 16853 6273 16865 6307
rect 16899 6304 16911 6307
rect 17310 6304 17316 6316
rect 16899 6276 17316 6304
rect 16899 6273 16911 6276
rect 16853 6267 16911 6273
rect 17310 6264 17316 6276
rect 17368 6264 17374 6316
rect 19153 6307 19211 6313
rect 19153 6273 19165 6307
rect 19199 6304 19211 6307
rect 20162 6304 20168 6316
rect 19199 6276 20168 6304
rect 19199 6273 19211 6276
rect 19153 6267 19211 6273
rect 20162 6264 20168 6276
rect 20220 6264 20226 6316
rect 20257 6307 20315 6313
rect 20257 6273 20269 6307
rect 20303 6304 20315 6307
rect 20622 6304 20628 6316
rect 20303 6276 20628 6304
rect 20303 6273 20315 6276
rect 20257 6267 20315 6273
rect 20622 6264 20628 6276
rect 20680 6264 20686 6316
rect 20898 6304 20904 6316
rect 20859 6276 20904 6304
rect 20898 6264 20904 6276
rect 20956 6304 20962 6316
rect 30561 6307 30619 6313
rect 20956 6276 22094 6304
rect 20956 6264 20962 6276
rect 15764 6208 15976 6236
rect 17681 6239 17739 6245
rect 17681 6205 17693 6239
rect 17727 6205 17739 6239
rect 18138 6236 18144 6248
rect 18099 6208 18144 6236
rect 17681 6199 17739 6205
rect 14752 6140 15332 6168
rect 2498 6100 2504 6112
rect 2459 6072 2504 6100
rect 2498 6060 2504 6072
rect 2556 6060 2562 6112
rect 3050 6060 3056 6112
rect 3108 6100 3114 6112
rect 3329 6103 3387 6109
rect 3329 6100 3341 6103
rect 3108 6072 3341 6100
rect 3108 6060 3114 6072
rect 3329 6069 3341 6072
rect 3375 6069 3387 6103
rect 3329 6063 3387 6069
rect 5626 6060 5632 6112
rect 5684 6100 5690 6112
rect 8386 6100 8392 6112
rect 5684 6072 8392 6100
rect 5684 6060 5690 6072
rect 8386 6060 8392 6072
rect 8444 6060 8450 6112
rect 8662 6100 8668 6112
rect 8623 6072 8668 6100
rect 8662 6060 8668 6072
rect 8720 6060 8726 6112
rect 10042 6060 10048 6112
rect 10100 6100 10106 6112
rect 10781 6103 10839 6109
rect 10781 6100 10793 6103
rect 10100 6072 10793 6100
rect 10100 6060 10106 6072
rect 10781 6069 10793 6072
rect 10827 6069 10839 6103
rect 10781 6063 10839 6069
rect 12434 6060 12440 6112
rect 12492 6100 12498 6112
rect 14752 6100 14780 6140
rect 15378 6128 15384 6180
rect 15436 6168 15442 6180
rect 17402 6168 17408 6180
rect 15436 6140 17408 6168
rect 15436 6128 15442 6140
rect 17402 6128 17408 6140
rect 17460 6128 17466 6180
rect 17696 6168 17724 6199
rect 18138 6196 18144 6208
rect 18196 6196 18202 6248
rect 19337 6239 19395 6245
rect 19337 6205 19349 6239
rect 19383 6236 19395 6239
rect 21082 6236 21088 6248
rect 19383 6208 21088 6236
rect 19383 6205 19395 6208
rect 19337 6199 19395 6205
rect 21082 6196 21088 6208
rect 21140 6196 21146 6248
rect 22066 6236 22094 6276
rect 30561 6273 30573 6307
rect 30607 6304 30619 6307
rect 35866 6304 35894 6412
rect 38105 6409 38117 6412
rect 38151 6409 38163 6443
rect 38105 6403 38163 6409
rect 38286 6304 38292 6316
rect 30607 6276 35894 6304
rect 38247 6276 38292 6304
rect 30607 6273 30619 6276
rect 30561 6267 30619 6273
rect 38286 6264 38292 6276
rect 38344 6264 38350 6316
rect 22557 6239 22615 6245
rect 22066 6208 22508 6236
rect 20622 6168 20628 6180
rect 17696 6140 20628 6168
rect 20622 6128 20628 6140
rect 20680 6128 20686 6180
rect 22480 6168 22508 6208
rect 22557 6205 22569 6239
rect 22603 6236 22615 6239
rect 23014 6236 23020 6248
rect 22603 6208 23020 6236
rect 22603 6205 22615 6208
rect 22557 6199 22615 6205
rect 23014 6196 23020 6208
rect 23072 6196 23078 6248
rect 23198 6236 23204 6248
rect 23159 6208 23204 6236
rect 23198 6196 23204 6208
rect 23256 6196 23262 6248
rect 23106 6168 23112 6180
rect 22480 6140 23112 6168
rect 23106 6128 23112 6140
rect 23164 6128 23170 6180
rect 30650 6168 30656 6180
rect 30611 6140 30656 6168
rect 30650 6128 30656 6140
rect 30708 6128 30714 6180
rect 12492 6072 14780 6100
rect 15197 6103 15255 6109
rect 12492 6060 12498 6072
rect 15197 6069 15209 6103
rect 15243 6100 15255 6103
rect 15930 6100 15936 6112
rect 15243 6072 15936 6100
rect 15243 6069 15255 6072
rect 15197 6063 15255 6069
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 16298 6100 16304 6112
rect 16259 6072 16304 6100
rect 16298 6060 16304 6072
rect 16356 6060 16362 6112
rect 16945 6103 17003 6109
rect 16945 6069 16957 6103
rect 16991 6100 17003 6103
rect 18598 6100 18604 6112
rect 16991 6072 18604 6100
rect 16991 6069 17003 6072
rect 16945 6063 17003 6069
rect 18598 6060 18604 6072
rect 18656 6060 18662 6112
rect 19518 6100 19524 6112
rect 19479 6072 19524 6100
rect 19518 6060 19524 6072
rect 19576 6060 19582 6112
rect 19794 6060 19800 6112
rect 19852 6100 19858 6112
rect 20898 6100 20904 6112
rect 19852 6072 20904 6100
rect 19852 6060 19858 6072
rect 20898 6060 20904 6072
rect 20956 6060 20962 6112
rect 21082 6060 21088 6112
rect 21140 6100 21146 6112
rect 22922 6100 22928 6112
rect 21140 6072 22928 6100
rect 21140 6060 21146 6072
rect 22922 6060 22928 6072
rect 22980 6060 22986 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 1578 5856 1584 5908
rect 1636 5896 1642 5908
rect 3329 5899 3387 5905
rect 3329 5896 3341 5899
rect 1636 5868 3341 5896
rect 1636 5856 1642 5868
rect 3329 5865 3341 5868
rect 3375 5896 3387 5899
rect 6914 5896 6920 5908
rect 3375 5868 6920 5896
rect 3375 5865 3387 5868
rect 3329 5859 3387 5865
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 7282 5856 7288 5908
rect 7340 5896 7346 5908
rect 10318 5896 10324 5908
rect 7340 5868 10324 5896
rect 7340 5856 7346 5868
rect 10318 5856 10324 5868
rect 10376 5856 10382 5908
rect 11057 5899 11115 5905
rect 11057 5865 11069 5899
rect 11103 5896 11115 5899
rect 11780 5899 11838 5905
rect 11780 5896 11792 5899
rect 11103 5868 11792 5896
rect 11103 5865 11115 5868
rect 11057 5859 11115 5865
rect 11780 5865 11792 5868
rect 11826 5896 11838 5899
rect 12434 5896 12440 5908
rect 11826 5868 12440 5896
rect 11826 5865 11838 5868
rect 11780 5859 11838 5865
rect 12434 5856 12440 5868
rect 12492 5856 12498 5908
rect 16298 5856 16304 5908
rect 16356 5896 16362 5908
rect 18417 5899 18475 5905
rect 18417 5896 18429 5899
rect 16356 5868 18429 5896
rect 16356 5856 16362 5868
rect 18417 5865 18429 5868
rect 18463 5896 18475 5899
rect 19518 5896 19524 5908
rect 18463 5868 19524 5896
rect 18463 5865 18475 5868
rect 18417 5859 18475 5865
rect 19518 5856 19524 5868
rect 19576 5856 19582 5908
rect 19610 5856 19616 5908
rect 19668 5896 19674 5908
rect 19668 5868 20024 5896
rect 19668 5856 19674 5868
rect 3973 5831 4031 5837
rect 3973 5797 3985 5831
rect 4019 5828 4031 5831
rect 4062 5828 4068 5840
rect 4019 5800 4068 5828
rect 4019 5797 4031 5800
rect 3973 5791 4031 5797
rect 4062 5788 4068 5800
rect 4120 5788 4126 5840
rect 7837 5831 7895 5837
rect 4172 5800 5396 5828
rect 1857 5763 1915 5769
rect 1857 5729 1869 5763
rect 1903 5760 1915 5763
rect 4172 5760 4200 5800
rect 5258 5760 5264 5772
rect 1903 5732 4200 5760
rect 4724 5732 5120 5760
rect 5219 5732 5264 5760
rect 1903 5729 1915 5732
rect 1857 5723 1915 5729
rect 1578 5692 1584 5704
rect 1539 5664 1584 5692
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 4157 5695 4215 5701
rect 4157 5661 4169 5695
rect 4203 5692 4215 5695
rect 4724 5692 4752 5732
rect 4203 5664 4752 5692
rect 4801 5695 4859 5701
rect 4203 5661 4215 5664
rect 4157 5655 4215 5661
rect 4801 5661 4813 5695
rect 4847 5661 4859 5695
rect 4801 5655 4859 5661
rect 2866 5584 2872 5636
rect 2924 5584 2930 5636
rect 3786 5584 3792 5636
rect 3844 5624 3850 5636
rect 4816 5624 4844 5655
rect 3844 5596 4844 5624
rect 3844 5584 3850 5596
rect 4617 5559 4675 5565
rect 4617 5525 4629 5559
rect 4663 5556 4675 5559
rect 4890 5556 4896 5568
rect 4663 5528 4896 5556
rect 4663 5525 4675 5528
rect 4617 5519 4675 5525
rect 4890 5516 4896 5528
rect 4948 5516 4954 5568
rect 5092 5556 5120 5732
rect 5258 5720 5264 5732
rect 5316 5720 5322 5772
rect 5368 5760 5396 5800
rect 7837 5797 7849 5831
rect 7883 5828 7895 5831
rect 7883 5800 8800 5828
rect 7883 5797 7895 5800
rect 7837 5791 7895 5797
rect 6546 5760 6552 5772
rect 5368 5732 6552 5760
rect 6546 5720 6552 5732
rect 6604 5720 6610 5772
rect 8478 5760 8484 5772
rect 6656 5732 8484 5760
rect 6656 5678 6684 5732
rect 8478 5720 8484 5732
rect 8536 5720 8542 5772
rect 6822 5652 6828 5704
rect 6880 5692 6886 5704
rect 7745 5695 7803 5701
rect 7745 5692 7757 5695
rect 6880 5664 7757 5692
rect 6880 5652 6886 5664
rect 7745 5661 7757 5664
rect 7791 5661 7803 5695
rect 8386 5692 8392 5704
rect 8347 5664 8392 5692
rect 7745 5655 7803 5661
rect 8386 5652 8392 5664
rect 8444 5652 8450 5704
rect 8772 5692 8800 5800
rect 18156 5800 18460 5828
rect 8846 5720 8852 5772
rect 8904 5760 8910 5772
rect 9309 5763 9367 5769
rect 9309 5760 9321 5763
rect 8904 5732 9321 5760
rect 8904 5720 8910 5732
rect 9309 5729 9321 5732
rect 9355 5729 9367 5763
rect 9309 5723 9367 5729
rect 9585 5763 9643 5769
rect 9585 5729 9597 5763
rect 9631 5760 9643 5763
rect 11517 5763 11575 5769
rect 9631 5732 11192 5760
rect 9631 5729 9643 5732
rect 9585 5723 9643 5729
rect 8772 5664 9168 5692
rect 5537 5627 5595 5633
rect 5537 5593 5549 5627
rect 5583 5624 5595 5627
rect 5626 5624 5632 5636
rect 5583 5596 5632 5624
rect 5583 5593 5595 5596
rect 5537 5587 5595 5593
rect 5626 5584 5632 5596
rect 5684 5584 5690 5636
rect 7282 5624 7288 5636
rect 7243 5596 7288 5624
rect 7282 5584 7288 5596
rect 7340 5584 7346 5636
rect 9030 5624 9036 5636
rect 8404 5596 9036 5624
rect 8404 5556 8432 5596
rect 9030 5584 9036 5596
rect 9088 5584 9094 5636
rect 9140 5624 9168 5664
rect 9674 5624 9680 5636
rect 9140 5596 9680 5624
rect 9674 5584 9680 5596
rect 9732 5584 9738 5636
rect 10594 5584 10600 5636
rect 10652 5584 10658 5636
rect 5092 5528 8432 5556
rect 8481 5559 8539 5565
rect 8481 5525 8493 5559
rect 8527 5556 8539 5559
rect 11054 5556 11060 5568
rect 8527 5528 11060 5556
rect 8527 5525 8539 5528
rect 8481 5519 8539 5525
rect 11054 5516 11060 5528
rect 11112 5516 11118 5568
rect 11164 5556 11192 5732
rect 11517 5729 11529 5763
rect 11563 5760 11575 5763
rect 13446 5760 13452 5772
rect 11563 5732 13452 5760
rect 11563 5729 11575 5732
rect 11517 5723 11575 5729
rect 13446 5720 13452 5732
rect 13504 5720 13510 5772
rect 16022 5760 16028 5772
rect 14200 5732 16028 5760
rect 14200 5692 14228 5732
rect 16022 5720 16028 5732
rect 16080 5720 16086 5772
rect 16577 5763 16635 5769
rect 16577 5729 16589 5763
rect 16623 5760 16635 5763
rect 17402 5760 17408 5772
rect 16623 5732 17408 5760
rect 16623 5729 16635 5732
rect 16577 5723 16635 5729
rect 17402 5720 17408 5732
rect 17460 5720 17466 5772
rect 17586 5760 17592 5772
rect 17547 5732 17592 5760
rect 17586 5720 17592 5732
rect 17644 5720 17650 5772
rect 18156 5760 18184 5800
rect 17972 5732 18184 5760
rect 18432 5760 18460 5800
rect 19242 5788 19248 5840
rect 19300 5828 19306 5840
rect 19996 5828 20024 5868
rect 20254 5856 20260 5908
rect 20312 5896 20318 5908
rect 20441 5899 20499 5905
rect 20441 5896 20453 5899
rect 20312 5868 20453 5896
rect 20312 5856 20318 5868
rect 20441 5865 20453 5868
rect 20487 5865 20499 5899
rect 20441 5859 20499 5865
rect 20622 5856 20628 5908
rect 20680 5896 20686 5908
rect 22278 5896 22284 5908
rect 20680 5868 22284 5896
rect 20680 5856 20686 5868
rect 22278 5856 22284 5868
rect 22336 5856 22342 5908
rect 22370 5856 22376 5908
rect 22428 5896 22434 5908
rect 24486 5896 24492 5908
rect 22428 5868 24492 5896
rect 22428 5856 22434 5868
rect 24486 5856 24492 5868
rect 24544 5856 24550 5908
rect 23661 5831 23719 5837
rect 23661 5828 23673 5831
rect 19300 5800 19932 5828
rect 19996 5800 23673 5828
rect 19300 5788 19306 5800
rect 18432 5732 19840 5760
rect 13096 5664 14228 5692
rect 14277 5695 14335 5701
rect 12250 5584 12256 5636
rect 12308 5584 12314 5636
rect 13096 5556 13124 5664
rect 14277 5661 14289 5695
rect 14323 5661 14335 5695
rect 14277 5655 14335 5661
rect 13446 5584 13452 5636
rect 13504 5624 13510 5636
rect 14292 5624 14320 5655
rect 15654 5652 15660 5704
rect 15712 5652 15718 5704
rect 14550 5624 14556 5636
rect 13504 5596 14320 5624
rect 14511 5596 14556 5624
rect 13504 5584 13510 5596
rect 14550 5584 14556 5596
rect 14608 5584 14614 5636
rect 16669 5627 16727 5633
rect 16669 5593 16681 5627
rect 16715 5624 16727 5627
rect 17972 5624 18000 5732
rect 18049 5695 18107 5701
rect 18049 5661 18061 5695
rect 18095 5661 18107 5695
rect 18049 5655 18107 5661
rect 18233 5695 18291 5701
rect 18233 5661 18245 5695
rect 18279 5692 18291 5695
rect 19429 5695 19487 5701
rect 18279 5664 19380 5692
rect 18279 5661 18291 5664
rect 18233 5655 18291 5661
rect 16715 5596 18000 5624
rect 18064 5624 18092 5655
rect 19150 5624 19156 5636
rect 18064 5596 19156 5624
rect 16715 5593 16727 5596
rect 16669 5587 16727 5593
rect 19150 5584 19156 5596
rect 19208 5584 19214 5636
rect 13262 5556 13268 5568
rect 11164 5528 13124 5556
rect 13223 5528 13268 5556
rect 13262 5516 13268 5528
rect 13320 5516 13326 5568
rect 14090 5516 14096 5568
rect 14148 5556 14154 5568
rect 16025 5559 16083 5565
rect 16025 5556 16037 5559
rect 14148 5528 16037 5556
rect 14148 5516 14154 5528
rect 16025 5525 16037 5528
rect 16071 5556 16083 5559
rect 19058 5556 19064 5568
rect 16071 5528 19064 5556
rect 16071 5525 16083 5528
rect 16025 5519 16083 5525
rect 19058 5516 19064 5528
rect 19116 5516 19122 5568
rect 19352 5556 19380 5664
rect 19429 5661 19441 5695
rect 19475 5692 19487 5695
rect 19610 5692 19616 5704
rect 19475 5664 19616 5692
rect 19475 5661 19487 5664
rect 19429 5655 19487 5661
rect 19610 5652 19616 5664
rect 19668 5652 19674 5704
rect 19702 5624 19708 5636
rect 19663 5596 19708 5624
rect 19702 5584 19708 5596
rect 19760 5584 19766 5636
rect 19812 5624 19840 5732
rect 19904 5692 19932 5800
rect 23661 5797 23673 5800
rect 23707 5797 23719 5831
rect 23661 5791 23719 5797
rect 20254 5720 20260 5772
rect 20312 5760 20318 5772
rect 21729 5763 21787 5769
rect 21729 5760 21741 5763
rect 20312 5732 21741 5760
rect 20312 5720 20318 5732
rect 21729 5729 21741 5732
rect 21775 5729 21787 5763
rect 22278 5760 22284 5772
rect 22239 5732 22284 5760
rect 21729 5723 21787 5729
rect 22278 5720 22284 5732
rect 22336 5720 22342 5772
rect 22646 5720 22652 5772
rect 22704 5760 22710 5772
rect 22704 5732 23152 5760
rect 22704 5720 22710 5732
rect 20349 5695 20407 5701
rect 20349 5692 20361 5695
rect 19904 5664 20361 5692
rect 20349 5661 20361 5664
rect 20395 5661 20407 5695
rect 20349 5655 20407 5661
rect 20806 5652 20812 5704
rect 20864 5692 20870 5704
rect 20993 5695 21051 5701
rect 20993 5692 21005 5695
rect 20864 5664 21005 5692
rect 20864 5652 20870 5664
rect 20993 5661 21005 5664
rect 21039 5692 21051 5695
rect 21266 5692 21272 5704
rect 21039 5664 21272 5692
rect 21039 5661 21051 5664
rect 20993 5655 21051 5661
rect 21266 5652 21272 5664
rect 21324 5652 21330 5704
rect 21358 5652 21364 5704
rect 21416 5692 21422 5704
rect 21637 5695 21695 5701
rect 21637 5692 21649 5695
rect 21416 5664 21649 5692
rect 21416 5652 21422 5664
rect 21637 5661 21649 5664
rect 21683 5661 21695 5695
rect 21637 5655 21695 5661
rect 21818 5652 21824 5704
rect 21876 5692 21882 5704
rect 22925 5695 22983 5701
rect 22925 5692 22937 5695
rect 21876 5664 22937 5692
rect 21876 5652 21882 5664
rect 22925 5661 22937 5664
rect 22971 5661 22983 5695
rect 23124 5692 23152 5732
rect 23198 5720 23204 5772
rect 23256 5760 23262 5772
rect 23256 5732 25728 5760
rect 23256 5720 23262 5732
rect 25700 5701 25728 5732
rect 23569 5695 23627 5701
rect 23569 5692 23581 5695
rect 23124 5664 23581 5692
rect 22925 5655 22983 5661
rect 23569 5661 23581 5664
rect 23615 5661 23627 5695
rect 23569 5655 23627 5661
rect 25685 5695 25743 5701
rect 25685 5661 25697 5695
rect 25731 5661 25743 5695
rect 25685 5655 25743 5661
rect 23017 5627 23075 5633
rect 23017 5624 23029 5627
rect 19812 5596 23029 5624
rect 23017 5593 23029 5596
rect 23063 5593 23075 5627
rect 23017 5587 23075 5593
rect 21085 5559 21143 5565
rect 21085 5556 21097 5559
rect 19352 5528 21097 5556
rect 21085 5525 21097 5528
rect 21131 5525 21143 5559
rect 21085 5519 21143 5525
rect 21174 5516 21180 5568
rect 21232 5556 21238 5568
rect 25222 5556 25228 5568
rect 21232 5528 25228 5556
rect 21232 5516 21238 5528
rect 25222 5516 25228 5528
rect 25280 5516 25286 5568
rect 25777 5559 25835 5565
rect 25777 5525 25789 5559
rect 25823 5556 25835 5559
rect 26418 5556 26424 5568
rect 25823 5528 26424 5556
rect 25823 5525 25835 5528
rect 25777 5519 25835 5525
rect 26418 5516 26424 5528
rect 26476 5516 26482 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 3421 5355 3479 5361
rect 3421 5321 3433 5355
rect 3467 5352 3479 5355
rect 3510 5352 3516 5364
rect 3467 5324 3516 5352
rect 3467 5321 3479 5324
rect 3421 5315 3479 5321
rect 3510 5312 3516 5324
rect 3568 5312 3574 5364
rect 4614 5312 4620 5364
rect 4672 5312 4678 5364
rect 11054 5312 11060 5364
rect 11112 5352 11118 5364
rect 19978 5352 19984 5364
rect 11112 5324 15976 5352
rect 11112 5312 11118 5324
rect 4632 5284 4660 5312
rect 2746 5256 4660 5284
rect 6917 5287 6975 5293
rect 1394 5176 1400 5228
rect 1452 5216 1458 5228
rect 1581 5219 1639 5225
rect 1581 5216 1593 5219
rect 1452 5188 1593 5216
rect 1452 5176 1458 5188
rect 1581 5185 1593 5188
rect 1627 5185 1639 5219
rect 1581 5179 1639 5185
rect 1857 5151 1915 5157
rect 1857 5117 1869 5151
rect 1903 5117 1915 5151
rect 1857 5111 1915 5117
rect 1872 5012 1900 5111
rect 2746 5012 2774 5256
rect 6917 5253 6929 5287
rect 6963 5284 6975 5287
rect 7006 5284 7012 5296
rect 6963 5256 7012 5284
rect 6963 5253 6975 5256
rect 6917 5247 6975 5253
rect 7006 5244 7012 5256
rect 7064 5244 7070 5296
rect 7745 5287 7803 5293
rect 7745 5253 7757 5287
rect 7791 5284 7803 5287
rect 8846 5284 8852 5296
rect 7791 5256 8852 5284
rect 7791 5253 7803 5256
rect 7745 5247 7803 5253
rect 8312 5228 8340 5256
rect 8846 5244 8852 5256
rect 8904 5244 8910 5296
rect 11698 5244 11704 5296
rect 11756 5284 11762 5296
rect 12069 5287 12127 5293
rect 12069 5284 12081 5287
rect 11756 5256 12081 5284
rect 11756 5244 11762 5256
rect 12069 5253 12081 5256
rect 12115 5253 12127 5287
rect 12069 5247 12127 5253
rect 12897 5287 12955 5293
rect 12897 5253 12909 5287
rect 12943 5284 12955 5287
rect 13354 5284 13360 5296
rect 12943 5256 13360 5284
rect 12943 5253 12955 5256
rect 12897 5247 12955 5253
rect 13354 5244 13360 5256
rect 13412 5284 13418 5296
rect 13722 5284 13728 5296
rect 13412 5256 13728 5284
rect 13412 5244 13418 5256
rect 13722 5244 13728 5256
rect 13780 5244 13786 5296
rect 15746 5284 15752 5296
rect 14950 5256 15752 5284
rect 15746 5244 15752 5256
rect 15804 5244 15810 5296
rect 3329 5219 3387 5225
rect 3329 5185 3341 5219
rect 3375 5216 3387 5219
rect 3602 5216 3608 5228
rect 3375 5188 3608 5216
rect 3375 5185 3387 5188
rect 3329 5179 3387 5185
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 8294 5216 8300 5228
rect 5382 5188 7880 5216
rect 8207 5188 8300 5216
rect 3973 5151 4031 5157
rect 3973 5117 3985 5151
rect 4019 5117 4031 5151
rect 3973 5111 4031 5117
rect 4249 5151 4307 5157
rect 4249 5117 4261 5151
rect 4295 5148 4307 5151
rect 6730 5148 6736 5160
rect 4295 5120 6736 5148
rect 4295 5117 4307 5120
rect 4249 5111 4307 5117
rect 3326 5040 3332 5092
rect 3384 5080 3390 5092
rect 3988 5080 4016 5111
rect 6730 5108 6736 5120
rect 6788 5108 6794 5160
rect 3384 5052 4016 5080
rect 3384 5040 3390 5052
rect 1872 4984 2774 5012
rect 3988 5012 4016 5052
rect 5258 5012 5264 5024
rect 3988 4984 5264 5012
rect 5258 4972 5264 4984
rect 5316 4972 5322 5024
rect 5534 4972 5540 5024
rect 5592 5012 5598 5024
rect 5721 5015 5779 5021
rect 5721 5012 5733 5015
rect 5592 4984 5733 5012
rect 5592 4972 5598 4984
rect 5721 4981 5733 4984
rect 5767 4981 5779 5015
rect 7852 5012 7880 5188
rect 8294 5176 8300 5188
rect 8352 5176 8358 5228
rect 8570 5148 8576 5160
rect 8531 5120 8576 5148
rect 8570 5108 8576 5120
rect 8628 5108 8634 5160
rect 9692 5080 9720 5202
rect 9858 5176 9864 5228
rect 9916 5216 9922 5228
rect 10318 5216 10324 5228
rect 9916 5188 10324 5216
rect 9916 5176 9922 5188
rect 10318 5176 10324 5188
rect 10376 5176 10382 5228
rect 10962 5216 10968 5228
rect 10923 5188 10968 5216
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 11146 5176 11152 5228
rect 11204 5216 11210 5228
rect 13449 5219 13507 5225
rect 13449 5216 13461 5219
rect 11204 5188 13461 5216
rect 11204 5176 11210 5188
rect 13449 5185 13461 5188
rect 13495 5185 13507 5219
rect 13449 5179 13507 5185
rect 15841 5219 15899 5225
rect 15841 5185 15853 5219
rect 15887 5216 15899 5219
rect 15948 5216 15976 5324
rect 16960 5324 19984 5352
rect 16960 5293 16988 5324
rect 19978 5312 19984 5324
rect 20036 5312 20042 5364
rect 20162 5312 20168 5364
rect 20220 5352 20226 5364
rect 22278 5352 22284 5364
rect 20220 5324 22284 5352
rect 20220 5312 20226 5324
rect 22278 5312 22284 5324
rect 22336 5312 22342 5364
rect 22370 5312 22376 5364
rect 22428 5352 22434 5364
rect 23845 5355 23903 5361
rect 23845 5352 23857 5355
rect 22428 5324 23857 5352
rect 22428 5312 22434 5324
rect 23845 5321 23857 5324
rect 23891 5321 23903 5355
rect 23845 5315 23903 5321
rect 16945 5287 17003 5293
rect 16945 5253 16957 5287
rect 16991 5253 17003 5287
rect 16945 5247 17003 5253
rect 17034 5244 17040 5296
rect 17092 5284 17098 5296
rect 17092 5256 17137 5284
rect 17092 5244 17098 5256
rect 17218 5244 17224 5296
rect 17276 5284 17282 5296
rect 17276 5256 17908 5284
rect 17276 5244 17282 5256
rect 15887 5188 15976 5216
rect 17880 5216 17908 5256
rect 17954 5244 17960 5296
rect 18012 5284 18018 5296
rect 18509 5287 18567 5293
rect 18509 5284 18521 5287
rect 18012 5256 18521 5284
rect 18012 5244 18018 5256
rect 18509 5253 18521 5256
rect 18555 5253 18567 5287
rect 18509 5247 18567 5253
rect 18601 5287 18659 5293
rect 18601 5253 18613 5287
rect 18647 5284 18659 5287
rect 19334 5284 19340 5296
rect 18647 5256 19340 5284
rect 18647 5253 18659 5256
rect 18601 5247 18659 5253
rect 19334 5244 19340 5256
rect 19392 5244 19398 5296
rect 19518 5244 19524 5296
rect 19576 5284 19582 5296
rect 20073 5287 20131 5293
rect 20073 5284 20085 5287
rect 19576 5256 20085 5284
rect 19576 5244 19582 5256
rect 20073 5253 20085 5256
rect 20119 5253 20131 5287
rect 20073 5247 20131 5253
rect 20254 5244 20260 5296
rect 20312 5284 20318 5296
rect 21542 5284 21548 5296
rect 20312 5256 21548 5284
rect 20312 5244 20318 5256
rect 21542 5244 21548 5256
rect 21600 5244 21606 5296
rect 21634 5244 21640 5296
rect 21692 5284 21698 5296
rect 22097 5287 22155 5293
rect 22097 5284 22109 5287
rect 21692 5256 22109 5284
rect 21692 5244 21698 5256
rect 22097 5253 22109 5256
rect 22143 5253 22155 5287
rect 22097 5247 22155 5253
rect 22186 5244 22192 5296
rect 22244 5284 22250 5296
rect 22244 5256 22289 5284
rect 22244 5244 22250 5256
rect 22554 5244 22560 5296
rect 22612 5284 22618 5296
rect 22612 5256 23244 5284
rect 22612 5244 22618 5256
rect 18230 5216 18236 5228
rect 17880 5188 18236 5216
rect 15887 5185 15899 5188
rect 15841 5179 15899 5185
rect 18230 5176 18236 5188
rect 18288 5176 18294 5228
rect 19150 5176 19156 5228
rect 19208 5216 19214 5228
rect 19702 5216 19708 5228
rect 19208 5188 19708 5216
rect 19208 5176 19214 5188
rect 19702 5176 19708 5188
rect 19760 5176 19766 5228
rect 21082 5216 21088 5228
rect 21043 5188 21088 5216
rect 21082 5176 21088 5188
rect 21140 5176 21146 5228
rect 22741 5219 22799 5225
rect 22741 5185 22753 5219
rect 22787 5216 22799 5219
rect 23106 5216 23112 5228
rect 22787 5188 23112 5216
rect 22787 5185 22799 5188
rect 22741 5179 22799 5185
rect 10045 5151 10103 5157
rect 10045 5117 10057 5151
rect 10091 5148 10103 5151
rect 12158 5148 12164 5160
rect 10091 5120 12164 5148
rect 10091 5117 10103 5120
rect 10045 5111 10103 5117
rect 12158 5108 12164 5120
rect 12216 5108 12222 5160
rect 13725 5151 13783 5157
rect 13725 5117 13737 5151
rect 13771 5148 13783 5151
rect 14090 5148 14096 5160
rect 13771 5120 14096 5148
rect 13771 5117 13783 5120
rect 13725 5111 13783 5117
rect 14090 5108 14096 5120
rect 14148 5108 14154 5160
rect 14182 5108 14188 5160
rect 14240 5148 14246 5160
rect 15470 5148 15476 5160
rect 14240 5120 15476 5148
rect 14240 5108 14246 5120
rect 15470 5108 15476 5120
rect 15528 5108 15534 5160
rect 15657 5151 15715 5157
rect 15657 5117 15669 5151
rect 15703 5148 15715 5151
rect 16482 5148 16488 5160
rect 15703 5120 16488 5148
rect 15703 5117 15715 5120
rect 15657 5111 15715 5117
rect 16482 5108 16488 5120
rect 16540 5108 16546 5160
rect 17862 5148 17868 5160
rect 17823 5120 17868 5148
rect 17862 5108 17868 5120
rect 17920 5108 17926 5160
rect 18598 5108 18604 5160
rect 18656 5148 18662 5160
rect 18785 5151 18843 5157
rect 18785 5148 18797 5151
rect 18656 5120 18797 5148
rect 18656 5108 18662 5120
rect 18785 5117 18797 5120
rect 18831 5117 18843 5151
rect 18785 5111 18843 5117
rect 19426 5108 19432 5160
rect 19484 5148 19490 5160
rect 19981 5151 20039 5157
rect 19981 5148 19993 5151
rect 19484 5120 19993 5148
rect 19484 5108 19490 5120
rect 19981 5117 19993 5120
rect 20027 5117 20039 5151
rect 19981 5111 20039 5117
rect 20625 5151 20683 5157
rect 20625 5117 20637 5151
rect 20671 5148 20683 5151
rect 22756 5148 22784 5179
rect 23106 5176 23112 5188
rect 23164 5176 23170 5228
rect 23216 5225 23244 5256
rect 26142 5244 26148 5296
rect 26200 5284 26206 5296
rect 26200 5256 30420 5284
rect 26200 5244 26206 5256
rect 23201 5219 23259 5225
rect 23201 5185 23213 5219
rect 23247 5185 23259 5219
rect 23201 5179 23259 5185
rect 24029 5219 24087 5225
rect 24029 5185 24041 5219
rect 24075 5185 24087 5219
rect 26418 5216 26424 5228
rect 26379 5188 26424 5216
rect 24029 5179 24087 5185
rect 20671 5120 22784 5148
rect 20671 5117 20683 5120
rect 20625 5111 20683 5117
rect 23014 5108 23020 5160
rect 23072 5148 23078 5160
rect 24044 5148 24072 5179
rect 26418 5176 26424 5188
rect 26476 5176 26482 5228
rect 30392 5225 30420 5256
rect 29549 5219 29607 5225
rect 29549 5185 29561 5219
rect 29595 5185 29607 5219
rect 29549 5179 29607 5185
rect 30377 5219 30435 5225
rect 30377 5185 30389 5219
rect 30423 5185 30435 5219
rect 30377 5179 30435 5185
rect 23072 5120 24072 5148
rect 29564 5148 29592 5179
rect 37918 5176 37924 5228
rect 37976 5216 37982 5228
rect 38013 5219 38071 5225
rect 38013 5216 38025 5219
rect 37976 5188 38025 5216
rect 37976 5176 37982 5188
rect 38013 5185 38025 5188
rect 38059 5185 38071 5219
rect 38013 5179 38071 5185
rect 38102 5148 38108 5160
rect 29564 5120 38108 5148
rect 23072 5108 23078 5120
rect 38102 5108 38108 5120
rect 38160 5108 38166 5160
rect 13170 5080 13176 5092
rect 9692 5052 13176 5080
rect 13170 5040 13176 5052
rect 13228 5040 13234 5092
rect 15194 5080 15200 5092
rect 15107 5052 15200 5080
rect 15194 5040 15200 5052
rect 15252 5080 15258 5092
rect 18138 5080 18144 5092
rect 15252 5052 18144 5080
rect 15252 5040 15258 5052
rect 18138 5040 18144 5052
rect 18196 5040 18202 5092
rect 20346 5080 20352 5092
rect 18248 5052 20352 5080
rect 18248 5024 18276 5052
rect 20346 5040 20352 5052
rect 20404 5040 20410 5092
rect 21542 5040 21548 5092
rect 21600 5080 21606 5092
rect 21910 5080 21916 5092
rect 21600 5052 21916 5080
rect 21600 5040 21606 5052
rect 21910 5040 21916 5052
rect 21968 5080 21974 5092
rect 21968 5052 29684 5080
rect 21968 5040 21974 5052
rect 10410 5012 10416 5024
rect 7852 4984 10416 5012
rect 5721 4975 5779 4981
rect 10410 4972 10416 4984
rect 10468 4972 10474 5024
rect 11057 5015 11115 5021
rect 11057 4981 11069 5015
rect 11103 5012 11115 5015
rect 14182 5012 14188 5024
rect 11103 4984 14188 5012
rect 11103 4981 11115 4984
rect 11057 4975 11115 4981
rect 14182 4972 14188 4984
rect 14240 4972 14246 5024
rect 16301 5015 16359 5021
rect 16301 4981 16313 5015
rect 16347 5012 16359 5015
rect 18230 5012 18236 5024
rect 16347 4984 18236 5012
rect 16347 4981 16359 4984
rect 16301 4975 16359 4981
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 18322 4972 18328 5024
rect 18380 5012 18386 5024
rect 21177 5015 21235 5021
rect 21177 5012 21189 5015
rect 18380 4984 21189 5012
rect 18380 4972 18386 4984
rect 21177 4981 21189 4984
rect 21223 4981 21235 5015
rect 21177 4975 21235 4981
rect 21726 4972 21732 5024
rect 21784 5012 21790 5024
rect 23293 5015 23351 5021
rect 23293 5012 23305 5015
rect 21784 4984 23305 5012
rect 21784 4972 21790 4984
rect 23293 4981 23305 4984
rect 23339 4981 23351 5015
rect 23293 4975 23351 4981
rect 26237 5015 26295 5021
rect 26237 4981 26249 5015
rect 26283 5012 26295 5015
rect 29454 5012 29460 5024
rect 26283 4984 29460 5012
rect 26283 4981 26295 4984
rect 26237 4975 26295 4981
rect 29454 4972 29460 4984
rect 29512 4972 29518 5024
rect 29656 5021 29684 5052
rect 29641 5015 29699 5021
rect 29641 4981 29653 5015
rect 29687 4981 29699 5015
rect 29641 4975 29699 4981
rect 30193 5015 30251 5021
rect 30193 4981 30205 5015
rect 30239 5012 30251 5015
rect 33042 5012 33048 5024
rect 30239 4984 33048 5012
rect 30239 4981 30251 4984
rect 30193 4975 30251 4981
rect 33042 4972 33048 4984
rect 33100 4972 33106 5024
rect 38194 5012 38200 5024
rect 38155 4984 38200 5012
rect 38194 4972 38200 4984
rect 38252 4972 38258 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 1936 4811 1994 4817
rect 1936 4777 1948 4811
rect 1982 4808 1994 4811
rect 3142 4808 3148 4820
rect 1982 4780 3148 4808
rect 1982 4777 1994 4780
rect 1936 4771 1994 4777
rect 3142 4768 3148 4780
rect 3200 4768 3206 4820
rect 3970 4768 3976 4820
rect 4028 4808 4034 4820
rect 4065 4811 4123 4817
rect 4065 4808 4077 4811
rect 4028 4780 4077 4808
rect 4028 4768 4034 4780
rect 4065 4777 4077 4780
rect 4111 4777 4123 4811
rect 7374 4808 7380 4820
rect 4065 4771 4123 4777
rect 6196 4780 7380 4808
rect 3694 4700 3700 4752
rect 3752 4740 3758 4752
rect 6196 4740 6224 4780
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 9940 4811 9998 4817
rect 9940 4777 9952 4811
rect 9986 4808 9998 4811
rect 13262 4808 13268 4820
rect 9986 4780 13268 4808
rect 9986 4777 9998 4780
rect 9940 4771 9998 4777
rect 13262 4768 13268 4780
rect 13320 4768 13326 4820
rect 13832 4780 16712 4808
rect 3752 4712 6224 4740
rect 3752 4700 3758 4712
rect 13354 4700 13360 4752
rect 13412 4740 13418 4752
rect 13725 4743 13783 4749
rect 13725 4740 13737 4743
rect 13412 4712 13737 4740
rect 13412 4700 13418 4712
rect 13725 4709 13737 4712
rect 13771 4709 13783 4743
rect 13725 4703 13783 4709
rect 1578 4632 1584 4684
rect 1636 4672 1642 4684
rect 1673 4675 1731 4681
rect 1673 4672 1685 4675
rect 1636 4644 1685 4672
rect 1636 4632 1642 4644
rect 1673 4641 1685 4644
rect 1719 4672 1731 4675
rect 3326 4672 3332 4684
rect 1719 4644 3332 4672
rect 1719 4641 1731 4644
rect 1673 4635 1731 4641
rect 3326 4632 3332 4644
rect 3384 4632 3390 4684
rect 5258 4632 5264 4684
rect 5316 4672 5322 4684
rect 6089 4675 6147 4681
rect 6089 4672 6101 4675
rect 5316 4644 6101 4672
rect 5316 4632 5322 4644
rect 6089 4641 6101 4644
rect 6135 4641 6147 4675
rect 6089 4635 6147 4641
rect 6365 4675 6423 4681
rect 6365 4641 6377 4675
rect 6411 4672 6423 4675
rect 7098 4672 7104 4684
rect 6411 4644 7104 4672
rect 6411 4641 6423 4644
rect 6365 4635 6423 4641
rect 7098 4632 7104 4644
rect 7156 4632 7162 4684
rect 9398 4632 9404 4684
rect 9456 4672 9462 4684
rect 9677 4675 9735 4681
rect 9677 4672 9689 4675
rect 9456 4644 9689 4672
rect 9456 4632 9462 4644
rect 9677 4641 9689 4644
rect 9723 4672 9735 4675
rect 11146 4672 11152 4684
rect 9723 4644 11152 4672
rect 9723 4641 9735 4644
rect 9677 4635 9735 4641
rect 11146 4632 11152 4644
rect 11204 4672 11210 4684
rect 11977 4675 12035 4681
rect 11977 4672 11989 4675
rect 11204 4644 11989 4672
rect 11204 4632 11210 4644
rect 11977 4641 11989 4644
rect 12023 4641 12035 4675
rect 13832 4672 13860 4780
rect 16022 4740 16028 4752
rect 15983 4712 16028 4740
rect 16022 4700 16028 4712
rect 16080 4700 16086 4752
rect 11977 4635 12035 4641
rect 13372 4644 13860 4672
rect 3602 4564 3608 4616
rect 3660 4604 3666 4616
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 3660 4576 3985 4604
rect 3660 4564 3666 4576
rect 3973 4573 3985 4576
rect 4019 4604 4031 4607
rect 4801 4607 4859 4613
rect 4801 4604 4813 4607
rect 4019 4576 4813 4604
rect 4019 4573 4031 4576
rect 3973 4567 4031 4573
rect 4801 4573 4813 4576
rect 4847 4604 4859 4607
rect 5445 4607 5503 4613
rect 5445 4604 5457 4607
rect 4847 4576 5457 4604
rect 4847 4573 4859 4576
rect 4801 4567 4859 4573
rect 5445 4573 5457 4576
rect 5491 4573 5503 4607
rect 5445 4567 5503 4573
rect 11054 4564 11060 4616
rect 11112 4564 11118 4616
rect 13372 4590 13400 4644
rect 14182 4632 14188 4684
rect 14240 4672 14246 4684
rect 16577 4675 16635 4681
rect 16577 4672 16589 4675
rect 14240 4644 16589 4672
rect 14240 4632 14246 4644
rect 16577 4641 16589 4644
rect 16623 4641 16635 4675
rect 16684 4672 16712 4780
rect 17034 4768 17040 4820
rect 17092 4808 17098 4820
rect 23201 4811 23259 4817
rect 23201 4808 23213 4811
rect 17092 4780 23213 4808
rect 17092 4768 17098 4780
rect 23201 4777 23213 4780
rect 23247 4777 23259 4811
rect 23842 4808 23848 4820
rect 23803 4780 23848 4808
rect 23201 4771 23259 4777
rect 23842 4768 23848 4780
rect 23900 4768 23906 4820
rect 17129 4743 17187 4749
rect 17129 4709 17141 4743
rect 17175 4740 17187 4743
rect 17218 4740 17224 4752
rect 17175 4712 17224 4740
rect 17175 4709 17187 4712
rect 17129 4703 17187 4709
rect 17218 4700 17224 4712
rect 17276 4700 17282 4752
rect 17586 4700 17592 4752
rect 17644 4740 17650 4752
rect 24673 4743 24731 4749
rect 24673 4740 24685 4743
rect 17644 4712 24685 4740
rect 17644 4700 17650 4712
rect 24673 4709 24685 4712
rect 24719 4709 24731 4743
rect 24673 4703 24731 4709
rect 18230 4672 18236 4684
rect 16684 4644 17264 4672
rect 18191 4644 18236 4672
rect 16577 4635 16635 4641
rect 13722 4564 13728 4616
rect 13780 4604 13786 4616
rect 14277 4607 14335 4613
rect 14277 4604 14289 4607
rect 13780 4576 14289 4604
rect 13780 4564 13786 4576
rect 14277 4573 14289 4576
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 4893 4539 4951 4545
rect 4893 4536 4905 4539
rect 3174 4508 4905 4536
rect 4893 4505 4905 4508
rect 4939 4505 4951 4539
rect 7926 4536 7932 4548
rect 7590 4508 7932 4536
rect 4893 4499 4951 4505
rect 7926 4496 7932 4508
rect 7984 4496 7990 4548
rect 8110 4536 8116 4548
rect 8071 4508 8116 4536
rect 8110 4496 8116 4508
rect 8168 4496 8174 4548
rect 12158 4496 12164 4548
rect 12216 4536 12222 4548
rect 12253 4539 12311 4545
rect 12253 4536 12265 4539
rect 12216 4508 12265 4536
rect 12216 4496 12222 4508
rect 12253 4505 12265 4508
rect 12299 4505 12311 4539
rect 12253 4499 12311 4505
rect 13630 4496 13636 4548
rect 13688 4536 13694 4548
rect 14553 4539 14611 4545
rect 14553 4536 14565 4539
rect 13688 4508 14565 4536
rect 13688 4496 13694 4508
rect 14553 4505 14565 4508
rect 14599 4505 14611 4539
rect 14553 4499 14611 4505
rect 15562 4496 15568 4548
rect 15620 4496 15626 4548
rect 16574 4536 16580 4548
rect 15856 4508 16580 4536
rect 3421 4471 3479 4477
rect 3421 4437 3433 4471
rect 3467 4468 3479 4471
rect 3510 4468 3516 4480
rect 3467 4440 3516 4468
rect 3467 4437 3479 4440
rect 3421 4431 3479 4437
rect 3510 4428 3516 4440
rect 3568 4428 3574 4480
rect 4614 4428 4620 4480
rect 4672 4468 4678 4480
rect 5537 4471 5595 4477
rect 5537 4468 5549 4471
rect 4672 4440 5549 4468
rect 4672 4428 4678 4440
rect 5537 4437 5549 4440
rect 5583 4437 5595 4471
rect 5537 4431 5595 4437
rect 5994 4428 6000 4480
rect 6052 4468 6058 4480
rect 9674 4468 9680 4480
rect 6052 4440 9680 4468
rect 6052 4428 6058 4440
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 9950 4428 9956 4480
rect 10008 4468 10014 4480
rect 11422 4468 11428 4480
rect 10008 4440 11428 4468
rect 10008 4428 10014 4440
rect 11422 4428 11428 4440
rect 11480 4428 11486 4480
rect 13170 4428 13176 4480
rect 13228 4468 13234 4480
rect 15856 4468 15884 4508
rect 16574 4496 16580 4508
rect 16632 4496 16638 4548
rect 16669 4539 16727 4545
rect 16669 4505 16681 4539
rect 16715 4505 16727 4539
rect 17236 4536 17264 4644
rect 18230 4632 18236 4644
rect 18288 4632 18294 4684
rect 18506 4672 18512 4684
rect 18467 4644 18512 4672
rect 18506 4632 18512 4644
rect 18564 4632 18570 4684
rect 18874 4632 18880 4684
rect 18932 4672 18938 4684
rect 19613 4675 19671 4681
rect 18932 4644 19564 4672
rect 18932 4632 18938 4644
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4573 19487 4607
rect 19536 4604 19564 4644
rect 19613 4641 19625 4675
rect 19659 4672 19671 4675
rect 21269 4675 21327 4681
rect 21269 4672 21281 4675
rect 19659 4644 21281 4672
rect 19659 4641 19671 4644
rect 19613 4635 19671 4641
rect 21269 4641 21281 4644
rect 21315 4641 21327 4675
rect 21269 4635 21327 4641
rect 21836 4644 22876 4672
rect 20346 4606 20352 4616
rect 19996 4604 20352 4606
rect 19536 4578 20352 4604
rect 19536 4576 20024 4578
rect 19429 4567 19487 4573
rect 17236 4508 18277 4536
rect 16669 4499 16727 4505
rect 13228 4440 15884 4468
rect 16684 4468 16712 4499
rect 18046 4468 18052 4480
rect 16684 4440 18052 4468
rect 13228 4428 13234 4440
rect 18046 4428 18052 4440
rect 18104 4428 18110 4480
rect 18249 4468 18277 4508
rect 18322 4496 18328 4548
rect 18380 4536 18386 4548
rect 19444 4536 19472 4567
rect 20346 4564 20352 4578
rect 20404 4564 20410 4616
rect 20530 4604 20536 4616
rect 20491 4576 20536 4604
rect 20530 4564 20536 4576
rect 20588 4604 20594 4616
rect 20806 4604 20812 4616
rect 20588 4576 20812 4604
rect 20588 4564 20594 4576
rect 20806 4564 20812 4576
rect 20864 4564 20870 4616
rect 21174 4604 21180 4616
rect 21135 4576 21180 4604
rect 21174 4564 21180 4576
rect 21232 4564 21238 4616
rect 21836 4613 21864 4644
rect 21821 4607 21879 4613
rect 21821 4573 21833 4607
rect 21867 4573 21879 4607
rect 21821 4567 21879 4573
rect 19702 4536 19708 4548
rect 18380 4508 18425 4536
rect 19444 4508 19708 4536
rect 18380 4496 18386 4508
rect 19702 4496 19708 4508
rect 19760 4496 19766 4548
rect 20073 4539 20131 4545
rect 20073 4505 20085 4539
rect 20119 4536 20131 4539
rect 20162 4536 20168 4548
rect 20119 4508 20168 4536
rect 20119 4505 20131 4508
rect 20073 4499 20131 4505
rect 20162 4496 20168 4508
rect 20220 4496 20226 4548
rect 20254 4496 20260 4548
rect 20312 4536 20318 4548
rect 22465 4539 22523 4545
rect 22465 4536 22477 4539
rect 20312 4508 22477 4536
rect 20312 4496 20318 4508
rect 22465 4505 22477 4508
rect 22511 4505 22523 4539
rect 22848 4536 22876 4644
rect 23106 4604 23112 4616
rect 23067 4576 23112 4604
rect 23106 4564 23112 4576
rect 23164 4564 23170 4616
rect 23750 4604 23756 4616
rect 23711 4576 23756 4604
rect 23750 4564 23756 4576
rect 23808 4564 23814 4616
rect 24394 4564 24400 4616
rect 24452 4604 24458 4616
rect 24581 4607 24639 4613
rect 24581 4604 24593 4607
rect 24452 4576 24593 4604
rect 24452 4564 24458 4576
rect 24581 4573 24593 4576
rect 24627 4573 24639 4607
rect 24581 4567 24639 4573
rect 25225 4607 25283 4613
rect 25225 4573 25237 4607
rect 25271 4604 25283 4607
rect 27798 4604 27804 4616
rect 25271 4576 27804 4604
rect 25271 4573 25283 4576
rect 25225 4567 25283 4573
rect 27798 4564 27804 4576
rect 27856 4564 27862 4616
rect 37734 4564 37740 4616
rect 37792 4604 37798 4616
rect 38013 4607 38071 4613
rect 38013 4604 38025 4607
rect 37792 4576 38025 4604
rect 37792 4564 37798 4576
rect 38013 4573 38025 4576
rect 38059 4573 38071 4607
rect 38013 4567 38071 4573
rect 23566 4536 23572 4548
rect 22848 4508 23572 4536
rect 22465 4499 22523 4505
rect 23566 4496 23572 4508
rect 23624 4496 23630 4548
rect 25317 4539 25375 4545
rect 25317 4536 25329 4539
rect 23676 4508 25329 4536
rect 19794 4468 19800 4480
rect 18249 4440 19800 4468
rect 19794 4428 19800 4440
rect 19852 4428 19858 4480
rect 20346 4428 20352 4480
rect 20404 4468 20410 4480
rect 20625 4471 20683 4477
rect 20625 4468 20637 4471
rect 20404 4440 20637 4468
rect 20404 4428 20410 4440
rect 20625 4437 20637 4440
rect 20671 4437 20683 4471
rect 20625 4431 20683 4437
rect 20714 4428 20720 4480
rect 20772 4468 20778 4480
rect 21913 4471 21971 4477
rect 21913 4468 21925 4471
rect 20772 4440 21925 4468
rect 20772 4428 20778 4440
rect 21913 4437 21925 4440
rect 21959 4437 21971 4471
rect 21913 4431 21971 4437
rect 22278 4428 22284 4480
rect 22336 4468 22342 4480
rect 23676 4468 23704 4508
rect 25317 4505 25329 4508
rect 25363 4505 25375 4539
rect 25317 4499 25375 4505
rect 22336 4440 23704 4468
rect 37829 4471 37887 4477
rect 22336 4428 22342 4440
rect 37829 4437 37841 4471
rect 37875 4468 37887 4471
rect 38010 4468 38016 4480
rect 37875 4440 38016 4468
rect 37875 4437 37887 4440
rect 37829 4431 37887 4437
rect 38010 4428 38016 4440
rect 38068 4428 38074 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 8294 4264 8300 4276
rect 3988 4236 6040 4264
rect 1670 4196 1676 4208
rect 1631 4168 1676 4196
rect 1670 4156 1676 4168
rect 1728 4156 1734 4208
rect 3510 4156 3516 4208
rect 3568 4196 3574 4208
rect 3612 4199 3670 4205
rect 3612 4196 3624 4199
rect 3568 4168 3624 4196
rect 3568 4156 3574 4168
rect 3612 4165 3624 4168
rect 3658 4196 3670 4199
rect 3988 4196 4016 4236
rect 3658 4168 4016 4196
rect 3658 4165 3670 4168
rect 3612 4159 3670 4165
rect 4614 4156 4620 4208
rect 4672 4156 4678 4208
rect 6012 4196 6040 4236
rect 7208 4236 8300 4264
rect 7098 4196 7104 4208
rect 6012 4168 7104 4196
rect 1857 4131 1915 4137
rect 1857 4097 1869 4131
rect 1903 4128 1915 4131
rect 2038 4128 2044 4140
rect 1903 4100 2044 4128
rect 1903 4097 1915 4100
rect 1857 4091 1915 4097
rect 2038 4088 2044 4100
rect 2096 4088 2102 4140
rect 2869 4131 2927 4137
rect 2869 4097 2881 4131
rect 2915 4097 2927 4131
rect 3326 4128 3332 4140
rect 3287 4100 3332 4128
rect 2869 4091 2927 4097
rect 2884 4060 2912 4091
rect 3326 4088 3332 4100
rect 3384 4088 3390 4140
rect 6012 4137 6040 4168
rect 7098 4156 7104 4168
rect 7156 4156 7162 4208
rect 5997 4131 6055 4137
rect 5997 4097 6009 4131
rect 6043 4097 6055 4131
rect 6546 4128 6552 4140
rect 6507 4100 6552 4128
rect 5997 4091 6055 4097
rect 6546 4088 6552 4100
rect 6604 4088 6610 4140
rect 7208 4137 7236 4236
rect 8294 4224 8300 4236
rect 8352 4224 8358 4276
rect 9214 4224 9220 4276
rect 9272 4264 9278 4276
rect 10502 4264 10508 4276
rect 9272 4236 10508 4264
rect 9272 4224 9278 4236
rect 10502 4224 10508 4236
rect 10560 4224 10566 4276
rect 11422 4224 11428 4276
rect 11480 4264 11486 4276
rect 18601 4267 18659 4273
rect 11480 4236 18460 4264
rect 11480 4224 11486 4236
rect 9582 4196 9588 4208
rect 8694 4168 9588 4196
rect 9582 4156 9588 4168
rect 9640 4156 9646 4208
rect 9674 4156 9680 4208
rect 9732 4196 9738 4208
rect 13446 4196 13452 4208
rect 9732 4168 10166 4196
rect 13280 4168 13452 4196
rect 9732 4156 9738 4168
rect 7193 4131 7251 4137
rect 7193 4097 7205 4131
rect 7239 4097 7251 4131
rect 9398 4128 9404 4140
rect 9359 4100 9404 4128
rect 7193 4091 7251 4097
rect 9398 4088 9404 4100
rect 9456 4088 9462 4140
rect 11514 4088 11520 4140
rect 11572 4128 11578 4140
rect 13280 4137 13308 4168
rect 13446 4156 13452 4168
rect 13504 4156 13510 4208
rect 13541 4199 13599 4205
rect 13541 4165 13553 4199
rect 13587 4196 13599 4199
rect 13814 4196 13820 4208
rect 13587 4168 13820 4196
rect 13587 4165 13599 4168
rect 13541 4159 13599 4165
rect 13814 4156 13820 4168
rect 13872 4156 13878 4208
rect 13998 4156 14004 4208
rect 14056 4156 14062 4208
rect 16574 4156 16580 4208
rect 16632 4196 16638 4208
rect 17402 4196 17408 4208
rect 16632 4168 17408 4196
rect 16632 4156 16638 4168
rect 17402 4156 17408 4168
rect 17460 4156 17466 4208
rect 18432 4196 18460 4236
rect 18601 4233 18613 4267
rect 18647 4264 18659 4267
rect 19150 4264 19156 4276
rect 18647 4236 19156 4264
rect 18647 4233 18659 4236
rect 18601 4227 18659 4233
rect 19150 4224 19156 4236
rect 19208 4264 19214 4276
rect 19208 4236 19564 4264
rect 19208 4224 19214 4236
rect 19536 4196 19564 4236
rect 19610 4224 19616 4276
rect 19668 4264 19674 4276
rect 20625 4267 20683 4273
rect 20625 4264 20637 4267
rect 19668 4236 20637 4264
rect 19668 4224 19674 4236
rect 20625 4233 20637 4236
rect 20671 4233 20683 4267
rect 23106 4264 23112 4276
rect 20625 4227 20683 4233
rect 20732 4236 23112 4264
rect 20732 4196 20760 4236
rect 23106 4224 23112 4236
rect 23164 4224 23170 4276
rect 23658 4224 23664 4276
rect 23716 4264 23722 4276
rect 24394 4264 24400 4276
rect 23716 4236 24400 4264
rect 23716 4224 23722 4236
rect 24394 4224 24400 4236
rect 24452 4224 24458 4276
rect 18432 4168 19380 4196
rect 19536 4168 20760 4196
rect 11977 4131 12035 4137
rect 11977 4128 11989 4131
rect 11572 4100 11989 4128
rect 11572 4088 11578 4100
rect 11977 4097 11989 4100
rect 12023 4097 12035 4131
rect 11977 4091 12035 4097
rect 12621 4131 12679 4137
rect 12621 4097 12633 4131
rect 12667 4097 12679 4131
rect 12621 4091 12679 4097
rect 13265 4131 13323 4137
rect 13265 4097 13277 4131
rect 13311 4097 13323 4131
rect 13265 4091 13323 4097
rect 6454 4060 6460 4072
rect 2884 4032 6460 4060
rect 6454 4020 6460 4032
rect 6512 4020 6518 4072
rect 7469 4063 7527 4069
rect 7469 4029 7481 4063
rect 7515 4060 7527 4063
rect 8110 4060 8116 4072
rect 7515 4032 8116 4060
rect 7515 4029 7527 4032
rect 7469 4023 7527 4029
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 9677 4063 9735 4069
rect 9677 4029 9689 4063
rect 9723 4060 9735 4063
rect 12526 4060 12532 4072
rect 9723 4032 12532 4060
rect 9723 4029 9735 4032
rect 9677 4023 9735 4029
rect 12526 4020 12532 4032
rect 12584 4020 12590 4072
rect 5077 3995 5135 4001
rect 5077 3961 5089 3995
rect 5123 3992 5135 3995
rect 5442 3992 5448 4004
rect 5123 3964 5448 3992
rect 5123 3961 5135 3964
rect 5077 3955 5135 3961
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 5902 3952 5908 4004
rect 5960 3992 5966 4004
rect 6641 3995 6699 4001
rect 6641 3992 6653 3995
rect 5960 3964 6653 3992
rect 5960 3952 5966 3964
rect 6641 3961 6653 3964
rect 6687 3961 6699 3995
rect 6641 3955 6699 3961
rect 11606 3952 11612 4004
rect 11664 3992 11670 4004
rect 12066 3992 12072 4004
rect 11664 3964 11836 3992
rect 12027 3964 12072 3992
rect 11664 3952 11670 3964
rect 2685 3927 2743 3933
rect 2685 3893 2697 3927
rect 2731 3924 2743 3927
rect 3970 3924 3976 3936
rect 2731 3896 3976 3924
rect 2731 3893 2743 3896
rect 2685 3887 2743 3893
rect 3970 3884 3976 3896
rect 4028 3884 4034 3936
rect 4614 3884 4620 3936
rect 4672 3924 4678 3936
rect 5534 3924 5540 3936
rect 4672 3896 5540 3924
rect 4672 3884 4678 3896
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 5626 3884 5632 3936
rect 5684 3924 5690 3936
rect 5813 3927 5871 3933
rect 5813 3924 5825 3927
rect 5684 3896 5825 3924
rect 5684 3884 5690 3896
rect 5813 3893 5825 3896
rect 5859 3893 5871 3927
rect 5813 3887 5871 3893
rect 7098 3884 7104 3936
rect 7156 3924 7162 3936
rect 8941 3927 8999 3933
rect 8941 3924 8953 3927
rect 7156 3896 8953 3924
rect 7156 3884 7162 3896
rect 8941 3893 8953 3896
rect 8987 3924 8999 3927
rect 9858 3924 9864 3936
rect 8987 3896 9864 3924
rect 8987 3893 8999 3896
rect 8941 3887 8999 3893
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 11149 3927 11207 3933
rect 11149 3893 11161 3927
rect 11195 3924 11207 3927
rect 11698 3924 11704 3936
rect 11195 3896 11704 3924
rect 11195 3893 11207 3896
rect 11149 3887 11207 3893
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 11808 3924 11836 3964
rect 12066 3952 12072 3964
rect 12124 3952 12130 4004
rect 12158 3952 12164 4004
rect 12216 3992 12222 4004
rect 12636 3992 12664 4091
rect 14826 4088 14832 4140
rect 14884 4128 14890 4140
rect 14884 4100 15332 4128
rect 14884 4088 14890 4100
rect 12713 4063 12771 4069
rect 12713 4029 12725 4063
rect 12759 4060 12771 4063
rect 15194 4060 15200 4072
rect 12759 4032 15200 4060
rect 12759 4029 12771 4032
rect 12713 4023 12771 4029
rect 15194 4020 15200 4032
rect 15252 4020 15258 4072
rect 15304 4069 15332 4100
rect 15470 4088 15476 4140
rect 15528 4128 15534 4140
rect 16117 4131 16175 4137
rect 16117 4128 16129 4131
rect 15528 4100 16129 4128
rect 15528 4088 15534 4100
rect 16117 4097 16129 4100
rect 16163 4097 16175 4131
rect 16117 4091 16175 4097
rect 16206 4088 16212 4140
rect 16264 4128 16270 4140
rect 16758 4128 16764 4140
rect 16264 4100 16309 4128
rect 16684 4100 16764 4128
rect 16264 4088 16270 4100
rect 15289 4063 15347 4069
rect 15289 4029 15301 4063
rect 15335 4060 15347 4063
rect 16684 4060 16712 4100
rect 16758 4088 16764 4100
rect 16816 4088 16822 4140
rect 18230 4088 18236 4140
rect 18288 4088 18294 4140
rect 19245 4131 19303 4137
rect 19245 4097 19257 4131
rect 19291 4097 19303 4131
rect 19352 4128 19380 4168
rect 20806 4156 20812 4208
rect 20864 4196 20870 4208
rect 23198 4196 23204 4208
rect 20864 4168 23204 4196
rect 20864 4156 20870 4168
rect 23198 4156 23204 4168
rect 23256 4196 23262 4208
rect 23256 4168 23336 4196
rect 23256 4156 23262 4168
rect 19889 4131 19947 4137
rect 19889 4128 19901 4131
rect 19352 4100 19901 4128
rect 19245 4091 19303 4097
rect 19889 4097 19901 4100
rect 19935 4097 19947 4131
rect 19889 4091 19947 4097
rect 16850 4060 16856 4072
rect 15335 4032 16712 4060
rect 16811 4032 16856 4060
rect 15335 4029 15347 4032
rect 15289 4023 15347 4029
rect 16850 4020 16856 4032
rect 16908 4020 16914 4072
rect 17129 4063 17187 4069
rect 17129 4060 17141 4063
rect 16960 4032 17141 4060
rect 12216 3964 12664 3992
rect 12216 3952 12222 3964
rect 14550 3952 14556 4004
rect 14608 3992 14614 4004
rect 16022 3992 16028 4004
rect 14608 3964 16028 3992
rect 14608 3952 14614 3964
rect 16022 3952 16028 3964
rect 16080 3952 16086 4004
rect 16114 3952 16120 4004
rect 16172 3992 16178 4004
rect 16960 3992 16988 4032
rect 17129 4029 17141 4032
rect 17175 4029 17187 4063
rect 17129 4023 17187 4029
rect 18138 4020 18144 4072
rect 18196 4060 18202 4072
rect 19260 4060 19288 4091
rect 19978 4088 19984 4140
rect 20036 4128 20042 4140
rect 20036 4100 20081 4128
rect 20036 4088 20042 4100
rect 20254 4088 20260 4140
rect 20312 4128 20318 4140
rect 20533 4131 20591 4137
rect 20533 4128 20545 4131
rect 20312 4100 20545 4128
rect 20312 4088 20318 4100
rect 20533 4097 20545 4100
rect 20579 4097 20591 4131
rect 21177 4131 21235 4137
rect 21177 4128 21189 4131
rect 20533 4091 20591 4097
rect 20640 4100 21189 4128
rect 20640 4060 20668 4100
rect 21177 4097 21189 4100
rect 21223 4097 21235 4131
rect 22002 4128 22008 4140
rect 21963 4100 22008 4128
rect 21177 4091 21235 4097
rect 22002 4088 22008 4100
rect 22060 4088 22066 4140
rect 22278 4088 22284 4140
rect 22336 4128 22342 4140
rect 23308 4137 23336 4168
rect 22649 4131 22707 4137
rect 22649 4128 22661 4131
rect 22336 4100 22661 4128
rect 22336 4088 22342 4100
rect 22649 4097 22661 4100
rect 22695 4097 22707 4131
rect 22649 4091 22707 4097
rect 23293 4131 23351 4137
rect 23293 4097 23305 4131
rect 23339 4097 23351 4131
rect 23293 4091 23351 4097
rect 23566 4088 23572 4140
rect 23624 4128 23630 4140
rect 23937 4131 23995 4137
rect 23937 4128 23949 4131
rect 23624 4100 23949 4128
rect 23624 4088 23630 4100
rect 23937 4097 23949 4100
rect 23983 4128 23995 4131
rect 24581 4131 24639 4137
rect 24581 4128 24593 4131
rect 23983 4100 24593 4128
rect 23983 4097 23995 4100
rect 23937 4091 23995 4097
rect 24581 4097 24593 4100
rect 24627 4097 24639 4131
rect 24581 4091 24639 4097
rect 24670 4088 24676 4140
rect 24728 4128 24734 4140
rect 25225 4131 25283 4137
rect 24728 4100 24773 4128
rect 24728 4088 24734 4100
rect 25225 4097 25237 4131
rect 25271 4097 25283 4131
rect 26050 4128 26056 4140
rect 26011 4100 26056 4128
rect 25225 4091 25283 4097
rect 18196 4032 19288 4060
rect 20456 4032 20668 4060
rect 18196 4020 18202 4032
rect 20456 3992 20484 4032
rect 20806 4020 20812 4072
rect 20864 4060 20870 4072
rect 21269 4063 21327 4069
rect 21269 4060 21281 4063
rect 20864 4032 21281 4060
rect 20864 4020 20870 4032
rect 21269 4029 21281 4032
rect 21315 4029 21327 4063
rect 21269 4023 21327 4029
rect 21542 4020 21548 4072
rect 21600 4060 21606 4072
rect 24029 4063 24087 4069
rect 24029 4060 24041 4063
rect 21600 4032 24041 4060
rect 21600 4020 21606 4032
rect 24029 4029 24041 4032
rect 24075 4029 24087 4063
rect 24029 4023 24087 4029
rect 22738 3992 22744 4004
rect 16172 3964 16988 3992
rect 18156 3964 20484 3992
rect 22699 3964 22744 3992
rect 16172 3952 16178 3964
rect 12618 3924 12624 3936
rect 11808 3896 12624 3924
rect 12618 3884 12624 3896
rect 12676 3884 12682 3936
rect 12986 3884 12992 3936
rect 13044 3924 13050 3936
rect 18156 3924 18184 3964
rect 22738 3952 22744 3964
rect 22796 3952 22802 4004
rect 25240 3992 25268 4091
rect 26050 4088 26056 4100
rect 26108 4088 26114 4140
rect 38286 4128 38292 4140
rect 38247 4100 38292 4128
rect 38286 4088 38292 4100
rect 38344 4088 38350 4140
rect 25774 3992 25780 4004
rect 23216 3964 25780 3992
rect 13044 3896 18184 3924
rect 19337 3927 19395 3933
rect 13044 3884 13050 3896
rect 19337 3893 19349 3927
rect 19383 3924 19395 3927
rect 20990 3924 20996 3936
rect 19383 3896 20996 3924
rect 19383 3893 19395 3896
rect 19337 3887 19395 3893
rect 20990 3884 20996 3896
rect 21048 3884 21054 3936
rect 21082 3884 21088 3936
rect 21140 3924 21146 3936
rect 22097 3927 22155 3933
rect 22097 3924 22109 3927
rect 21140 3896 22109 3924
rect 21140 3884 21146 3896
rect 22097 3893 22109 3896
rect 22143 3893 22155 3927
rect 22097 3887 22155 3893
rect 22554 3884 22560 3936
rect 22612 3924 22618 3936
rect 23216 3924 23244 3964
rect 25774 3952 25780 3964
rect 25832 3952 25838 4004
rect 31386 3952 31392 4004
rect 31444 3992 31450 4004
rect 38105 3995 38163 4001
rect 38105 3992 38117 3995
rect 31444 3964 38117 3992
rect 31444 3952 31450 3964
rect 38105 3961 38117 3964
rect 38151 3961 38163 3995
rect 38105 3955 38163 3961
rect 23382 3924 23388 3936
rect 22612 3896 23244 3924
rect 23343 3896 23388 3924
rect 22612 3884 22618 3896
rect 23382 3884 23388 3896
rect 23440 3884 23446 3936
rect 25314 3924 25320 3936
rect 25275 3896 25320 3924
rect 25314 3884 25320 3896
rect 25372 3884 25378 3936
rect 25869 3927 25927 3933
rect 25869 3893 25881 3927
rect 25915 3924 25927 3927
rect 27430 3924 27436 3936
rect 25915 3896 27436 3924
rect 25915 3893 25927 3896
rect 25869 3887 25927 3893
rect 27430 3884 27436 3896
rect 27488 3884 27494 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 1949 3723 2007 3729
rect 1949 3689 1961 3723
rect 1995 3720 2007 3723
rect 6546 3720 6552 3732
rect 1995 3692 6552 3720
rect 1995 3689 2007 3692
rect 1949 3683 2007 3689
rect 6546 3680 6552 3692
rect 6604 3680 6610 3732
rect 11606 3720 11612 3732
rect 6932 3692 11612 3720
rect 3878 3652 3884 3664
rect 2148 3624 3884 3652
rect 2148 3525 2176 3624
rect 3878 3612 3884 3624
rect 3936 3612 3942 3664
rect 6932 3652 6960 3692
rect 11606 3680 11612 3692
rect 11664 3680 11670 3732
rect 11698 3680 11704 3732
rect 11756 3720 11762 3732
rect 13354 3720 13360 3732
rect 11756 3692 13360 3720
rect 11756 3680 11762 3692
rect 13354 3680 13360 3692
rect 13412 3680 13418 3732
rect 13446 3680 13452 3732
rect 13504 3720 13510 3732
rect 16022 3720 16028 3732
rect 13504 3692 15608 3720
rect 15983 3692 16028 3720
rect 13504 3680 13510 3692
rect 3988 3624 6132 3652
rect 3988 3584 4016 3624
rect 3436 3556 4016 3584
rect 3436 3525 3464 3556
rect 4062 3544 4068 3596
rect 4120 3584 4126 3596
rect 5810 3584 5816 3596
rect 4120 3556 5816 3584
rect 4120 3544 4126 3556
rect 5810 3544 5816 3556
rect 5868 3544 5874 3596
rect 2133 3519 2191 3525
rect 2133 3485 2145 3519
rect 2179 3485 2191 3519
rect 2133 3479 2191 3485
rect 2777 3519 2835 3525
rect 2777 3485 2789 3519
rect 2823 3485 2835 3519
rect 2777 3479 2835 3485
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3485 3479 3519
rect 3421 3479 3479 3485
rect 4249 3519 4307 3525
rect 4249 3485 4261 3519
rect 4295 3516 4307 3519
rect 4614 3516 4620 3528
rect 4295 3488 4620 3516
rect 4295 3485 4307 3488
rect 4249 3479 4307 3485
rect 2792 3448 2820 3479
rect 4614 3476 4620 3488
rect 4672 3476 4678 3528
rect 4890 3516 4896 3528
rect 4851 3488 4896 3516
rect 4890 3476 4896 3488
rect 4948 3476 4954 3528
rect 4154 3448 4160 3460
rect 2792 3420 4160 3448
rect 4154 3408 4160 3420
rect 4212 3408 4218 3460
rect 4338 3448 4344 3460
rect 4299 3420 4344 3448
rect 4338 3408 4344 3420
rect 4396 3408 4402 3460
rect 2593 3383 2651 3389
rect 2593 3349 2605 3383
rect 2639 3380 2651 3383
rect 3142 3380 3148 3392
rect 2639 3352 3148 3380
rect 2639 3349 2651 3352
rect 2593 3343 2651 3349
rect 3142 3340 3148 3352
rect 3200 3340 3206 3392
rect 3237 3383 3295 3389
rect 3237 3349 3249 3383
rect 3283 3380 3295 3383
rect 4614 3380 4620 3392
rect 3283 3352 4620 3380
rect 3283 3349 3295 3352
rect 3237 3343 3295 3349
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 4985 3383 5043 3389
rect 4985 3349 4997 3383
rect 5031 3380 5043 3383
rect 5166 3380 5172 3392
rect 5031 3352 5172 3380
rect 5031 3349 5043 3352
rect 4985 3343 5043 3349
rect 5166 3340 5172 3352
rect 5224 3340 5230 3392
rect 5534 3380 5540 3392
rect 5495 3352 5540 3380
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 6104 3380 6132 3624
rect 6196 3624 6960 3652
rect 6196 3593 6224 3624
rect 8110 3612 8116 3664
rect 8168 3652 8174 3664
rect 8168 3624 11376 3652
rect 8168 3612 8174 3624
rect 6181 3587 6239 3593
rect 6181 3553 6193 3587
rect 6227 3553 6239 3587
rect 6181 3547 6239 3553
rect 6825 3587 6883 3593
rect 6825 3553 6837 3587
rect 6871 3584 6883 3587
rect 8294 3584 8300 3596
rect 6871 3556 8300 3584
rect 6871 3553 6883 3556
rect 6825 3547 6883 3553
rect 8294 3544 8300 3556
rect 8352 3544 8358 3596
rect 8386 3544 8392 3596
rect 8444 3584 8450 3596
rect 8573 3587 8631 3593
rect 8573 3584 8585 3587
rect 8444 3556 8585 3584
rect 8444 3544 8450 3556
rect 8573 3553 8585 3556
rect 8619 3553 8631 3587
rect 8573 3547 8631 3553
rect 8662 3544 8668 3596
rect 8720 3584 8726 3596
rect 9766 3584 9772 3596
rect 8720 3556 9772 3584
rect 8720 3544 8726 3556
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 10045 3587 10103 3593
rect 10045 3553 10057 3587
rect 10091 3584 10103 3587
rect 10870 3584 10876 3596
rect 10091 3556 10876 3584
rect 10091 3553 10103 3556
rect 10045 3547 10103 3553
rect 10870 3544 10876 3556
rect 10928 3544 10934 3596
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 11241 3587 11299 3593
rect 11241 3584 11253 3587
rect 11204 3556 11253 3584
rect 11204 3544 11210 3556
rect 11241 3553 11253 3556
rect 11287 3553 11299 3587
rect 11348 3584 11376 3624
rect 12526 3612 12532 3664
rect 12584 3652 12590 3664
rect 14182 3652 14188 3664
rect 12584 3624 14188 3652
rect 12584 3612 12590 3624
rect 14182 3612 14188 3624
rect 14240 3612 14246 3664
rect 15580 3652 15608 3692
rect 16022 3680 16028 3692
rect 16080 3720 16086 3732
rect 17586 3720 17592 3732
rect 16080 3692 17592 3720
rect 16080 3680 16086 3692
rect 17586 3680 17592 3692
rect 17644 3680 17650 3732
rect 17770 3680 17776 3732
rect 17828 3720 17834 3732
rect 18141 3723 18199 3729
rect 18141 3720 18153 3723
rect 17828 3692 18153 3720
rect 17828 3680 17834 3692
rect 18141 3689 18153 3692
rect 18187 3689 18199 3723
rect 18141 3683 18199 3689
rect 18322 3680 18328 3732
rect 18380 3720 18386 3732
rect 18785 3723 18843 3729
rect 18785 3720 18797 3723
rect 18380 3692 18797 3720
rect 18380 3680 18386 3692
rect 18785 3689 18797 3692
rect 18831 3689 18843 3723
rect 18785 3683 18843 3689
rect 19058 3680 19064 3732
rect 19116 3720 19122 3732
rect 19518 3720 19524 3732
rect 19116 3692 19524 3720
rect 19116 3680 19122 3692
rect 19518 3680 19524 3692
rect 19576 3680 19582 3732
rect 20257 3723 20315 3729
rect 20257 3689 20269 3723
rect 20303 3720 20315 3723
rect 22186 3720 22192 3732
rect 20303 3692 22192 3720
rect 20303 3689 20315 3692
rect 20257 3683 20315 3689
rect 22186 3680 22192 3692
rect 22244 3680 22250 3732
rect 22830 3720 22836 3732
rect 22791 3692 22836 3720
rect 22830 3680 22836 3692
rect 22888 3680 22894 3732
rect 24578 3680 24584 3732
rect 24636 3720 24642 3732
rect 24673 3723 24731 3729
rect 24673 3720 24685 3723
rect 24636 3692 24685 3720
rect 24636 3680 24642 3692
rect 24673 3689 24685 3692
rect 24719 3689 24731 3723
rect 24673 3683 24731 3689
rect 25222 3680 25228 3732
rect 25280 3720 25286 3732
rect 25317 3723 25375 3729
rect 25317 3720 25329 3723
rect 25280 3692 25329 3720
rect 25280 3680 25286 3692
rect 25317 3689 25329 3692
rect 25363 3689 25375 3723
rect 37458 3720 37464 3732
rect 37419 3692 37464 3720
rect 25317 3683 25375 3689
rect 37458 3680 37464 3692
rect 37516 3680 37522 3732
rect 38102 3720 38108 3732
rect 38063 3692 38108 3720
rect 38102 3680 38108 3692
rect 38160 3680 38166 3732
rect 15580 3624 18092 3652
rect 13630 3584 13636 3596
rect 11348 3556 13636 3584
rect 11241 3547 11299 3553
rect 13630 3544 13636 3556
rect 13688 3544 13694 3596
rect 13722 3544 13728 3596
rect 13780 3584 13786 3596
rect 14277 3587 14335 3593
rect 14277 3584 14289 3587
rect 13780 3556 14289 3584
rect 13780 3544 13786 3556
rect 14277 3553 14289 3556
rect 14323 3584 14335 3587
rect 16850 3584 16856 3596
rect 14323 3556 16856 3584
rect 14323 3553 14335 3556
rect 14277 3547 14335 3553
rect 16850 3544 16856 3556
rect 16908 3544 16914 3596
rect 9306 3516 9312 3528
rect 9267 3488 9312 3516
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 9858 3476 9864 3528
rect 9916 3516 9922 3528
rect 9953 3519 10011 3525
rect 9953 3516 9965 3519
rect 9916 3488 9965 3516
rect 9916 3476 9922 3488
rect 9953 3485 9965 3488
rect 9999 3485 10011 3519
rect 9953 3479 10011 3485
rect 10597 3519 10655 3525
rect 10597 3485 10609 3519
rect 10643 3516 10655 3519
rect 10643 3488 11192 3516
rect 10643 3485 10655 3488
rect 10597 3479 10655 3485
rect 11164 3460 11192 3488
rect 13078 3476 13084 3528
rect 13136 3516 13142 3528
rect 13265 3519 13323 3525
rect 13265 3516 13277 3519
rect 13136 3488 13277 3516
rect 13136 3476 13142 3488
rect 13265 3485 13277 3488
rect 13311 3485 13323 3519
rect 13265 3479 13323 3485
rect 13354 3476 13360 3528
rect 13412 3516 13418 3528
rect 18064 3525 18092 3624
rect 18230 3612 18236 3664
rect 18288 3652 18294 3664
rect 18288 3624 21680 3652
rect 18288 3612 18294 3624
rect 21082 3584 21088 3596
rect 18432 3556 21088 3584
rect 18049 3519 18107 3525
rect 13412 3488 14320 3516
rect 13412 3476 13418 3488
rect 7098 3448 7104 3460
rect 7059 3420 7104 3448
rect 7098 3408 7104 3420
rect 7156 3408 7162 3460
rect 9122 3448 9128 3460
rect 8326 3420 9128 3448
rect 9122 3408 9128 3420
rect 9180 3408 9186 3460
rect 9232 3420 10824 3448
rect 7006 3380 7012 3392
rect 6104 3352 7012 3380
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 7190 3340 7196 3392
rect 7248 3380 7254 3392
rect 9232 3380 9260 3420
rect 7248 3352 9260 3380
rect 9401 3383 9459 3389
rect 7248 3340 7254 3352
rect 9401 3349 9413 3383
rect 9447 3380 9459 3383
rect 9674 3380 9680 3392
rect 9447 3352 9680 3380
rect 9447 3349 9459 3352
rect 9401 3343 9459 3349
rect 9674 3340 9680 3352
rect 9732 3340 9738 3392
rect 9766 3340 9772 3392
rect 9824 3380 9830 3392
rect 10134 3380 10140 3392
rect 9824 3352 10140 3380
rect 9824 3340 9830 3352
rect 10134 3340 10140 3352
rect 10192 3340 10198 3392
rect 10226 3340 10232 3392
rect 10284 3380 10290 3392
rect 10689 3383 10747 3389
rect 10689 3380 10701 3383
rect 10284 3352 10701 3380
rect 10284 3340 10290 3352
rect 10689 3349 10701 3352
rect 10735 3349 10747 3383
rect 10796 3380 10824 3420
rect 11146 3408 11152 3460
rect 11204 3408 11210 3460
rect 11422 3408 11428 3460
rect 11480 3448 11486 3460
rect 11517 3451 11575 3457
rect 11517 3448 11529 3451
rect 11480 3420 11529 3448
rect 11480 3408 11486 3420
rect 11517 3417 11529 3420
rect 11563 3417 11575 3451
rect 13538 3448 13544 3460
rect 12742 3420 13544 3448
rect 11517 3411 11575 3417
rect 13538 3408 13544 3420
rect 13596 3408 13602 3460
rect 14292 3448 14320 3488
rect 17512 3488 18000 3516
rect 14553 3451 14611 3457
rect 14553 3448 14565 3451
rect 14292 3420 14565 3448
rect 14553 3417 14565 3420
rect 14599 3448 14611 3451
rect 14826 3448 14832 3460
rect 14599 3420 14832 3448
rect 14599 3417 14611 3420
rect 14553 3411 14611 3417
rect 14826 3408 14832 3420
rect 14884 3408 14890 3460
rect 16390 3448 16396 3460
rect 15778 3420 16396 3448
rect 16390 3408 16396 3420
rect 16448 3408 16454 3460
rect 16574 3448 16580 3460
rect 16535 3420 16580 3448
rect 16574 3408 16580 3420
rect 16632 3408 16638 3460
rect 16669 3451 16727 3457
rect 16669 3417 16681 3451
rect 16715 3448 16727 3451
rect 17512 3448 17540 3488
rect 16715 3420 17540 3448
rect 17589 3451 17647 3457
rect 16715 3417 16727 3420
rect 16669 3411 16727 3417
rect 17589 3417 17601 3451
rect 17635 3448 17647 3451
rect 17770 3448 17776 3460
rect 17635 3420 17776 3448
rect 17635 3417 17647 3420
rect 17589 3411 17647 3417
rect 17770 3408 17776 3420
rect 17828 3408 17834 3460
rect 17972 3448 18000 3488
rect 18049 3485 18061 3519
rect 18095 3485 18107 3519
rect 18049 3479 18107 3485
rect 18432 3448 18460 3556
rect 21082 3544 21088 3556
rect 21140 3544 21146 3596
rect 21652 3584 21680 3624
rect 23382 3612 23388 3664
rect 23440 3652 23446 3664
rect 27246 3652 27252 3664
rect 23440 3624 27252 3652
rect 23440 3612 23446 3624
rect 27246 3612 27252 3624
rect 27304 3612 27310 3664
rect 26605 3587 26663 3593
rect 26605 3584 26617 3587
rect 21652 3556 26617 3584
rect 26605 3553 26617 3556
rect 26651 3553 26663 3587
rect 26605 3547 26663 3553
rect 18690 3516 18696 3528
rect 18651 3488 18696 3516
rect 18690 3476 18696 3488
rect 18748 3476 18754 3528
rect 19429 3519 19487 3525
rect 19429 3485 19441 3519
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 17972 3420 18460 3448
rect 18506 3408 18512 3460
rect 18564 3448 18570 3460
rect 19444 3448 19472 3479
rect 19518 3476 19524 3528
rect 19576 3516 19582 3528
rect 20165 3519 20223 3525
rect 20165 3516 20177 3519
rect 19576 3488 20177 3516
rect 19576 3476 19582 3488
rect 20165 3485 20177 3488
rect 20211 3485 20223 3519
rect 20165 3479 20223 3485
rect 20714 3476 20720 3528
rect 20772 3516 20778 3528
rect 20809 3519 20867 3525
rect 20809 3516 20821 3519
rect 20772 3488 20821 3516
rect 20772 3476 20778 3488
rect 20809 3485 20821 3488
rect 20855 3485 20867 3519
rect 21450 3516 21456 3528
rect 21411 3488 21456 3516
rect 20809 3479 20867 3485
rect 21450 3476 21456 3488
rect 21508 3476 21514 3528
rect 22094 3476 22100 3528
rect 22152 3516 22158 3528
rect 22152 3488 22197 3516
rect 22152 3476 22158 3488
rect 22646 3476 22652 3528
rect 22704 3516 22710 3528
rect 22741 3519 22799 3525
rect 22741 3516 22753 3519
rect 22704 3488 22753 3516
rect 22704 3476 22710 3488
rect 22741 3485 22753 3488
rect 22787 3485 22799 3519
rect 22741 3479 22799 3485
rect 23385 3519 23443 3525
rect 23385 3485 23397 3519
rect 23431 3516 23443 3519
rect 23566 3516 23572 3528
rect 23431 3488 23572 3516
rect 23431 3485 23443 3488
rect 23385 3479 23443 3485
rect 23566 3476 23572 3488
rect 23624 3516 23630 3528
rect 24581 3519 24639 3525
rect 24581 3516 24593 3519
rect 23624 3488 24593 3516
rect 23624 3476 23630 3488
rect 24581 3485 24593 3488
rect 24627 3485 24639 3519
rect 24581 3479 24639 3485
rect 24670 3476 24676 3528
rect 24728 3516 24734 3528
rect 25225 3519 25283 3525
rect 25225 3516 25237 3519
rect 24728 3488 25237 3516
rect 24728 3476 24734 3488
rect 25225 3485 25237 3488
rect 25271 3485 25283 3519
rect 25225 3479 25283 3485
rect 25774 3476 25780 3528
rect 25832 3516 25838 3528
rect 25869 3519 25927 3525
rect 25869 3516 25881 3519
rect 25832 3488 25881 3516
rect 25832 3476 25838 3488
rect 25869 3485 25881 3488
rect 25915 3516 25927 3519
rect 26513 3519 26571 3525
rect 26513 3516 26525 3519
rect 25915 3488 26525 3516
rect 25915 3485 25927 3488
rect 25869 3479 25927 3485
rect 26513 3485 26525 3488
rect 26559 3485 26571 3519
rect 37642 3516 37648 3528
rect 37603 3488 37648 3516
rect 26513 3479 26571 3485
rect 37642 3476 37648 3488
rect 37700 3476 37706 3528
rect 38102 3476 38108 3528
rect 38160 3516 38166 3528
rect 38289 3519 38347 3525
rect 38289 3516 38301 3519
rect 38160 3488 38301 3516
rect 38160 3476 38166 3488
rect 38289 3485 38301 3488
rect 38335 3485 38347 3519
rect 38289 3479 38347 3485
rect 18564 3420 19472 3448
rect 19705 3451 19763 3457
rect 18564 3408 18570 3420
rect 19705 3417 19717 3451
rect 19751 3448 19763 3451
rect 20622 3448 20628 3460
rect 19751 3420 20628 3448
rect 19751 3417 19763 3420
rect 19705 3411 19763 3417
rect 20622 3408 20628 3420
rect 20680 3408 20686 3460
rect 22278 3448 22284 3460
rect 20824 3420 22284 3448
rect 20824 3380 20852 3420
rect 22278 3408 22284 3420
rect 22336 3408 22342 3460
rect 24026 3408 24032 3460
rect 24084 3448 24090 3460
rect 25961 3451 26019 3457
rect 25961 3448 25973 3451
rect 24084 3420 25973 3448
rect 24084 3408 24090 3420
rect 25961 3417 25973 3420
rect 26007 3417 26019 3451
rect 25961 3411 26019 3417
rect 26142 3408 26148 3460
rect 26200 3448 26206 3460
rect 33594 3448 33600 3460
rect 26200 3420 33600 3448
rect 26200 3408 26206 3420
rect 33594 3408 33600 3420
rect 33652 3408 33658 3460
rect 10796 3352 20852 3380
rect 10689 3343 10747 3349
rect 20898 3340 20904 3392
rect 20956 3380 20962 3392
rect 21542 3380 21548 3392
rect 20956 3352 21001 3380
rect 21503 3352 21548 3380
rect 20956 3340 20962 3352
rect 21542 3340 21548 3352
rect 21600 3340 21606 3392
rect 21910 3340 21916 3392
rect 21968 3380 21974 3392
rect 22189 3383 22247 3389
rect 22189 3380 22201 3383
rect 21968 3352 22201 3380
rect 21968 3340 21974 3352
rect 22189 3349 22201 3352
rect 22235 3349 22247 3383
rect 22189 3343 22247 3349
rect 23477 3383 23535 3389
rect 23477 3349 23489 3383
rect 23523 3380 23535 3383
rect 23566 3380 23572 3392
rect 23523 3352 23572 3380
rect 23523 3349 23535 3352
rect 23477 3343 23535 3349
rect 23566 3340 23572 3352
rect 23624 3340 23630 3392
rect 24394 3340 24400 3392
rect 24452 3380 24458 3392
rect 26234 3380 26240 3392
rect 24452 3352 26240 3380
rect 24452 3340 24458 3352
rect 26234 3340 26240 3352
rect 26292 3340 26298 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 3418 3176 3424 3188
rect 3379 3148 3424 3176
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 4706 3136 4712 3188
rect 4764 3176 4770 3188
rect 5445 3179 5503 3185
rect 5445 3176 5457 3179
rect 4764 3148 5457 3176
rect 4764 3136 4770 3148
rect 5445 3145 5457 3148
rect 5491 3145 5503 3179
rect 5445 3139 5503 3145
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 20806 3176 20812 3188
rect 5592 3148 15700 3176
rect 5592 3136 5598 3148
rect 1946 3068 1952 3120
rect 2004 3108 2010 3120
rect 3786 3108 3792 3120
rect 2004 3080 3792 3108
rect 2004 3068 2010 3080
rect 3786 3068 3792 3080
rect 3844 3068 3850 3120
rect 4154 3068 4160 3120
rect 4212 3108 4218 3120
rect 5350 3108 5356 3120
rect 4212 3080 5356 3108
rect 4212 3068 4218 3080
rect 5350 3068 5356 3080
rect 5408 3068 5414 3120
rect 8110 3108 8116 3120
rect 5460 3080 8116 3108
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3040 1639 3043
rect 2498 3040 2504 3052
rect 1627 3012 2504 3040
rect 1627 3009 1639 3012
rect 1581 3003 1639 3009
rect 2498 3000 2504 3012
rect 2556 3000 2562 3052
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3009 2927 3043
rect 2869 3003 2927 3009
rect 3329 3043 3387 3049
rect 3329 3009 3341 3043
rect 3375 3040 3387 3043
rect 3694 3040 3700 3052
rect 3375 3012 3700 3040
rect 3375 3009 3387 3012
rect 3329 3003 3387 3009
rect 2884 2972 2912 3003
rect 3694 3000 3700 3012
rect 3752 3000 3758 3052
rect 3970 3040 3976 3052
rect 3931 3012 3976 3040
rect 3970 3000 3976 3012
rect 4028 3000 4034 3052
rect 4617 3043 4675 3049
rect 4617 3009 4629 3043
rect 4663 3009 4675 3043
rect 4617 3003 4675 3009
rect 4632 2972 4660 3003
rect 4982 3000 4988 3052
rect 5040 3040 5046 3052
rect 5166 3040 5172 3052
rect 5040 3012 5172 3040
rect 5040 3000 5046 3012
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 5460 3049 5488 3080
rect 8110 3068 8116 3080
rect 8168 3068 8174 3120
rect 9490 3108 9496 3120
rect 8220 3080 9496 3108
rect 5445 3043 5503 3049
rect 5445 3009 5457 3043
rect 5491 3009 5503 3043
rect 5445 3003 5503 3009
rect 7009 3043 7067 3049
rect 7009 3009 7021 3043
rect 7055 3040 7067 3043
rect 7558 3040 7564 3052
rect 7055 3012 7564 3040
rect 7055 3009 7067 3012
rect 7009 3003 7067 3009
rect 7558 3000 7564 3012
rect 7616 3040 7622 3052
rect 7653 3043 7711 3049
rect 7653 3040 7665 3043
rect 7616 3012 7665 3040
rect 7616 3000 7622 3012
rect 7653 3009 7665 3012
rect 7699 3009 7711 3043
rect 7653 3003 7711 3009
rect 7742 3000 7748 3052
rect 7800 3040 7806 3052
rect 7800 3012 7845 3040
rect 7800 3000 7806 3012
rect 6914 2972 6920 2984
rect 2884 2944 4568 2972
rect 4632 2944 6920 2972
rect 4062 2904 4068 2916
rect 4023 2876 4068 2904
rect 4062 2864 4068 2876
rect 4120 2864 4126 2916
rect 4540 2904 4568 2944
rect 6914 2932 6920 2944
rect 6972 2932 6978 2984
rect 8220 2972 8248 3080
rect 9490 3068 9496 3080
rect 9548 3068 9554 3120
rect 9674 3068 9680 3120
rect 9732 3068 9738 3120
rect 10686 3068 10692 3120
rect 10744 3108 10750 3120
rect 12253 3111 12311 3117
rect 12253 3108 12265 3111
rect 10744 3080 12265 3108
rect 10744 3068 10750 3080
rect 12253 3077 12265 3080
rect 12299 3077 12311 3111
rect 13354 3108 13360 3120
rect 12253 3071 12311 3077
rect 13188 3080 13360 3108
rect 8297 3043 8355 3049
rect 8297 3009 8309 3043
rect 8343 3009 8355 3043
rect 8297 3003 8355 3009
rect 7024 2944 8248 2972
rect 8312 2972 8340 3003
rect 8386 3000 8392 3052
rect 8444 3040 8450 3052
rect 8941 3043 8999 3049
rect 8941 3040 8953 3043
rect 8444 3012 8953 3040
rect 8444 3000 8450 3012
rect 8941 3009 8953 3012
rect 8987 3009 8999 3043
rect 8941 3003 8999 3009
rect 11146 3000 11152 3052
rect 11204 3040 11210 3052
rect 11882 3040 11888 3052
rect 11204 3012 11888 3040
rect 11204 3000 11210 3012
rect 11882 3000 11888 3012
rect 11940 3040 11946 3052
rect 12158 3040 12164 3052
rect 11940 3012 12164 3040
rect 11940 3000 11946 3012
rect 12158 3000 12164 3012
rect 12216 3000 12222 3052
rect 13188 3049 13216 3080
rect 13354 3068 13360 3080
rect 13412 3068 13418 3120
rect 13446 3068 13452 3120
rect 13504 3108 13510 3120
rect 15470 3108 15476 3120
rect 13504 3080 13549 3108
rect 14674 3080 15476 3108
rect 13504 3068 13510 3080
rect 15470 3068 15476 3080
rect 15528 3068 15534 3120
rect 15672 3117 15700 3148
rect 15764 3148 20812 3176
rect 15764 3117 15792 3148
rect 20806 3136 20812 3148
rect 20864 3136 20870 3188
rect 22002 3176 22008 3188
rect 20916 3148 22008 3176
rect 15657 3111 15715 3117
rect 15657 3077 15669 3111
rect 15703 3077 15715 3111
rect 15657 3071 15715 3077
rect 15749 3111 15807 3117
rect 15749 3077 15761 3111
rect 15795 3077 15807 3111
rect 15749 3071 15807 3077
rect 16574 3068 16580 3120
rect 16632 3108 16638 3120
rect 17037 3111 17095 3117
rect 17037 3108 17049 3111
rect 16632 3080 17049 3108
rect 16632 3068 16638 3080
rect 17037 3077 17049 3080
rect 17083 3077 17095 3111
rect 17037 3071 17095 3077
rect 17678 3068 17684 3120
rect 17736 3108 17742 3120
rect 18141 3111 18199 3117
rect 18141 3108 18153 3111
rect 17736 3080 18153 3108
rect 17736 3068 17742 3080
rect 18141 3077 18153 3080
rect 18187 3077 18199 3111
rect 18141 3071 18199 3077
rect 18877 3111 18935 3117
rect 18877 3077 18889 3111
rect 18923 3108 18935 3111
rect 19978 3108 19984 3120
rect 18923 3080 19984 3108
rect 18923 3077 18935 3080
rect 18877 3071 18935 3077
rect 19978 3068 19984 3080
rect 20036 3068 20042 3120
rect 20070 3068 20076 3120
rect 20128 3108 20134 3120
rect 20349 3111 20407 3117
rect 20349 3108 20361 3111
rect 20128 3080 20361 3108
rect 20128 3068 20134 3080
rect 20349 3077 20361 3080
rect 20395 3077 20407 3111
rect 20349 3071 20407 3077
rect 20441 3111 20499 3117
rect 20441 3077 20453 3111
rect 20487 3108 20499 3111
rect 20622 3108 20628 3120
rect 20487 3080 20628 3108
rect 20487 3077 20499 3080
rect 20441 3071 20499 3077
rect 20622 3068 20628 3080
rect 20680 3068 20686 3120
rect 20714 3068 20720 3120
rect 20772 3108 20778 3120
rect 20916 3108 20944 3148
rect 22002 3136 22008 3148
rect 22060 3136 22066 3188
rect 22646 3176 22652 3188
rect 22607 3148 22652 3176
rect 22646 3136 22652 3148
rect 22704 3136 22710 3188
rect 22756 3148 25912 3176
rect 20772 3080 20944 3108
rect 20993 3111 21051 3117
rect 20772 3068 20778 3080
rect 20993 3077 21005 3111
rect 21039 3108 21051 3111
rect 22756 3108 22784 3148
rect 21039 3080 22784 3108
rect 21039 3077 21051 3080
rect 20993 3071 21051 3077
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3009 13231 3043
rect 13173 3003 13231 3009
rect 16301 3043 16359 3049
rect 16301 3009 16313 3043
rect 16347 3040 16359 3043
rect 16666 3040 16672 3052
rect 16347 3012 16672 3040
rect 16347 3009 16359 3012
rect 16301 3003 16359 3009
rect 16666 3000 16672 3012
rect 16724 3000 16730 3052
rect 18046 3040 18052 3052
rect 18007 3012 18052 3040
rect 18046 3000 18052 3012
rect 18104 3000 18110 3052
rect 8662 2972 8668 2984
rect 8312 2944 8668 2972
rect 7024 2904 7052 2944
rect 8662 2932 8668 2944
rect 8720 2932 8726 2984
rect 9217 2975 9275 2981
rect 9217 2941 9229 2975
rect 9263 2972 9275 2975
rect 9950 2972 9956 2984
rect 9263 2944 9956 2972
rect 9263 2941 9275 2944
rect 9217 2935 9275 2941
rect 9950 2932 9956 2944
rect 10008 2932 10014 2984
rect 13998 2972 14004 2984
rect 10244 2944 14004 2972
rect 4540 2876 7052 2904
rect 7101 2907 7159 2913
rect 7101 2873 7113 2907
rect 7147 2904 7159 2907
rect 7147 2876 9076 2904
rect 7147 2873 7159 2876
rect 7101 2867 7159 2873
rect 658 2796 664 2848
rect 716 2836 722 2848
rect 1765 2839 1823 2845
rect 1765 2836 1777 2839
rect 716 2808 1777 2836
rect 716 2796 722 2808
rect 1765 2805 1777 2808
rect 1811 2805 1823 2839
rect 2682 2836 2688 2848
rect 2643 2808 2688 2836
rect 1765 2799 1823 2805
rect 2682 2796 2688 2808
rect 2740 2796 2746 2848
rect 4709 2839 4767 2845
rect 4709 2805 4721 2839
rect 4755 2836 4767 2839
rect 5994 2836 6000 2848
rect 4755 2808 6000 2836
rect 4755 2805 4767 2808
rect 4709 2799 4767 2805
rect 5994 2796 6000 2808
rect 6052 2796 6058 2848
rect 8389 2839 8447 2845
rect 8389 2805 8401 2839
rect 8435 2836 8447 2839
rect 8478 2836 8484 2848
rect 8435 2808 8484 2836
rect 8435 2805 8447 2808
rect 8389 2799 8447 2805
rect 8478 2796 8484 2808
rect 8536 2796 8542 2848
rect 9048 2836 9076 2876
rect 10244 2836 10272 2944
rect 13998 2932 14004 2944
rect 14056 2932 14062 2984
rect 16945 2975 17003 2981
rect 16945 2972 16957 2975
rect 15580 2944 16957 2972
rect 10318 2864 10324 2916
rect 10376 2904 10382 2916
rect 10689 2907 10747 2913
rect 10689 2904 10701 2907
rect 10376 2876 10701 2904
rect 10376 2864 10382 2876
rect 10689 2873 10701 2876
rect 10735 2873 10747 2907
rect 15580 2904 15608 2944
rect 16945 2941 16957 2944
rect 16991 2941 17003 2975
rect 16945 2935 17003 2941
rect 17221 2975 17279 2981
rect 17221 2941 17233 2975
rect 17267 2972 17279 2975
rect 18598 2972 18604 2984
rect 17267 2944 18604 2972
rect 17267 2941 17279 2944
rect 17221 2935 17279 2941
rect 10689 2867 10747 2873
rect 14476 2876 15608 2904
rect 9048 2808 10272 2836
rect 11606 2796 11612 2848
rect 11664 2836 11670 2848
rect 14476 2836 14504 2876
rect 16298 2864 16304 2916
rect 16356 2904 16362 2916
rect 17236 2904 17264 2935
rect 18598 2932 18604 2944
rect 18656 2932 18662 2984
rect 18782 2972 18788 2984
rect 18743 2944 18788 2972
rect 18782 2932 18788 2944
rect 18840 2932 18846 2984
rect 18874 2932 18880 2984
rect 18932 2972 18938 2984
rect 19061 2975 19119 2981
rect 19061 2972 19073 2975
rect 18932 2944 19073 2972
rect 18932 2932 18938 2944
rect 19061 2941 19073 2944
rect 19107 2941 19119 2975
rect 19061 2935 19119 2941
rect 19242 2932 19248 2984
rect 19300 2972 19306 2984
rect 21008 2972 21036 3071
rect 22189 3043 22247 3049
rect 22189 3009 22201 3043
rect 22235 3040 22247 3043
rect 22462 3040 22468 3052
rect 22235 3012 22468 3040
rect 22235 3009 22247 3012
rect 22189 3003 22247 3009
rect 22462 3000 22468 3012
rect 22520 3000 22526 3052
rect 22833 3043 22891 3049
rect 22833 3009 22845 3043
rect 22879 3009 22891 3043
rect 22833 3003 22891 3009
rect 19300 2944 21036 2972
rect 19300 2932 19306 2944
rect 21910 2932 21916 2984
rect 21968 2972 21974 2984
rect 22848 2972 22876 3003
rect 23198 3000 23204 3052
rect 23256 3040 23262 3052
rect 23293 3043 23351 3049
rect 23293 3040 23305 3043
rect 23256 3012 23305 3040
rect 23256 3000 23262 3012
rect 23293 3009 23305 3012
rect 23339 3040 23351 3043
rect 23937 3043 23995 3049
rect 23937 3040 23949 3043
rect 23339 3012 23949 3040
rect 23339 3009 23351 3012
rect 23293 3003 23351 3009
rect 23937 3009 23949 3012
rect 23983 3040 23995 3043
rect 24578 3040 24584 3052
rect 23983 3012 24584 3040
rect 23983 3009 23995 3012
rect 23937 3003 23995 3009
rect 24578 3000 24584 3012
rect 24636 3000 24642 3052
rect 24765 3043 24823 3049
rect 24765 3009 24777 3043
rect 24811 3009 24823 3043
rect 25406 3040 25412 3052
rect 25367 3012 25412 3040
rect 24765 3003 24823 3009
rect 21968 2944 22876 2972
rect 21968 2932 21974 2944
rect 22922 2932 22928 2984
rect 22980 2972 22986 2984
rect 24780 2972 24808 3003
rect 25406 3000 25412 3012
rect 25464 3000 25470 3052
rect 25884 3049 25912 3148
rect 27154 3136 27160 3188
rect 27212 3176 27218 3188
rect 37461 3179 37519 3185
rect 37461 3176 37473 3179
rect 27212 3148 37473 3176
rect 27212 3136 27218 3148
rect 37461 3145 37473 3148
rect 37507 3145 37519 3179
rect 37461 3139 37519 3145
rect 27246 3108 27252 3120
rect 27207 3080 27252 3108
rect 27246 3068 27252 3080
rect 27304 3068 27310 3120
rect 36722 3068 36728 3120
rect 36780 3108 36786 3120
rect 36780 3080 37688 3108
rect 36780 3068 36786 3080
rect 25869 3043 25927 3049
rect 25869 3009 25881 3043
rect 25915 3009 25927 3043
rect 25869 3003 25927 3009
rect 26234 3000 26240 3052
rect 26292 3040 26298 3052
rect 27157 3043 27215 3049
rect 27157 3040 27169 3043
rect 26292 3012 27169 3040
rect 26292 3000 26298 3012
rect 27157 3009 27169 3012
rect 27203 3009 27215 3043
rect 33594 3040 33600 3052
rect 33555 3012 33600 3040
rect 27157 3003 27215 3009
rect 33594 3000 33600 3012
rect 33652 3000 33658 3052
rect 36906 3040 36912 3052
rect 36867 3012 36912 3040
rect 36906 3000 36912 3012
rect 36964 3000 36970 3052
rect 37660 3049 37688 3080
rect 37645 3043 37703 3049
rect 37645 3009 37657 3043
rect 37691 3009 37703 3043
rect 38286 3040 38292 3052
rect 38247 3012 38292 3040
rect 37645 3003 37703 3009
rect 38286 3000 38292 3012
rect 38344 3000 38350 3052
rect 25961 2975 26019 2981
rect 25961 2972 25973 2975
rect 22980 2944 24716 2972
rect 24780 2944 25973 2972
rect 22980 2932 22986 2944
rect 16356 2876 17264 2904
rect 16356 2864 16362 2876
rect 17586 2864 17592 2916
rect 17644 2904 17650 2916
rect 20254 2904 20260 2916
rect 17644 2876 20260 2904
rect 17644 2864 17650 2876
rect 20254 2864 20260 2876
rect 20312 2864 20318 2916
rect 22005 2907 22063 2913
rect 22005 2873 22017 2907
rect 22051 2904 22063 2907
rect 22646 2904 22652 2916
rect 22051 2876 22652 2904
rect 22051 2873 22063 2876
rect 22005 2867 22063 2873
rect 22646 2864 22652 2876
rect 22704 2864 22710 2916
rect 22738 2864 22744 2916
rect 22796 2904 22802 2916
rect 24581 2907 24639 2913
rect 24581 2904 24593 2907
rect 22796 2876 24593 2904
rect 22796 2864 22802 2876
rect 24581 2873 24593 2876
rect 24627 2873 24639 2907
rect 24688 2904 24716 2944
rect 25961 2941 25973 2944
rect 26007 2941 26019 2975
rect 25961 2935 26019 2941
rect 30742 2932 30748 2984
rect 30800 2972 30806 2984
rect 30800 2944 38148 2972
rect 30800 2932 30806 2944
rect 25866 2904 25872 2916
rect 24688 2876 25872 2904
rect 24581 2867 24639 2873
rect 25866 2864 25872 2876
rect 25924 2864 25930 2916
rect 30558 2864 30564 2916
rect 30616 2904 30622 2916
rect 38120 2913 38148 2944
rect 36725 2907 36783 2913
rect 36725 2904 36737 2907
rect 30616 2876 36737 2904
rect 30616 2864 30622 2876
rect 36725 2873 36737 2876
rect 36771 2873 36783 2907
rect 36725 2867 36783 2873
rect 38105 2907 38163 2913
rect 38105 2873 38117 2907
rect 38151 2873 38163 2907
rect 38105 2867 38163 2873
rect 11664 2808 14504 2836
rect 14921 2839 14979 2845
rect 11664 2796 11670 2808
rect 14921 2805 14933 2839
rect 14967 2836 14979 2839
rect 15102 2836 15108 2848
rect 14967 2808 15108 2836
rect 14967 2805 14979 2808
rect 14921 2799 14979 2805
rect 15102 2796 15108 2808
rect 15160 2796 15166 2848
rect 17954 2796 17960 2848
rect 18012 2836 18018 2848
rect 21266 2836 21272 2848
rect 18012 2808 21272 2836
rect 18012 2796 18018 2808
rect 21266 2796 21272 2808
rect 21324 2796 21330 2848
rect 22094 2796 22100 2848
rect 22152 2836 22158 2848
rect 23385 2839 23443 2845
rect 23385 2836 23397 2839
rect 22152 2808 23397 2836
rect 22152 2796 22158 2808
rect 23385 2805 23397 2808
rect 23431 2805 23443 2839
rect 23385 2799 23443 2805
rect 23474 2796 23480 2848
rect 23532 2836 23538 2848
rect 24029 2839 24087 2845
rect 24029 2836 24041 2839
rect 23532 2808 24041 2836
rect 23532 2796 23538 2808
rect 24029 2805 24041 2808
rect 24075 2805 24087 2839
rect 24029 2799 24087 2805
rect 24486 2796 24492 2848
rect 24544 2836 24550 2848
rect 25225 2839 25283 2845
rect 25225 2836 25237 2839
rect 24544 2808 25237 2836
rect 24544 2796 24550 2808
rect 25225 2805 25237 2808
rect 25271 2805 25283 2839
rect 25225 2799 25283 2805
rect 33502 2796 33508 2848
rect 33560 2836 33566 2848
rect 33781 2839 33839 2845
rect 33781 2836 33793 2839
rect 33560 2808 33793 2836
rect 33560 2796 33566 2808
rect 33781 2805 33793 2808
rect 33827 2805 33839 2839
rect 33781 2799 33839 2805
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 1486 2592 1492 2644
rect 1544 2632 1550 2644
rect 1765 2635 1823 2641
rect 1765 2632 1777 2635
rect 1544 2604 1777 2632
rect 1544 2592 1550 2604
rect 1765 2601 1777 2604
rect 1811 2601 1823 2635
rect 1765 2595 1823 2601
rect 9122 2592 9128 2644
rect 9180 2632 9186 2644
rect 10321 2635 10379 2641
rect 10321 2632 10333 2635
rect 9180 2604 10333 2632
rect 9180 2592 9186 2604
rect 10321 2601 10333 2604
rect 10367 2601 10379 2635
rect 10321 2595 10379 2601
rect 11238 2592 11244 2644
rect 11296 2632 11302 2644
rect 11885 2635 11943 2641
rect 11885 2632 11897 2635
rect 11296 2604 11897 2632
rect 11296 2592 11302 2604
rect 11885 2601 11897 2604
rect 11931 2601 11943 2635
rect 11885 2595 11943 2601
rect 11974 2592 11980 2644
rect 12032 2632 12038 2644
rect 14540 2635 14598 2641
rect 12032 2604 14412 2632
rect 12032 2592 12038 2604
rect 14 2524 20 2576
rect 72 2564 78 2576
rect 3237 2567 3295 2573
rect 3237 2564 3249 2567
rect 72 2536 3249 2564
rect 72 2524 78 2536
rect 3237 2533 3249 2536
rect 3283 2533 3295 2567
rect 3237 2527 3295 2533
rect 7742 2524 7748 2576
rect 7800 2564 7806 2576
rect 9306 2564 9312 2576
rect 7800 2536 9312 2564
rect 7800 2524 7806 2536
rect 9306 2524 9312 2536
rect 9364 2524 9370 2576
rect 9677 2567 9735 2573
rect 9677 2533 9689 2567
rect 9723 2564 9735 2567
rect 11054 2564 11060 2576
rect 9723 2536 11060 2564
rect 9723 2533 9735 2536
rect 9677 2527 9735 2533
rect 11054 2524 11060 2536
rect 11112 2524 11118 2576
rect 13906 2564 13912 2576
rect 12820 2536 13912 2564
rect 5626 2496 5632 2508
rect 4172 2468 5632 2496
rect 2222 2388 2228 2440
rect 2280 2428 2286 2440
rect 2317 2431 2375 2437
rect 2317 2428 2329 2431
rect 2280 2400 2329 2428
rect 2280 2388 2286 2400
rect 2317 2397 2329 2400
rect 2363 2397 2375 2431
rect 3050 2428 3056 2440
rect 3011 2400 3056 2428
rect 2317 2391 2375 2397
rect 3050 2388 3056 2400
rect 3108 2388 3114 2440
rect 4172 2437 4200 2468
rect 5626 2456 5632 2468
rect 5684 2456 5690 2508
rect 6914 2456 6920 2508
rect 6972 2496 6978 2508
rect 9324 2496 9352 2524
rect 6972 2468 8294 2496
rect 9324 2468 9620 2496
rect 6972 2456 6978 2468
rect 4157 2431 4215 2437
rect 4157 2397 4169 2431
rect 4203 2397 4215 2431
rect 4614 2428 4620 2440
rect 4575 2400 4620 2428
rect 4157 2391 4215 2397
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 5258 2428 5264 2440
rect 5219 2400 5264 2428
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 7101 2431 7159 2437
rect 7101 2397 7113 2431
rect 7147 2428 7159 2431
rect 7742 2428 7748 2440
rect 7147 2400 7748 2428
rect 7147 2397 7159 2400
rect 7101 2391 7159 2397
rect 7742 2388 7748 2400
rect 7800 2388 7806 2440
rect 8266 2428 8294 2468
rect 9592 2439 9620 2468
rect 8389 2431 8447 2437
rect 8389 2428 8401 2431
rect 8266 2400 8401 2428
rect 8389 2397 8401 2400
rect 8435 2428 8447 2431
rect 9577 2433 9635 2439
rect 8435 2400 9536 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 1670 2360 1676 2372
rect 1631 2332 1676 2360
rect 1670 2320 1676 2332
rect 1728 2320 1734 2372
rect 7193 2363 7251 2369
rect 7193 2329 7205 2363
rect 7239 2360 7251 2363
rect 9398 2360 9404 2372
rect 7239 2332 9404 2360
rect 7239 2329 7251 2332
rect 7193 2323 7251 2329
rect 9398 2320 9404 2332
rect 9456 2320 9462 2372
rect 2498 2292 2504 2304
rect 2459 2264 2504 2292
rect 2498 2252 2504 2264
rect 2556 2252 2562 2304
rect 3970 2292 3976 2304
rect 3931 2264 3976 2292
rect 3970 2252 3976 2264
rect 4028 2252 4034 2304
rect 4706 2292 4712 2304
rect 4667 2264 4712 2292
rect 4706 2252 4712 2264
rect 4764 2252 4770 2304
rect 5166 2252 5172 2304
rect 5224 2292 5230 2304
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 5224 2264 5457 2292
rect 5224 2252 5230 2264
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 7834 2292 7840 2304
rect 7795 2264 7840 2292
rect 5445 2255 5503 2261
rect 7834 2252 7840 2264
rect 7892 2252 7898 2304
rect 8478 2292 8484 2304
rect 8439 2264 8484 2292
rect 8478 2252 8484 2264
rect 8536 2252 8542 2304
rect 9508 2292 9536 2400
rect 9577 2399 9589 2433
rect 9623 2399 9635 2433
rect 9577 2393 9635 2399
rect 10134 2388 10140 2440
rect 10192 2428 10198 2440
rect 10229 2431 10287 2437
rect 10229 2428 10241 2431
rect 10192 2400 10241 2428
rect 10192 2388 10198 2400
rect 10229 2397 10241 2400
rect 10275 2397 10287 2431
rect 10870 2428 10876 2440
rect 10831 2400 10876 2428
rect 10229 2391 10287 2397
rect 10870 2388 10876 2400
rect 10928 2388 10934 2440
rect 12820 2437 12848 2536
rect 13906 2524 13912 2536
rect 13964 2524 13970 2576
rect 13722 2456 13728 2508
rect 13780 2496 13786 2508
rect 14277 2499 14335 2505
rect 14277 2496 14289 2499
rect 13780 2468 14289 2496
rect 13780 2456 13786 2468
rect 14277 2465 14289 2468
rect 14323 2465 14335 2499
rect 14384 2496 14412 2604
rect 14540 2601 14552 2635
rect 14586 2632 14598 2635
rect 15930 2632 15936 2644
rect 14586 2604 15936 2632
rect 14586 2601 14598 2604
rect 14540 2595 14598 2601
rect 15930 2592 15936 2604
rect 15988 2592 15994 2644
rect 16025 2635 16083 2641
rect 16025 2601 16037 2635
rect 16071 2632 16083 2635
rect 16758 2632 16764 2644
rect 16071 2604 16764 2632
rect 16071 2601 16083 2604
rect 16025 2595 16083 2601
rect 16758 2592 16764 2604
rect 16816 2592 16822 2644
rect 16945 2635 17003 2641
rect 16945 2601 16957 2635
rect 16991 2632 17003 2635
rect 17310 2632 17316 2644
rect 16991 2604 17316 2632
rect 16991 2601 17003 2604
rect 16945 2595 17003 2601
rect 17310 2592 17316 2604
rect 17368 2592 17374 2644
rect 17402 2592 17408 2644
rect 17460 2632 17466 2644
rect 19521 2635 19579 2641
rect 19521 2632 19533 2635
rect 17460 2604 19533 2632
rect 17460 2592 17466 2604
rect 19521 2601 19533 2604
rect 19567 2601 19579 2635
rect 19521 2595 19579 2601
rect 20162 2592 20168 2644
rect 20220 2632 20226 2644
rect 20441 2635 20499 2641
rect 20441 2632 20453 2635
rect 20220 2604 20453 2632
rect 20220 2592 20226 2604
rect 20441 2601 20453 2604
rect 20487 2601 20499 2635
rect 20441 2595 20499 2601
rect 21177 2635 21235 2641
rect 21177 2601 21189 2635
rect 21223 2632 21235 2635
rect 21358 2632 21364 2644
rect 21223 2604 21364 2632
rect 21223 2601 21235 2604
rect 21177 2595 21235 2601
rect 21358 2592 21364 2604
rect 21416 2592 21422 2644
rect 22005 2635 22063 2641
rect 22005 2601 22017 2635
rect 22051 2632 22063 2635
rect 25222 2632 25228 2644
rect 22051 2604 25228 2632
rect 22051 2601 22063 2604
rect 22005 2595 22063 2601
rect 25222 2592 25228 2604
rect 25280 2592 25286 2644
rect 27798 2632 27804 2644
rect 27759 2604 27804 2632
rect 27798 2592 27804 2604
rect 27856 2592 27862 2644
rect 28626 2632 28632 2644
rect 28587 2604 28632 2632
rect 28626 2592 28632 2604
rect 28684 2592 28690 2644
rect 30098 2592 30104 2644
rect 30156 2632 30162 2644
rect 30469 2635 30527 2641
rect 30469 2632 30481 2635
rect 30156 2604 30481 2632
rect 30156 2592 30162 2604
rect 30469 2601 30481 2604
rect 30515 2601 30527 2635
rect 30469 2595 30527 2601
rect 16114 2524 16120 2576
rect 16172 2564 16178 2576
rect 18417 2567 18475 2573
rect 18417 2564 18429 2567
rect 16172 2536 18429 2564
rect 16172 2524 16178 2536
rect 18417 2533 18429 2536
rect 18463 2533 18475 2567
rect 22738 2564 22744 2576
rect 18417 2527 18475 2533
rect 19812 2536 22744 2564
rect 16574 2496 16580 2508
rect 14384 2468 16580 2496
rect 14277 2459 14335 2465
rect 16574 2456 16580 2468
rect 16632 2456 16638 2508
rect 19812 2496 19840 2536
rect 22738 2524 22744 2536
rect 22796 2524 22802 2576
rect 23382 2564 23388 2576
rect 23343 2536 23388 2564
rect 23382 2524 23388 2536
rect 23440 2524 23446 2576
rect 27430 2524 27436 2576
rect 27488 2564 27494 2576
rect 27488 2536 35894 2564
rect 27488 2524 27494 2536
rect 17512 2468 19840 2496
rect 20257 2499 20315 2505
rect 12805 2431 12863 2437
rect 12805 2397 12817 2431
rect 12851 2397 12863 2431
rect 13446 2428 13452 2440
rect 13407 2400 13452 2428
rect 12805 2391 12863 2397
rect 13446 2388 13452 2400
rect 13504 2388 13510 2440
rect 17512 2437 17540 2468
rect 20257 2465 20269 2499
rect 20303 2496 20315 2499
rect 21542 2496 21548 2508
rect 20303 2468 21548 2496
rect 20303 2465 20315 2468
rect 20257 2459 20315 2465
rect 21542 2456 21548 2468
rect 21600 2456 21606 2508
rect 21652 2468 23612 2496
rect 16853 2431 16911 2437
rect 16853 2397 16865 2431
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 17497 2431 17555 2437
rect 17497 2397 17509 2431
rect 17543 2397 17555 2431
rect 18230 2428 18236 2440
rect 18191 2400 18236 2428
rect 17497 2391 17555 2397
rect 11514 2360 11520 2372
rect 9646 2332 11520 2360
rect 9646 2292 9674 2332
rect 11514 2320 11520 2332
rect 11572 2320 11578 2372
rect 11606 2320 11612 2372
rect 11664 2360 11670 2372
rect 11793 2363 11851 2369
rect 11793 2360 11805 2363
rect 11664 2332 11805 2360
rect 11664 2320 11670 2332
rect 11793 2329 11805 2332
rect 11839 2329 11851 2363
rect 11793 2323 11851 2329
rect 12158 2320 12164 2372
rect 12216 2360 12222 2372
rect 16758 2360 16764 2372
rect 12216 2332 14964 2360
rect 15778 2332 16764 2360
rect 12216 2320 12222 2332
rect 9508 2264 9674 2292
rect 10962 2252 10968 2304
rect 11020 2292 11026 2304
rect 11057 2295 11115 2301
rect 11057 2292 11069 2295
rect 11020 2264 11069 2292
rect 11020 2252 11026 2264
rect 11057 2261 11069 2264
rect 11103 2261 11115 2295
rect 11057 2255 11115 2261
rect 12897 2295 12955 2301
rect 12897 2261 12909 2295
rect 12943 2292 12955 2295
rect 13538 2292 13544 2304
rect 12943 2264 13544 2292
rect 12943 2261 12955 2264
rect 12897 2255 12955 2261
rect 13538 2252 13544 2264
rect 13596 2252 13602 2304
rect 13633 2295 13691 2301
rect 13633 2261 13645 2295
rect 13679 2292 13691 2295
rect 14826 2292 14832 2304
rect 13679 2264 14832 2292
rect 13679 2261 13691 2264
rect 13633 2255 13691 2261
rect 14826 2252 14832 2264
rect 14884 2252 14890 2304
rect 14936 2292 14964 2332
rect 16758 2320 16764 2332
rect 16816 2320 16822 2372
rect 16868 2360 16896 2391
rect 18230 2388 18236 2400
rect 18288 2388 18294 2440
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 18340 2400 19441 2428
rect 18340 2360 18368 2400
rect 16868 2332 18368 2360
rect 16868 2292 16896 2332
rect 14936 2264 16896 2292
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17460 2264 17693 2292
rect 17460 2252 17466 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 19260 2292 19288 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 20070 2428 20076 2440
rect 20031 2400 20076 2428
rect 19429 2391 19487 2397
rect 20070 2388 20076 2400
rect 20128 2388 20134 2440
rect 20622 2388 20628 2440
rect 20680 2428 20686 2440
rect 21361 2431 21419 2437
rect 21361 2428 21373 2431
rect 20680 2400 21373 2428
rect 20680 2388 20686 2400
rect 21361 2397 21373 2400
rect 21407 2397 21419 2431
rect 21361 2391 21419 2397
rect 19334 2320 19340 2372
rect 19392 2360 19398 2372
rect 21652 2360 21680 2468
rect 22002 2388 22008 2440
rect 22060 2428 22066 2440
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 22060 2400 22201 2428
rect 22060 2388 22066 2400
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22646 2428 22652 2440
rect 22607 2400 22652 2428
rect 22189 2391 22247 2397
rect 22646 2388 22652 2400
rect 22704 2388 22710 2440
rect 23584 2437 23612 2468
rect 24118 2456 24124 2508
rect 24176 2496 24182 2508
rect 32585 2499 32643 2505
rect 32585 2496 32597 2499
rect 24176 2468 32597 2496
rect 24176 2456 24182 2468
rect 32585 2465 32597 2468
rect 32631 2465 32643 2499
rect 32585 2459 32643 2465
rect 23569 2431 23627 2437
rect 23569 2397 23581 2431
rect 23615 2397 23627 2431
rect 24578 2428 24584 2440
rect 24539 2400 24584 2428
rect 23569 2391 23627 2397
rect 24578 2388 24584 2400
rect 24636 2388 24642 2440
rect 25222 2428 25228 2440
rect 25183 2400 25228 2428
rect 25222 2388 25228 2400
rect 25280 2388 25286 2440
rect 25866 2388 25872 2440
rect 25924 2428 25930 2440
rect 25961 2431 26019 2437
rect 25961 2428 25973 2431
rect 25924 2400 25973 2428
rect 25924 2388 25930 2400
rect 25961 2397 25973 2400
rect 26007 2397 26019 2431
rect 27338 2428 27344 2440
rect 27299 2400 27344 2428
rect 25961 2391 26019 2397
rect 27338 2388 27344 2400
rect 27396 2388 27402 2440
rect 27985 2431 28043 2437
rect 27985 2397 27997 2431
rect 28031 2397 28043 2431
rect 27985 2391 28043 2397
rect 19392 2332 21680 2360
rect 19392 2320 19398 2332
rect 27062 2320 27068 2372
rect 27120 2360 27126 2372
rect 28000 2360 28028 2391
rect 29454 2388 29460 2440
rect 29512 2428 29518 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29512 2400 29745 2428
rect 29512 2388 29518 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 30282 2388 30288 2440
rect 30340 2428 30346 2440
rect 30653 2431 30711 2437
rect 30653 2428 30665 2431
rect 30340 2400 30665 2428
rect 30340 2388 30346 2400
rect 30653 2397 30665 2400
rect 30699 2397 30711 2431
rect 30653 2391 30711 2397
rect 31570 2388 31576 2440
rect 31628 2428 31634 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 31628 2400 32321 2428
rect 31628 2388 31634 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 33042 2388 33048 2440
rect 33100 2428 33106 2440
rect 33597 2431 33655 2437
rect 33597 2428 33609 2431
rect 33100 2400 33609 2428
rect 33100 2388 33106 2400
rect 33597 2397 33609 2400
rect 33643 2397 33655 2431
rect 33597 2391 33655 2397
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34848 2400 34897 2428
rect 34848 2388 34854 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 35866 2428 35894 2536
rect 36173 2431 36231 2437
rect 36173 2428 36185 2431
rect 35866 2400 36185 2428
rect 34885 2391 34943 2397
rect 36173 2397 36185 2400
rect 36219 2397 36231 2431
rect 38010 2428 38016 2440
rect 37971 2400 38016 2428
rect 36173 2391 36231 2397
rect 38010 2388 38016 2400
rect 38068 2388 38074 2440
rect 27120 2332 28028 2360
rect 27120 2320 27126 2332
rect 28350 2320 28356 2372
rect 28408 2360 28414 2372
rect 28537 2363 28595 2369
rect 28537 2360 28549 2363
rect 28408 2332 28549 2360
rect 28408 2320 28414 2332
rect 28537 2329 28549 2332
rect 28583 2329 28595 2363
rect 28537 2323 28595 2329
rect 22186 2292 22192 2304
rect 19260 2264 22192 2292
rect 17681 2255 17739 2261
rect 22186 2252 22192 2264
rect 22244 2252 22250 2304
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 22833 2295 22891 2301
rect 22833 2292 22845 2295
rect 22612 2264 22845 2292
rect 22612 2252 22618 2264
rect 22833 2261 22845 2264
rect 22879 2261 22891 2295
rect 24670 2292 24676 2304
rect 24631 2264 24676 2292
rect 22833 2255 22891 2261
rect 24670 2252 24676 2264
rect 24728 2252 24734 2304
rect 25130 2252 25136 2304
rect 25188 2292 25194 2304
rect 25409 2295 25467 2301
rect 25409 2292 25421 2295
rect 25188 2264 25421 2292
rect 25188 2252 25194 2264
rect 25409 2261 25421 2264
rect 25455 2261 25467 2295
rect 25409 2255 25467 2261
rect 25774 2252 25780 2304
rect 25832 2292 25838 2304
rect 26145 2295 26203 2301
rect 26145 2292 26157 2295
rect 25832 2264 26157 2292
rect 25832 2252 25838 2264
rect 26145 2261 26157 2264
rect 26191 2261 26203 2295
rect 27154 2292 27160 2304
rect 27115 2264 27160 2292
rect 26145 2255 26203 2261
rect 27154 2252 27160 2264
rect 27212 2252 27218 2304
rect 29638 2252 29644 2304
rect 29696 2292 29702 2304
rect 29917 2295 29975 2301
rect 29917 2292 29929 2295
rect 29696 2264 29929 2292
rect 29696 2252 29702 2264
rect 29917 2261 29929 2264
rect 29963 2261 29975 2295
rect 29917 2255 29975 2261
rect 32858 2252 32864 2304
rect 32916 2292 32922 2304
rect 33781 2295 33839 2301
rect 33781 2292 33793 2295
rect 32916 2264 33793 2292
rect 32916 2252 32922 2264
rect 33781 2261 33793 2264
rect 33827 2261 33839 2295
rect 33781 2255 33839 2261
rect 34790 2252 34796 2304
rect 34848 2292 34854 2304
rect 35069 2295 35127 2301
rect 35069 2292 35081 2295
rect 34848 2264 35081 2292
rect 34848 2252 34854 2264
rect 35069 2261 35081 2264
rect 35115 2261 35127 2295
rect 35069 2255 35127 2261
rect 36078 2252 36084 2304
rect 36136 2292 36142 2304
rect 36357 2295 36415 2301
rect 36357 2292 36369 2295
rect 36136 2264 36369 2292
rect 36136 2252 36142 2264
rect 36357 2261 36369 2264
rect 36403 2261 36415 2295
rect 36357 2255 36415 2261
rect 38197 2295 38255 2301
rect 38197 2261 38209 2295
rect 38243 2292 38255 2295
rect 39298 2292 39304 2304
rect 38243 2264 39304 2292
rect 38243 2261 38255 2264
rect 38197 2255 38255 2261
rect 39298 2252 39304 2264
rect 39356 2252 39362 2304
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 3970 2048 3976 2100
rect 4028 2088 4034 2100
rect 11974 2088 11980 2100
rect 4028 2060 11980 2088
rect 4028 2048 4034 2060
rect 11974 2048 11980 2060
rect 12032 2048 12038 2100
rect 18230 2048 18236 2100
rect 18288 2088 18294 2100
rect 22370 2088 22376 2100
rect 18288 2060 22376 2088
rect 18288 2048 18294 2060
rect 22370 2048 22376 2060
rect 22428 2048 22434 2100
rect 7834 1980 7840 2032
rect 7892 2020 7898 2032
rect 15562 2020 15568 2032
rect 7892 1992 15568 2020
rect 7892 1980 7898 1992
rect 15562 1980 15568 1992
rect 15620 1980 15626 2032
rect 16758 1980 16764 2032
rect 16816 2020 16822 2032
rect 25314 2020 25320 2032
rect 16816 1992 25320 2020
rect 16816 1980 16822 1992
rect 25314 1980 25320 1992
rect 25372 1980 25378 2032
rect 4982 1912 4988 1964
rect 5040 1952 5046 1964
rect 14458 1952 14464 1964
rect 5040 1924 14464 1952
rect 5040 1912 5046 1924
rect 14458 1912 14464 1924
rect 14516 1912 14522 1964
rect 15930 1912 15936 1964
rect 15988 1952 15994 1964
rect 19150 1952 19156 1964
rect 15988 1924 19156 1952
rect 15988 1912 15994 1924
rect 19150 1912 19156 1924
rect 19208 1912 19214 1964
rect 8478 1844 8484 1896
rect 8536 1884 8542 1896
rect 12526 1884 12532 1896
rect 8536 1856 12532 1884
rect 8536 1844 8542 1856
rect 12526 1844 12532 1856
rect 12584 1844 12590 1896
rect 24670 1884 24676 1896
rect 13464 1856 24676 1884
rect 10594 1776 10600 1828
rect 10652 1816 10658 1828
rect 13464 1816 13492 1856
rect 24670 1844 24676 1856
rect 24728 1844 24734 1896
rect 20070 1816 20076 1828
rect 10652 1788 13492 1816
rect 15764 1788 20076 1816
rect 10652 1776 10658 1788
rect 14458 1708 14464 1760
rect 14516 1748 14522 1760
rect 15764 1748 15792 1788
rect 20070 1776 20076 1788
rect 20128 1776 20134 1828
rect 14516 1720 15792 1748
rect 14516 1708 14522 1720
rect 18046 1708 18052 1760
rect 18104 1748 18110 1760
rect 27338 1748 27344 1760
rect 18104 1720 27344 1748
rect 18104 1708 18110 1720
rect 27338 1708 27344 1720
rect 27396 1708 27402 1760
rect 12526 1640 12532 1692
rect 12584 1680 12590 1692
rect 15654 1680 15660 1692
rect 12584 1652 15660 1680
rect 12584 1640 12590 1652
rect 15654 1640 15660 1652
rect 15712 1640 15718 1692
rect 16942 1640 16948 1692
rect 17000 1680 17006 1692
rect 22646 1680 22652 1692
rect 17000 1652 22652 1680
rect 17000 1640 17006 1652
rect 22646 1640 22652 1652
rect 22704 1640 22710 1692
rect 23842 1640 23848 1692
rect 23900 1680 23906 1692
rect 25406 1680 25412 1692
rect 23900 1652 25412 1680
rect 23900 1640 23906 1652
rect 25406 1640 25412 1652
rect 25464 1640 25470 1692
rect 13538 1572 13544 1624
rect 13596 1612 13602 1624
rect 22922 1612 22928 1624
rect 13596 1584 22928 1612
rect 13596 1572 13602 1584
rect 22922 1572 22928 1584
rect 22980 1572 22986 1624
rect 7282 1504 7288 1556
rect 7340 1544 7346 1556
rect 20438 1544 20444 1556
rect 7340 1516 20444 1544
rect 7340 1504 7346 1516
rect 20438 1504 20444 1516
rect 20496 1504 20502 1556
rect 4706 1436 4712 1488
rect 4764 1476 4770 1488
rect 18782 1476 18788 1488
rect 4764 1448 18788 1476
rect 4764 1436 4770 1448
rect 18782 1436 18788 1448
rect 18840 1436 18846 1488
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 1768 37451 1820 37460
rect 1768 37417 1777 37451
rect 1777 37417 1811 37451
rect 1811 37417 1820 37451
rect 1768 37408 1820 37417
rect 18512 37272 18564 37324
rect 21272 37272 21324 37324
rect 32772 37272 32824 37324
rect 2412 37204 2464 37256
rect 2780 37204 2832 37256
rect 3976 37247 4028 37256
rect 3976 37213 3985 37247
rect 3985 37213 4019 37247
rect 4019 37213 4028 37247
rect 3976 37204 4028 37213
rect 4620 37204 4672 37256
rect 5816 37204 5868 37256
rect 6460 37204 6512 37256
rect 7840 37247 7892 37256
rect 7840 37213 7849 37247
rect 7849 37213 7883 37247
rect 7883 37213 7892 37247
rect 7840 37204 7892 37213
rect 9772 37247 9824 37256
rect 9772 37213 9781 37247
rect 9781 37213 9815 37247
rect 9815 37213 9824 37247
rect 9772 37204 9824 37213
rect 6828 37136 6880 37188
rect 9496 37136 9548 37188
rect 12440 37204 12492 37256
rect 14188 37204 14240 37256
rect 14280 37247 14332 37256
rect 14280 37213 14289 37247
rect 14289 37213 14323 37247
rect 14323 37213 14332 37247
rect 14280 37204 14332 37213
rect 14832 37204 14884 37256
rect 18696 37247 18748 37256
rect 18696 37213 18705 37247
rect 18705 37213 18739 37247
rect 18739 37213 18748 37247
rect 18696 37204 18748 37213
rect 20076 37247 20128 37256
rect 20076 37213 20085 37247
rect 20085 37213 20119 37247
rect 20119 37213 20128 37247
rect 20076 37204 20128 37213
rect 21456 37204 21508 37256
rect 19064 37136 19116 37188
rect 21824 37136 21876 37188
rect 25136 37204 25188 37256
rect 26424 37204 26476 37256
rect 27896 37247 27948 37256
rect 27896 37213 27905 37247
rect 27905 37213 27939 37247
rect 27939 37213 27948 37247
rect 27896 37204 27948 37213
rect 28356 37204 28408 37256
rect 29644 37204 29696 37256
rect 30932 37204 30984 37256
rect 32312 37247 32364 37256
rect 32312 37213 32321 37247
rect 32321 37213 32355 37247
rect 32355 37213 32364 37247
rect 32312 37204 32364 37213
rect 32404 37204 32456 37256
rect 34796 37204 34848 37256
rect 36084 37204 36136 37256
rect 37372 37204 37424 37256
rect 28264 37136 28316 37188
rect 3240 37068 3292 37120
rect 4712 37111 4764 37120
rect 4712 37077 4721 37111
rect 4721 37077 4755 37111
rect 4755 37077 4764 37111
rect 4712 37068 4764 37077
rect 6368 37068 6420 37120
rect 6552 37111 6604 37120
rect 6552 37077 6561 37111
rect 6561 37077 6595 37111
rect 6595 37077 6604 37111
rect 6552 37068 6604 37077
rect 7748 37068 7800 37120
rect 9680 37068 9732 37120
rect 11060 37068 11112 37120
rect 12440 37111 12492 37120
rect 12440 37077 12449 37111
rect 12449 37077 12483 37111
rect 12483 37077 12492 37111
rect 12440 37068 12492 37077
rect 12900 37068 12952 37120
rect 13820 37068 13872 37120
rect 15476 37068 15528 37120
rect 17408 37068 17460 37120
rect 19984 37068 20036 37120
rect 24492 37068 24544 37120
rect 25320 37111 25372 37120
rect 25320 37077 25329 37111
rect 25329 37077 25363 37111
rect 25363 37077 25372 37111
rect 25320 37068 25372 37077
rect 27712 37068 27764 37120
rect 28632 37111 28684 37120
rect 28632 37077 28641 37111
rect 28641 37077 28675 37111
rect 28675 37077 28684 37111
rect 28632 37068 28684 37077
rect 28724 37068 28776 37120
rect 32220 37068 32272 37120
rect 33140 37068 33192 37120
rect 34520 37068 34572 37120
rect 36360 37111 36412 37120
rect 36360 37077 36369 37111
rect 36369 37077 36403 37111
rect 36403 37077 36412 37111
rect 36360 37068 36412 37077
rect 37648 37111 37700 37120
rect 37648 37077 37657 37111
rect 37657 37077 37691 37111
rect 37691 37077 37700 37111
rect 37648 37068 37700 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 1676 36864 1728 36916
rect 9036 36864 9088 36916
rect 14832 36907 14884 36916
rect 14832 36873 14841 36907
rect 14841 36873 14875 36907
rect 14875 36873 14884 36907
rect 14832 36864 14884 36873
rect 16764 36864 16816 36916
rect 20 36796 72 36848
rect 2504 36771 2556 36780
rect 2504 36737 2513 36771
rect 2513 36737 2547 36771
rect 2547 36737 2556 36771
rect 2504 36728 2556 36737
rect 7840 36796 7892 36848
rect 22836 36864 22888 36916
rect 32312 36864 32364 36916
rect 19340 36796 19392 36848
rect 38108 36839 38160 36848
rect 9128 36771 9180 36780
rect 9128 36737 9137 36771
rect 9137 36737 9171 36771
rect 9171 36737 9180 36771
rect 9128 36728 9180 36737
rect 14096 36771 14148 36780
rect 14096 36737 14105 36771
rect 14105 36737 14139 36771
rect 14139 36737 14148 36771
rect 14096 36728 14148 36737
rect 16856 36771 16908 36780
rect 16856 36737 16865 36771
rect 16865 36737 16899 36771
rect 16899 36737 16908 36771
rect 16856 36728 16908 36737
rect 22100 36728 22152 36780
rect 23204 36728 23256 36780
rect 4068 36660 4120 36712
rect 35440 36728 35492 36780
rect 38108 36805 38117 36839
rect 38117 36805 38151 36839
rect 38151 36805 38160 36839
rect 38108 36796 38160 36805
rect 39304 36728 39356 36780
rect 37648 36660 37700 36712
rect 14280 36592 14332 36644
rect 22100 36592 22152 36644
rect 33140 36592 33192 36644
rect 38384 36592 38436 36644
rect 2320 36567 2372 36576
rect 2320 36533 2329 36567
rect 2329 36533 2363 36567
rect 2363 36533 2372 36567
rect 2320 36524 2372 36533
rect 5816 36524 5868 36576
rect 20720 36524 20772 36576
rect 35532 36567 35584 36576
rect 35532 36533 35541 36567
rect 35541 36533 35575 36567
rect 35575 36533 35584 36567
rect 35532 36524 35584 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 20076 36320 20128 36372
rect 37188 36320 37240 36372
rect 27620 36184 27672 36236
rect 28724 36184 28776 36236
rect 1308 36116 1360 36168
rect 19984 36116 20036 36168
rect 38476 36184 38528 36236
rect 33232 36048 33284 36100
rect 2596 35980 2648 36032
rect 38200 36023 38252 36032
rect 38200 35989 38209 36023
rect 38209 35989 38243 36023
rect 38243 35989 38252 36023
rect 38200 35980 38252 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 38108 35683 38160 35692
rect 38108 35649 38117 35683
rect 38117 35649 38151 35683
rect 38151 35649 38160 35683
rect 38108 35640 38160 35649
rect 1584 35615 1636 35624
rect 1584 35581 1593 35615
rect 1593 35581 1627 35615
rect 1627 35581 1636 35615
rect 1584 35572 1636 35581
rect 7472 35572 7524 35624
rect 37648 35436 37700 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 3976 35232 4028 35284
rect 19984 35232 20036 35284
rect 1768 35071 1820 35080
rect 1768 35037 1777 35071
rect 1777 35037 1811 35071
rect 1811 35037 1820 35071
rect 1768 35028 1820 35037
rect 1860 35028 1912 35080
rect 19432 35071 19484 35080
rect 19432 35037 19441 35071
rect 19441 35037 19475 35071
rect 19475 35037 19484 35071
rect 19432 35028 19484 35037
rect 38660 35028 38712 35080
rect 2688 34892 2740 34944
rect 37280 34892 37332 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4068 34688 4120 34740
rect 5724 34552 5776 34604
rect 38568 34552 38620 34604
rect 38200 34391 38252 34400
rect 38200 34357 38209 34391
rect 38209 34357 38243 34391
rect 38243 34357 38252 34391
rect 38200 34348 38252 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 21824 34144 21876 34196
rect 21364 33940 21416 33992
rect 2412 33804 2464 33856
rect 17408 33804 17460 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4068 33464 4120 33516
rect 4712 33464 4764 33516
rect 1768 33371 1820 33380
rect 1768 33337 1777 33371
rect 1777 33337 1811 33371
rect 1811 33337 1820 33371
rect 1768 33328 1820 33337
rect 9312 33260 9364 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 33232 33099 33284 33108
rect 33232 33065 33241 33099
rect 33241 33065 33275 33099
rect 33275 33065 33284 33099
rect 33232 33056 33284 33065
rect 6552 32852 6604 32904
rect 13636 32852 13688 32904
rect 28264 32895 28316 32904
rect 28264 32861 28273 32895
rect 28273 32861 28307 32895
rect 28307 32861 28316 32895
rect 28264 32852 28316 32861
rect 30472 32852 30524 32904
rect 38108 32827 38160 32836
rect 38108 32793 38117 32827
rect 38117 32793 38151 32827
rect 38151 32793 38160 32827
rect 38108 32784 38160 32793
rect 10140 32716 10192 32768
rect 10784 32716 10836 32768
rect 28356 32759 28408 32768
rect 28356 32725 28365 32759
rect 28365 32725 28399 32759
rect 28399 32725 28408 32759
rect 28356 32716 28408 32725
rect 38200 32759 38252 32768
rect 38200 32725 38209 32759
rect 38209 32725 38243 32759
rect 38243 32725 38252 32759
rect 38200 32716 38252 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 9496 32512 9548 32564
rect 9772 32512 9824 32564
rect 9220 32419 9272 32428
rect 9220 32385 9229 32419
rect 9229 32385 9263 32419
rect 9263 32385 9272 32419
rect 9220 32376 9272 32385
rect 10784 32419 10836 32428
rect 10784 32385 10793 32419
rect 10793 32385 10827 32419
rect 10827 32385 10836 32419
rect 10784 32376 10836 32385
rect 20720 32419 20772 32428
rect 20720 32385 20729 32419
rect 20729 32385 20763 32419
rect 20763 32385 20772 32419
rect 20720 32376 20772 32385
rect 28632 32376 28684 32428
rect 38108 32419 38160 32428
rect 38108 32385 38117 32419
rect 38117 32385 38151 32419
rect 38151 32385 38160 32419
rect 38108 32376 38160 32385
rect 1768 32215 1820 32224
rect 1768 32181 1777 32215
rect 1777 32181 1811 32215
rect 1811 32181 1820 32215
rect 1768 32172 1820 32181
rect 2228 32215 2280 32224
rect 2228 32181 2237 32215
rect 2237 32181 2271 32215
rect 2271 32181 2280 32215
rect 2228 32172 2280 32181
rect 20628 32172 20680 32224
rect 23572 32215 23624 32224
rect 23572 32181 23581 32215
rect 23581 32181 23615 32215
rect 23615 32181 23624 32215
rect 23572 32172 23624 32181
rect 37924 32172 37976 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 2228 31968 2280 32020
rect 17224 31968 17276 32020
rect 18788 31968 18840 32020
rect 15384 31900 15436 31952
rect 23572 31900 23624 31952
rect 1860 31875 1912 31884
rect 1860 31841 1869 31875
rect 1869 31841 1903 31875
rect 1903 31841 1912 31875
rect 1860 31832 1912 31841
rect 2964 31832 3016 31884
rect 20720 31832 20772 31884
rect 1584 31807 1636 31816
rect 1584 31773 1593 31807
rect 1593 31773 1627 31807
rect 1627 31773 1636 31807
rect 1584 31764 1636 31773
rect 25320 31832 25372 31884
rect 27804 31832 27856 31884
rect 27620 31764 27672 31816
rect 35532 31764 35584 31816
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 33140 31288 33192 31340
rect 17592 31084 17644 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 9220 30880 9272 30932
rect 27896 30880 27948 30932
rect 9772 30812 9824 30864
rect 2596 30744 2648 30796
rect 2320 30676 2372 30728
rect 5816 30719 5868 30728
rect 5816 30685 5825 30719
rect 5825 30685 5859 30719
rect 5859 30685 5868 30719
rect 5816 30676 5868 30685
rect 6368 30676 6420 30728
rect 7656 30676 7708 30728
rect 12440 30676 12492 30728
rect 12900 30719 12952 30728
rect 12900 30685 12909 30719
rect 12909 30685 12943 30719
rect 12943 30685 12952 30719
rect 12900 30676 12952 30685
rect 26148 30719 26200 30728
rect 26148 30685 26157 30719
rect 26157 30685 26191 30719
rect 26191 30685 26200 30719
rect 26148 30676 26200 30685
rect 37280 30812 37332 30864
rect 9864 30608 9916 30660
rect 37464 30719 37516 30728
rect 37464 30685 37473 30719
rect 37473 30685 37507 30719
rect 37507 30685 37516 30719
rect 37464 30676 37516 30685
rect 5356 30540 5408 30592
rect 6552 30583 6604 30592
rect 6552 30549 6561 30583
rect 6561 30549 6595 30583
rect 6595 30549 6604 30583
rect 6552 30540 6604 30549
rect 10324 30540 10376 30592
rect 13360 30540 13412 30592
rect 28080 30583 28132 30592
rect 28080 30549 28089 30583
rect 28089 30549 28123 30583
rect 28123 30549 28132 30583
rect 28080 30540 28132 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 13268 30336 13320 30388
rect 14096 30336 14148 30388
rect 2688 30200 2740 30252
rect 5172 30132 5224 30184
rect 1768 30039 1820 30048
rect 1768 30005 1777 30039
rect 1777 30005 1811 30039
rect 1811 30005 1820 30039
rect 1768 29996 1820 30005
rect 4988 29996 5040 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 4068 29792 4120 29844
rect 30472 29792 30524 29844
rect 16764 29656 16816 29708
rect 32404 29656 32456 29708
rect 1768 29631 1820 29640
rect 1768 29597 1777 29631
rect 1777 29597 1811 29631
rect 1811 29597 1820 29631
rect 1768 29588 1820 29597
rect 5816 29588 5868 29640
rect 6828 29588 6880 29640
rect 16212 29588 16264 29640
rect 17960 29588 18012 29640
rect 37372 29588 37424 29640
rect 14280 29520 14332 29572
rect 4712 29452 4764 29504
rect 11888 29452 11940 29504
rect 17684 29495 17736 29504
rect 17684 29461 17693 29495
rect 17693 29461 17727 29495
rect 17727 29461 17736 29495
rect 17684 29452 17736 29461
rect 38200 29495 38252 29504
rect 38200 29461 38209 29495
rect 38209 29461 38243 29495
rect 38243 29461 38252 29495
rect 38200 29452 38252 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 5724 29248 5776 29300
rect 16856 29291 16908 29300
rect 16856 29257 16865 29291
rect 16865 29257 16899 29291
rect 16899 29257 16908 29291
rect 16856 29248 16908 29257
rect 2780 29112 2832 29164
rect 8300 29112 8352 29164
rect 11888 29155 11940 29164
rect 11888 29121 11897 29155
rect 11897 29121 11931 29155
rect 11931 29121 11940 29155
rect 11888 29112 11940 29121
rect 16672 29112 16724 29164
rect 17684 29155 17736 29164
rect 17684 29121 17693 29155
rect 17693 29121 17727 29155
rect 17727 29121 17736 29155
rect 17684 29112 17736 29121
rect 1584 29019 1636 29028
rect 1584 28985 1593 29019
rect 1593 28985 1627 29019
rect 1627 28985 1636 29019
rect 1584 28976 1636 28985
rect 10600 28976 10652 29028
rect 17500 28951 17552 28960
rect 17500 28917 17509 28951
rect 17509 28917 17543 28951
rect 17543 28917 17552 28951
rect 17500 28908 17552 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 16856 28636 16908 28688
rect 756 28568 808 28620
rect 1860 28543 1912 28552
rect 1860 28509 1869 28543
rect 1869 28509 1903 28543
rect 1903 28509 1912 28543
rect 1860 28500 1912 28509
rect 17500 28568 17552 28620
rect 15752 28500 15804 28552
rect 16212 28543 16264 28552
rect 16212 28509 16221 28543
rect 16221 28509 16255 28543
rect 16255 28509 16264 28543
rect 16212 28500 16264 28509
rect 16948 28500 17000 28552
rect 2872 28432 2924 28484
rect 2320 28364 2372 28416
rect 17500 28364 17552 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 5816 28203 5868 28212
rect 5816 28169 5825 28203
rect 5825 28169 5859 28203
rect 5859 28169 5868 28203
rect 5816 28160 5868 28169
rect 16948 28203 17000 28212
rect 16948 28169 16957 28203
rect 16957 28169 16991 28203
rect 16991 28169 17000 28203
rect 16948 28160 17000 28169
rect 21364 28203 21416 28212
rect 21364 28169 21373 28203
rect 21373 28169 21407 28203
rect 21407 28169 21416 28203
rect 21364 28160 21416 28169
rect 1952 28067 2004 28076
rect 1952 28033 1961 28067
rect 1961 28033 1995 28067
rect 1995 28033 2004 28067
rect 1952 28024 2004 28033
rect 2596 28067 2648 28076
rect 2596 28033 2605 28067
rect 2605 28033 2639 28067
rect 2639 28033 2648 28067
rect 2596 28024 2648 28033
rect 3424 28067 3476 28076
rect 3424 28033 3433 28067
rect 3433 28033 3467 28067
rect 3467 28033 3476 28067
rect 3424 28024 3476 28033
rect 4068 28067 4120 28076
rect 4068 28033 4077 28067
rect 4077 28033 4111 28067
rect 4111 28033 4120 28067
rect 4068 28024 4120 28033
rect 6460 28024 6512 28076
rect 8392 28024 8444 28076
rect 12624 28067 12676 28076
rect 12624 28033 12633 28067
rect 12633 28033 12667 28067
rect 12667 28033 12676 28067
rect 12624 28024 12676 28033
rect 17684 28067 17736 28076
rect 17684 28033 17693 28067
rect 17693 28033 17727 28067
rect 17727 28033 17736 28067
rect 17684 28024 17736 28033
rect 19248 28067 19300 28076
rect 19248 28033 19257 28067
rect 19257 28033 19291 28067
rect 19291 28033 19300 28067
rect 19248 28024 19300 28033
rect 1584 27888 1636 27940
rect 9680 27956 9732 28008
rect 16948 27956 17000 28008
rect 37464 27999 37516 28008
rect 37464 27965 37473 27999
rect 37473 27965 37507 27999
rect 37507 27965 37516 27999
rect 37464 27956 37516 27965
rect 37832 27956 37884 28008
rect 2044 27863 2096 27872
rect 2044 27829 2053 27863
rect 2053 27829 2087 27863
rect 2087 27829 2096 27863
rect 2044 27820 2096 27829
rect 3240 27863 3292 27872
rect 3240 27829 3249 27863
rect 3249 27829 3283 27863
rect 3283 27829 3292 27863
rect 3240 27820 3292 27829
rect 5080 27820 5132 27872
rect 8208 27820 8260 27872
rect 11152 27820 11204 27872
rect 17040 27820 17092 27872
rect 17868 27820 17920 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 17684 27616 17736 27668
rect 12072 27548 12124 27600
rect 6552 27480 6604 27532
rect 10600 27523 10652 27532
rect 10600 27489 10609 27523
rect 10609 27489 10643 27523
rect 10643 27489 10652 27523
rect 10600 27480 10652 27489
rect 15752 27480 15804 27532
rect 1860 27455 1912 27464
rect 1860 27421 1869 27455
rect 1869 27421 1903 27455
rect 1903 27421 1912 27455
rect 1860 27412 1912 27421
rect 2504 27455 2556 27464
rect 2504 27421 2513 27455
rect 2513 27421 2547 27455
rect 2547 27421 2556 27455
rect 2504 27412 2556 27421
rect 3240 27412 3292 27464
rect 8392 27412 8444 27464
rect 8944 27412 8996 27464
rect 3884 27344 3936 27396
rect 13176 27412 13228 27464
rect 17500 27480 17552 27532
rect 19248 27616 19300 27668
rect 37372 27591 37424 27600
rect 37372 27557 37381 27591
rect 37381 27557 37415 27591
rect 37415 27557 37424 27591
rect 37372 27548 37424 27557
rect 19340 27412 19392 27464
rect 22100 27455 22152 27464
rect 22100 27421 22109 27455
rect 22109 27421 22143 27455
rect 22143 27421 22152 27455
rect 37556 27455 37608 27464
rect 22100 27412 22152 27421
rect 37556 27421 37565 27455
rect 37565 27421 37599 27455
rect 37599 27421 37608 27455
rect 37556 27412 37608 27421
rect 38016 27455 38068 27464
rect 38016 27421 38025 27455
rect 38025 27421 38059 27455
rect 38059 27421 38068 27455
rect 38016 27412 38068 27421
rect 20352 27344 20404 27396
rect 1952 27319 2004 27328
rect 1952 27285 1961 27319
rect 1961 27285 1995 27319
rect 1995 27285 2004 27319
rect 1952 27276 2004 27285
rect 2136 27276 2188 27328
rect 3700 27276 3752 27328
rect 7840 27319 7892 27328
rect 7840 27285 7849 27319
rect 7849 27285 7883 27319
rect 7883 27285 7892 27319
rect 7840 27276 7892 27285
rect 10048 27276 10100 27328
rect 11980 27276 12032 27328
rect 12624 27276 12676 27328
rect 12716 27276 12768 27328
rect 18144 27319 18196 27328
rect 18144 27285 18153 27319
rect 18153 27285 18187 27319
rect 18187 27285 18196 27319
rect 18144 27276 18196 27285
rect 18788 27276 18840 27328
rect 22560 27276 22612 27328
rect 38200 27319 38252 27328
rect 38200 27285 38209 27319
rect 38209 27285 38243 27319
rect 38243 27285 38252 27319
rect 38200 27276 38252 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 2964 27072 3016 27124
rect 5172 27115 5224 27124
rect 1216 27004 1268 27056
rect 5172 27081 5181 27115
rect 5181 27081 5215 27115
rect 5215 27081 5224 27115
rect 5172 27072 5224 27081
rect 11152 27072 11204 27124
rect 12716 27047 12768 27056
rect 572 26936 624 26988
rect 1860 26979 1912 26988
rect 1860 26945 1869 26979
rect 1869 26945 1903 26979
rect 1903 26945 1912 26979
rect 1860 26936 1912 26945
rect 2964 26936 3016 26988
rect 3056 26868 3108 26920
rect 6828 26936 6880 26988
rect 12716 27013 12725 27047
rect 12725 27013 12759 27047
rect 12759 27013 12768 27047
rect 12716 27004 12768 27013
rect 11244 26936 11296 26988
rect 5264 26868 5316 26920
rect 848 26800 900 26852
rect 1124 26732 1176 26784
rect 3148 26732 3200 26784
rect 4620 26732 4672 26784
rect 7288 26732 7340 26784
rect 12164 26732 12216 26784
rect 12716 26868 12768 26920
rect 17500 27072 17552 27124
rect 28080 27072 28132 27124
rect 37556 27115 37608 27124
rect 37556 27081 37565 27115
rect 37565 27081 37599 27115
rect 37599 27081 37608 27115
rect 37556 27072 37608 27081
rect 17040 27047 17092 27056
rect 17040 27013 17049 27047
rect 17049 27013 17083 27047
rect 17083 27013 17092 27047
rect 17040 27004 17092 27013
rect 17960 27004 18012 27056
rect 22100 26936 22152 26988
rect 37280 26936 37332 26988
rect 18144 26868 18196 26920
rect 22468 26868 22520 26920
rect 28356 26868 28408 26920
rect 16856 26732 16908 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 8300 26571 8352 26580
rect 8300 26537 8309 26571
rect 8309 26537 8343 26571
rect 8343 26537 8352 26571
rect 8300 26528 8352 26537
rect 11244 26528 11296 26580
rect 12992 26528 13044 26580
rect 13176 26571 13228 26580
rect 13176 26537 13185 26571
rect 13185 26537 13219 26571
rect 13219 26537 13228 26571
rect 13176 26528 13228 26537
rect 14832 26528 14884 26580
rect 15844 26528 15896 26580
rect 664 26392 716 26444
rect 9588 26460 9640 26512
rect 12256 26460 12308 26512
rect 7840 26435 7892 26444
rect 1860 26367 1912 26376
rect 1860 26333 1869 26367
rect 1869 26333 1903 26367
rect 1903 26333 1912 26367
rect 1860 26324 1912 26333
rect 2504 26367 2556 26376
rect 2504 26333 2513 26367
rect 2513 26333 2547 26367
rect 2547 26333 2556 26367
rect 2504 26324 2556 26333
rect 2964 26324 3016 26376
rect 7840 26401 7849 26435
rect 7849 26401 7883 26435
rect 7883 26401 7892 26435
rect 7840 26392 7892 26401
rect 12072 26435 12124 26444
rect 12072 26401 12081 26435
rect 12081 26401 12115 26435
rect 12115 26401 12124 26435
rect 12072 26392 12124 26401
rect 12440 26435 12492 26444
rect 12440 26401 12449 26435
rect 12449 26401 12483 26435
rect 12483 26401 12492 26435
rect 20628 26435 20680 26444
rect 12440 26392 12492 26401
rect 5172 26367 5224 26376
rect 5172 26333 5181 26367
rect 5181 26333 5215 26367
rect 5215 26333 5224 26367
rect 5172 26324 5224 26333
rect 5448 26324 5500 26376
rect 6092 26324 6144 26376
rect 6920 26367 6972 26376
rect 6920 26333 6929 26367
rect 6929 26333 6963 26367
rect 6963 26333 6972 26367
rect 6920 26324 6972 26333
rect 11060 26324 11112 26376
rect 12992 26324 13044 26376
rect 14372 26367 14424 26376
rect 14372 26333 14381 26367
rect 14381 26333 14415 26367
rect 14415 26333 14424 26367
rect 14372 26324 14424 26333
rect 16120 26367 16172 26376
rect 16120 26333 16129 26367
rect 16129 26333 16163 26367
rect 16163 26333 16172 26367
rect 16120 26324 16172 26333
rect 20628 26401 20637 26435
rect 20637 26401 20671 26435
rect 20671 26401 20680 26435
rect 20628 26392 20680 26401
rect 34520 26460 34572 26512
rect 38292 26367 38344 26376
rect 38292 26333 38301 26367
rect 38301 26333 38335 26367
rect 38335 26333 38344 26367
rect 38292 26324 38344 26333
rect 1952 26299 2004 26308
rect 1952 26265 1961 26299
rect 1961 26265 1995 26299
rect 1995 26265 2004 26299
rect 1952 26256 2004 26265
rect 2688 26256 2740 26308
rect 11428 26256 11480 26308
rect 12164 26299 12216 26308
rect 12164 26265 12173 26299
rect 12173 26265 12207 26299
rect 12207 26265 12216 26299
rect 12164 26256 12216 26265
rect 20812 26256 20864 26308
rect 16580 26231 16632 26240
rect 16580 26197 16589 26231
rect 16589 26197 16623 26231
rect 16623 26197 16632 26231
rect 16580 26188 16632 26197
rect 17776 26231 17828 26240
rect 17776 26197 17785 26231
rect 17785 26197 17819 26231
rect 17819 26197 17828 26231
rect 17776 26188 17828 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 6828 25984 6880 26036
rect 2044 25916 2096 25968
rect 2688 25916 2740 25968
rect 1400 25848 1452 25900
rect 6000 25916 6052 25968
rect 17776 25959 17828 25968
rect 3976 25848 4028 25900
rect 4804 25891 4856 25900
rect 4804 25857 4813 25891
rect 4813 25857 4847 25891
rect 4847 25857 4856 25891
rect 4804 25848 4856 25857
rect 5632 25891 5684 25900
rect 5632 25857 5641 25891
rect 5641 25857 5675 25891
rect 5675 25857 5684 25891
rect 5632 25848 5684 25857
rect 6920 25848 6972 25900
rect 7748 25891 7800 25900
rect 5724 25780 5776 25832
rect 7748 25857 7757 25891
rect 7757 25857 7791 25891
rect 7791 25857 7800 25891
rect 7748 25848 7800 25857
rect 10692 25848 10744 25900
rect 14188 25848 14240 25900
rect 15016 25848 15068 25900
rect 17776 25925 17785 25959
rect 17785 25925 17819 25959
rect 17819 25925 17828 25959
rect 17776 25916 17828 25925
rect 17868 25959 17920 25968
rect 17868 25925 17877 25959
rect 17877 25925 17911 25959
rect 17911 25925 17920 25959
rect 17868 25916 17920 25925
rect 7840 25780 7892 25832
rect 9680 25823 9732 25832
rect 9680 25789 9689 25823
rect 9689 25789 9723 25823
rect 9723 25789 9732 25823
rect 9680 25780 9732 25789
rect 7012 25712 7064 25764
rect 16304 25780 16356 25832
rect 17960 25780 18012 25832
rect 2596 25644 2648 25696
rect 3332 25687 3384 25696
rect 3332 25653 3341 25687
rect 3341 25653 3375 25687
rect 3375 25653 3384 25687
rect 3332 25644 3384 25653
rect 3792 25644 3844 25696
rect 6184 25644 6236 25696
rect 6276 25644 6328 25696
rect 14096 25687 14148 25696
rect 14096 25653 14105 25687
rect 14105 25653 14139 25687
rect 14139 25653 14148 25687
rect 14096 25644 14148 25653
rect 14740 25687 14792 25696
rect 14740 25653 14749 25687
rect 14749 25653 14783 25687
rect 14783 25653 14792 25687
rect 14740 25644 14792 25653
rect 15292 25687 15344 25696
rect 15292 25653 15301 25687
rect 15301 25653 15335 25687
rect 15335 25653 15344 25687
rect 15292 25644 15344 25653
rect 18880 25644 18932 25696
rect 27804 25644 27856 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 2228 25236 2280 25288
rect 3608 25236 3660 25288
rect 7196 25440 7248 25492
rect 10692 25483 10744 25492
rect 10692 25449 10701 25483
rect 10701 25449 10735 25483
rect 10735 25449 10744 25483
rect 10692 25440 10744 25449
rect 20812 25440 20864 25492
rect 38016 25440 38068 25492
rect 7932 25372 7984 25424
rect 11428 25372 11480 25424
rect 6184 25347 6236 25356
rect 6184 25313 6193 25347
rect 6193 25313 6227 25347
rect 6227 25313 6236 25347
rect 6184 25304 6236 25313
rect 13636 25347 13688 25356
rect 13636 25313 13645 25347
rect 13645 25313 13679 25347
rect 13679 25313 13688 25347
rect 13636 25304 13688 25313
rect 1308 25168 1360 25220
rect 5632 25236 5684 25288
rect 6276 25236 6328 25288
rect 6368 25236 6420 25288
rect 9128 25279 9180 25288
rect 9128 25245 9137 25279
rect 9137 25245 9171 25279
rect 9171 25245 9180 25279
rect 9128 25236 9180 25245
rect 10876 25279 10928 25288
rect 10876 25245 10885 25279
rect 10885 25245 10919 25279
rect 10919 25245 10928 25279
rect 10876 25236 10928 25245
rect 15476 25236 15528 25288
rect 16120 25304 16172 25356
rect 16304 25347 16356 25356
rect 16304 25313 16313 25347
rect 16313 25313 16347 25347
rect 16347 25313 16356 25347
rect 16304 25304 16356 25313
rect 16948 25347 17000 25356
rect 16948 25313 16957 25347
rect 16957 25313 16991 25347
rect 16991 25313 17000 25347
rect 16948 25304 17000 25313
rect 19248 25236 19300 25288
rect 26148 25236 26200 25288
rect 30104 25279 30156 25288
rect 30104 25245 30113 25279
rect 30113 25245 30147 25279
rect 30147 25245 30156 25279
rect 30104 25236 30156 25245
rect 7748 25168 7800 25220
rect 8024 25168 8076 25220
rect 15292 25168 15344 25220
rect 16580 25168 16632 25220
rect 1768 25143 1820 25152
rect 1768 25109 1777 25143
rect 1777 25109 1811 25143
rect 1811 25109 1820 25143
rect 1768 25100 1820 25109
rect 1860 25100 1912 25152
rect 2872 25100 2924 25152
rect 4896 25100 4948 25152
rect 6736 25100 6788 25152
rect 8116 25143 8168 25152
rect 8116 25109 8125 25143
rect 8125 25109 8159 25143
rect 8159 25109 8168 25143
rect 8116 25100 8168 25109
rect 14372 25100 14424 25152
rect 14464 25100 14516 25152
rect 15200 25100 15252 25152
rect 17960 25100 18012 25152
rect 20812 25100 20864 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 2044 24760 2096 24812
rect 3884 24760 3936 24812
rect 4804 24896 4856 24948
rect 2412 24692 2464 24744
rect 2964 24692 3016 24744
rect 5540 24760 5592 24812
rect 8116 24760 8168 24812
rect 8208 24803 8260 24812
rect 8208 24769 8217 24803
rect 8217 24769 8251 24803
rect 8251 24769 8260 24803
rect 8208 24760 8260 24769
rect 6828 24692 6880 24744
rect 7012 24735 7064 24744
rect 7012 24701 7021 24735
rect 7021 24701 7055 24735
rect 7055 24701 7064 24735
rect 7012 24692 7064 24701
rect 7932 24692 7984 24744
rect 10140 24896 10192 24948
rect 10784 24896 10836 24948
rect 10048 24803 10100 24812
rect 10048 24769 10057 24803
rect 10057 24769 10091 24803
rect 10091 24769 10100 24803
rect 10048 24760 10100 24769
rect 10876 24760 10928 24812
rect 15292 24896 15344 24948
rect 14740 24828 14792 24880
rect 15200 24871 15252 24880
rect 15200 24837 15209 24871
rect 15209 24837 15243 24871
rect 15243 24837 15252 24871
rect 15200 24828 15252 24837
rect 17960 24871 18012 24880
rect 17960 24837 17969 24871
rect 17969 24837 18003 24871
rect 18003 24837 18012 24871
rect 17960 24828 18012 24837
rect 16948 24760 17000 24812
rect 11520 24692 11572 24744
rect 13360 24735 13412 24744
rect 13360 24701 13369 24735
rect 13369 24701 13403 24735
rect 13403 24701 13412 24735
rect 13360 24692 13412 24701
rect 14832 24692 14884 24744
rect 14924 24692 14976 24744
rect 15292 24692 15344 24744
rect 16212 24692 16264 24744
rect 32680 24760 32732 24812
rect 17592 24692 17644 24744
rect 17868 24735 17920 24744
rect 17868 24701 17877 24735
rect 17877 24701 17911 24735
rect 17911 24701 17920 24735
rect 17868 24692 17920 24701
rect 18696 24735 18748 24744
rect 18696 24701 18705 24735
rect 18705 24701 18739 24735
rect 18739 24701 18748 24735
rect 18696 24692 18748 24701
rect 940 24556 992 24608
rect 3424 24599 3476 24608
rect 3424 24565 3433 24599
rect 3433 24565 3467 24599
rect 3467 24565 3476 24599
rect 3424 24556 3476 24565
rect 8208 24624 8260 24676
rect 8300 24624 8352 24676
rect 8852 24624 8904 24676
rect 10692 24624 10744 24676
rect 10876 24624 10928 24676
rect 12716 24624 12768 24676
rect 17960 24624 18012 24676
rect 9128 24599 9180 24608
rect 9128 24565 9137 24599
rect 9137 24565 9171 24599
rect 9171 24565 9180 24599
rect 9128 24556 9180 24565
rect 9496 24556 9548 24608
rect 11060 24556 11112 24608
rect 12072 24556 12124 24608
rect 15292 24556 15344 24608
rect 15476 24556 15528 24608
rect 38200 24599 38252 24608
rect 38200 24565 38209 24599
rect 38209 24565 38243 24599
rect 38243 24565 38252 24599
rect 38200 24556 38252 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 6460 24352 6512 24404
rect 8852 24352 8904 24404
rect 9036 24352 9088 24404
rect 3976 24284 4028 24336
rect 1032 24080 1084 24132
rect 3516 24148 3568 24200
rect 3976 24191 4028 24200
rect 3976 24157 3985 24191
rect 3985 24157 4019 24191
rect 4019 24157 4028 24191
rect 3976 24148 4028 24157
rect 4804 24148 4856 24200
rect 5632 24080 5684 24132
rect 1768 24055 1820 24064
rect 1768 24021 1777 24055
rect 1777 24021 1811 24055
rect 1811 24021 1820 24055
rect 1768 24012 1820 24021
rect 2504 24012 2556 24064
rect 2964 24012 3016 24064
rect 5816 24012 5868 24064
rect 6828 24284 6880 24336
rect 7380 24284 7432 24336
rect 7564 24284 7616 24336
rect 12716 24352 12768 24404
rect 19064 24352 19116 24404
rect 20352 24395 20404 24404
rect 20352 24361 20361 24395
rect 20361 24361 20395 24395
rect 20395 24361 20404 24395
rect 20352 24352 20404 24361
rect 7012 24259 7064 24268
rect 7012 24225 7021 24259
rect 7021 24225 7055 24259
rect 7055 24225 7064 24259
rect 7012 24216 7064 24225
rect 7472 24216 7524 24268
rect 8760 24216 8812 24268
rect 15660 24284 15712 24336
rect 16488 24284 16540 24336
rect 23296 24284 23348 24336
rect 13636 24216 13688 24268
rect 14372 24259 14424 24268
rect 14372 24225 14381 24259
rect 14381 24225 14415 24259
rect 14415 24225 14424 24259
rect 14372 24216 14424 24225
rect 14832 24259 14884 24268
rect 14832 24225 14841 24259
rect 14841 24225 14875 24259
rect 14875 24225 14884 24259
rect 14832 24216 14884 24225
rect 15292 24216 15344 24268
rect 30104 24216 30156 24268
rect 6828 24148 6880 24200
rect 7656 24191 7708 24200
rect 7656 24157 7665 24191
rect 7665 24157 7699 24191
rect 7699 24157 7708 24191
rect 8208 24191 8260 24200
rect 7656 24148 7708 24157
rect 8208 24157 8217 24191
rect 8217 24157 8251 24191
rect 8251 24157 8260 24191
rect 8208 24148 8260 24157
rect 8668 24148 8720 24200
rect 10416 24148 10468 24200
rect 12532 24148 12584 24200
rect 6644 24080 6696 24132
rect 7196 24080 7248 24132
rect 8392 24123 8444 24132
rect 8392 24089 8401 24123
rect 8401 24089 8435 24123
rect 8435 24089 8444 24123
rect 8392 24080 8444 24089
rect 9220 24080 9272 24132
rect 12624 24080 12676 24132
rect 12808 24123 12860 24132
rect 12808 24089 12817 24123
rect 12817 24089 12851 24123
rect 12851 24089 12860 24123
rect 12808 24080 12860 24089
rect 14096 24080 14148 24132
rect 14464 24123 14516 24132
rect 14464 24089 14473 24123
rect 14473 24089 14507 24123
rect 14507 24089 14516 24123
rect 18420 24148 18472 24200
rect 18512 24191 18564 24200
rect 18512 24157 18521 24191
rect 18521 24157 18555 24191
rect 18555 24157 18564 24191
rect 18512 24148 18564 24157
rect 16396 24123 16448 24132
rect 14464 24080 14516 24089
rect 7472 24012 7524 24064
rect 10232 24012 10284 24064
rect 11060 24012 11112 24064
rect 13912 24012 13964 24064
rect 16396 24089 16405 24123
rect 16405 24089 16439 24123
rect 16439 24089 16448 24123
rect 16396 24080 16448 24089
rect 17776 24080 17828 24132
rect 21456 24148 21508 24200
rect 34520 24148 34572 24200
rect 37740 24148 37792 24200
rect 16580 24012 16632 24064
rect 31116 24055 31168 24064
rect 31116 24021 31125 24055
rect 31125 24021 31159 24055
rect 31159 24021 31168 24055
rect 31116 24012 31168 24021
rect 38200 24055 38252 24064
rect 38200 24021 38209 24055
rect 38209 24021 38243 24055
rect 38243 24021 38252 24055
rect 38200 24012 38252 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1676 23715 1728 23724
rect 1676 23681 1685 23715
rect 1685 23681 1719 23715
rect 1719 23681 1728 23715
rect 1676 23672 1728 23681
rect 3884 23808 3936 23860
rect 6644 23851 6696 23860
rect 3608 23672 3660 23724
rect 6092 23740 6144 23792
rect 6644 23817 6653 23851
rect 6653 23817 6687 23851
rect 6687 23817 6696 23851
rect 6644 23808 6696 23817
rect 6828 23808 6880 23860
rect 7748 23808 7800 23860
rect 11152 23808 11204 23860
rect 7012 23740 7064 23792
rect 4712 23715 4764 23724
rect 4712 23681 4721 23715
rect 4721 23681 4755 23715
rect 4755 23681 4764 23715
rect 5172 23715 5224 23724
rect 4712 23672 4764 23681
rect 5172 23681 5181 23715
rect 5181 23681 5215 23715
rect 5215 23681 5224 23715
rect 5172 23672 5224 23681
rect 6460 23672 6512 23724
rect 7288 23672 7340 23724
rect 12440 23740 12492 23792
rect 12532 23740 12584 23792
rect 12900 23740 12952 23792
rect 15384 23783 15436 23792
rect 7656 23672 7708 23724
rect 7564 23604 7616 23656
rect 9128 23672 9180 23724
rect 9312 23715 9364 23724
rect 9312 23681 9321 23715
rect 9321 23681 9355 23715
rect 9355 23681 9364 23715
rect 9312 23672 9364 23681
rect 9496 23715 9548 23724
rect 9496 23681 9505 23715
rect 9505 23681 9539 23715
rect 9539 23681 9548 23715
rect 9496 23672 9548 23681
rect 10600 23672 10652 23724
rect 11704 23715 11756 23724
rect 11704 23681 11713 23715
rect 11713 23681 11747 23715
rect 11747 23681 11756 23715
rect 11704 23672 11756 23681
rect 5816 23536 5868 23588
rect 10876 23604 10928 23656
rect 12624 23672 12676 23724
rect 15384 23749 15393 23783
rect 15393 23749 15427 23783
rect 15427 23749 15436 23783
rect 15384 23740 15436 23749
rect 16580 23740 16632 23792
rect 22100 23851 22152 23860
rect 22100 23817 22109 23851
rect 22109 23817 22143 23851
rect 22143 23817 22152 23851
rect 32680 23851 32732 23860
rect 22100 23808 22152 23817
rect 32680 23817 32689 23851
rect 32689 23817 32723 23851
rect 32723 23817 32732 23851
rect 32680 23808 32732 23817
rect 18972 23783 19024 23792
rect 18972 23749 18981 23783
rect 18981 23749 19015 23783
rect 19015 23749 19024 23783
rect 18972 23740 19024 23749
rect 23296 23715 23348 23724
rect 23296 23681 23305 23715
rect 23305 23681 23339 23715
rect 23339 23681 23348 23715
rect 23296 23672 23348 23681
rect 25412 23672 25464 23724
rect 32864 23715 32916 23724
rect 32864 23681 32873 23715
rect 32873 23681 32907 23715
rect 32907 23681 32916 23715
rect 32864 23672 32916 23681
rect 13912 23579 13964 23588
rect 2504 23468 2556 23520
rect 3884 23468 3936 23520
rect 4712 23468 4764 23520
rect 5264 23511 5316 23520
rect 5264 23477 5273 23511
rect 5273 23477 5307 23511
rect 5307 23477 5316 23511
rect 5264 23468 5316 23477
rect 6644 23468 6696 23520
rect 9772 23468 9824 23520
rect 11612 23468 11664 23520
rect 11796 23511 11848 23520
rect 11796 23477 11805 23511
rect 11805 23477 11839 23511
rect 11839 23477 11848 23511
rect 11796 23468 11848 23477
rect 13912 23545 13921 23579
rect 13921 23545 13955 23579
rect 13955 23545 13964 23579
rect 13912 23536 13964 23545
rect 14832 23604 14884 23656
rect 15660 23647 15712 23656
rect 15660 23613 15669 23647
rect 15669 23613 15703 23647
rect 15703 23613 15712 23647
rect 15660 23604 15712 23613
rect 18052 23647 18104 23656
rect 18052 23613 18061 23647
rect 18061 23613 18095 23647
rect 18095 23613 18104 23647
rect 18052 23604 18104 23613
rect 18880 23647 18932 23656
rect 18880 23613 18889 23647
rect 18889 23613 18923 23647
rect 18923 23613 18932 23647
rect 18880 23604 18932 23613
rect 18604 23536 18656 23588
rect 14464 23468 14516 23520
rect 16396 23468 16448 23520
rect 17316 23468 17368 23520
rect 18512 23468 18564 23520
rect 23940 23511 23992 23520
rect 23940 23477 23949 23511
rect 23949 23477 23983 23511
rect 23983 23477 23992 23511
rect 23940 23468 23992 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 6276 23264 6328 23316
rect 3516 23060 3568 23112
rect 4620 23060 4672 23112
rect 6644 23128 6696 23180
rect 9680 23128 9732 23180
rect 1860 23035 1912 23044
rect 1860 23001 1869 23035
rect 1869 23001 1903 23035
rect 1903 23001 1912 23035
rect 1860 22992 1912 23001
rect 3608 22992 3660 23044
rect 3976 22992 4028 23044
rect 6552 23060 6604 23112
rect 7012 23060 7064 23112
rect 7380 23060 7432 23112
rect 7748 23103 7800 23112
rect 7748 23069 7757 23103
rect 7757 23069 7791 23103
rect 7791 23069 7800 23103
rect 7748 23060 7800 23069
rect 8392 23103 8444 23112
rect 8392 23069 8401 23103
rect 8401 23069 8435 23103
rect 8435 23069 8444 23103
rect 8392 23060 8444 23069
rect 11336 23060 11388 23112
rect 13084 23196 13136 23248
rect 13360 23128 13412 23180
rect 16488 23196 16540 23248
rect 16764 23239 16816 23248
rect 16764 23205 16773 23239
rect 16773 23205 16807 23239
rect 16807 23205 16816 23239
rect 16764 23196 16816 23205
rect 14740 23171 14792 23180
rect 14740 23137 14749 23171
rect 14749 23137 14783 23171
rect 14783 23137 14792 23171
rect 14740 23128 14792 23137
rect 17408 23264 17460 23316
rect 18972 23264 19024 23316
rect 17316 23196 17368 23248
rect 18880 23128 18932 23180
rect 15016 23060 15068 23112
rect 7196 22992 7248 23044
rect 9588 23035 9640 23044
rect 9588 23001 9597 23035
rect 9597 23001 9631 23035
rect 9631 23001 9640 23035
rect 9588 22992 9640 23001
rect 1676 22924 1728 22976
rect 4068 22924 4120 22976
rect 4620 22924 4672 22976
rect 7472 22924 7524 22976
rect 7564 22924 7616 22976
rect 9404 22924 9456 22976
rect 11152 22967 11204 22976
rect 11152 22933 11161 22967
rect 11161 22933 11195 22967
rect 11195 22933 11204 22967
rect 11152 22924 11204 22933
rect 12716 22924 12768 22976
rect 14464 23035 14516 23044
rect 14464 23001 14473 23035
rect 14473 23001 14507 23035
rect 14507 23001 14516 23035
rect 17592 23060 17644 23112
rect 18328 23103 18380 23112
rect 18328 23069 18337 23103
rect 18337 23069 18371 23103
rect 18371 23069 18380 23103
rect 18328 23060 18380 23069
rect 16580 23035 16632 23044
rect 14464 22992 14516 23001
rect 16580 23001 16589 23035
rect 16589 23001 16623 23035
rect 16623 23001 16632 23035
rect 16580 22992 16632 23001
rect 17684 23035 17736 23044
rect 17684 23001 17693 23035
rect 17693 23001 17727 23035
rect 17727 23001 17736 23035
rect 17684 22992 17736 23001
rect 18144 22992 18196 23044
rect 19432 22992 19484 23044
rect 15200 22924 15252 22976
rect 18880 22924 18932 22976
rect 22376 22924 22428 22976
rect 22652 22924 22704 22976
rect 25412 23103 25464 23112
rect 25412 23069 25421 23103
rect 25421 23069 25455 23103
rect 25455 23069 25464 23103
rect 25412 23060 25464 23069
rect 37832 23060 37884 23112
rect 27988 22992 28040 23044
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 1860 22720 1912 22772
rect 6736 22720 6788 22772
rect 2688 22652 2740 22704
rect 2872 22695 2924 22704
rect 2872 22661 2881 22695
rect 2881 22661 2915 22695
rect 2915 22661 2924 22695
rect 2872 22652 2924 22661
rect 2964 22695 3016 22704
rect 2964 22661 2973 22695
rect 2973 22661 3007 22695
rect 3007 22661 3016 22695
rect 2964 22652 3016 22661
rect 6460 22652 6512 22704
rect 7472 22695 7524 22704
rect 7472 22661 7481 22695
rect 7481 22661 7515 22695
rect 7515 22661 7524 22695
rect 7472 22652 7524 22661
rect 12072 22720 12124 22772
rect 8484 22652 8536 22704
rect 9680 22652 9732 22704
rect 11060 22652 11112 22704
rect 11796 22652 11848 22704
rect 14648 22720 14700 22772
rect 21456 22652 21508 22704
rect 37832 22720 37884 22772
rect 38016 22720 38068 22772
rect 3608 22516 3660 22568
rect 2228 22491 2280 22500
rect 2228 22457 2237 22491
rect 2237 22457 2271 22491
rect 2271 22457 2280 22491
rect 2228 22448 2280 22457
rect 5080 22584 5132 22636
rect 6736 22627 6788 22636
rect 6736 22593 6745 22627
rect 6745 22593 6779 22627
rect 6779 22593 6788 22627
rect 6736 22584 6788 22593
rect 13268 22584 13320 22636
rect 16028 22584 16080 22636
rect 7748 22516 7800 22568
rect 8852 22516 8904 22568
rect 10324 22516 10376 22568
rect 6276 22448 6328 22500
rect 6460 22448 6512 22500
rect 9588 22448 9640 22500
rect 12072 22516 12124 22568
rect 12256 22559 12308 22568
rect 12256 22525 12265 22559
rect 12265 22525 12299 22559
rect 12299 22525 12308 22559
rect 12256 22516 12308 22525
rect 17316 22516 17368 22568
rect 18880 22559 18932 22568
rect 18880 22525 18889 22559
rect 18889 22525 18923 22559
rect 18923 22525 18932 22559
rect 18880 22516 18932 22525
rect 19156 22516 19208 22568
rect 22192 22516 22244 22568
rect 22376 22559 22428 22568
rect 22376 22525 22385 22559
rect 22385 22525 22419 22559
rect 22419 22525 22428 22559
rect 22376 22516 22428 22525
rect 23296 22516 23348 22568
rect 23848 22584 23900 22636
rect 37832 22584 37884 22636
rect 37924 22516 37976 22568
rect 5172 22380 5224 22432
rect 5816 22380 5868 22432
rect 6644 22380 6696 22432
rect 13820 22423 13872 22432
rect 13820 22389 13829 22423
rect 13829 22389 13863 22423
rect 13863 22389 13872 22423
rect 13820 22380 13872 22389
rect 18512 22448 18564 22500
rect 21364 22491 21416 22500
rect 21364 22457 21373 22491
rect 21373 22457 21407 22491
rect 21407 22457 21416 22491
rect 21364 22448 21416 22457
rect 34796 22448 34848 22500
rect 38200 22491 38252 22500
rect 38200 22457 38209 22491
rect 38209 22457 38243 22491
rect 38243 22457 38252 22491
rect 38200 22448 38252 22457
rect 22192 22380 22244 22432
rect 23204 22380 23256 22432
rect 23756 22423 23808 22432
rect 23756 22389 23765 22423
rect 23765 22389 23799 22423
rect 23799 22389 23808 22423
rect 23756 22380 23808 22389
rect 24768 22380 24820 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3608 22176 3660 22228
rect 16120 22176 16172 22228
rect 17500 22176 17552 22228
rect 17868 22176 17920 22228
rect 7472 22108 7524 22160
rect 8392 22108 8444 22160
rect 2044 22040 2096 22092
rect 2412 22083 2464 22092
rect 2412 22049 2421 22083
rect 2421 22049 2455 22083
rect 2455 22049 2464 22083
rect 2412 22040 2464 22049
rect 4620 22040 4672 22092
rect 4988 22083 5040 22092
rect 4988 22049 4997 22083
rect 4997 22049 5031 22083
rect 5031 22049 5040 22083
rect 4988 22040 5040 22049
rect 5816 22040 5868 22092
rect 6460 22040 6512 22092
rect 7748 22040 7800 22092
rect 11060 22108 11112 22160
rect 12072 22108 12124 22160
rect 9588 22040 9640 22092
rect 4160 21972 4212 22024
rect 4804 21972 4856 22024
rect 8392 22015 8444 22024
rect 8392 21981 8401 22015
rect 8401 21981 8435 22015
rect 8435 21981 8444 22015
rect 8392 21972 8444 21981
rect 2504 21947 2556 21956
rect 2504 21913 2513 21947
rect 2513 21913 2547 21947
rect 2547 21913 2556 21947
rect 2504 21904 2556 21913
rect 3608 21904 3660 21956
rect 4252 21836 4304 21888
rect 4344 21879 4396 21888
rect 4344 21845 4353 21879
rect 4353 21845 4387 21879
rect 4387 21845 4396 21879
rect 5816 21904 5868 21956
rect 9404 21947 9456 21956
rect 4344 21836 4396 21845
rect 5724 21836 5776 21888
rect 9404 21913 9413 21947
rect 9413 21913 9447 21947
rect 9447 21913 9456 21947
rect 9404 21904 9456 21913
rect 9496 21947 9548 21956
rect 9496 21913 9505 21947
rect 9505 21913 9539 21947
rect 9539 21913 9548 21947
rect 9496 21904 9548 21913
rect 7932 21836 7984 21888
rect 9956 21836 10008 21888
rect 11152 21904 11204 21956
rect 11336 21904 11388 21956
rect 12072 21972 12124 22024
rect 11888 21904 11940 21956
rect 17960 22108 18012 22160
rect 22928 22108 22980 22160
rect 14648 22083 14700 22092
rect 14648 22049 14657 22083
rect 14657 22049 14691 22083
rect 14691 22049 14700 22083
rect 14648 22040 14700 22049
rect 12440 21947 12492 21956
rect 12440 21913 12449 21947
rect 12449 21913 12483 21947
rect 12483 21913 12492 21947
rect 12440 21904 12492 21913
rect 12716 21904 12768 21956
rect 13544 21904 13596 21956
rect 14096 21972 14148 22024
rect 13728 21904 13780 21956
rect 23020 21972 23072 22024
rect 23296 21972 23348 22024
rect 38016 22015 38068 22024
rect 38016 21981 38025 22015
rect 38025 21981 38059 22015
rect 38059 21981 38068 22015
rect 38016 21972 38068 21981
rect 18144 21904 18196 21956
rect 15292 21879 15344 21888
rect 15292 21845 15301 21879
rect 15301 21845 15335 21879
rect 15335 21845 15344 21879
rect 15292 21836 15344 21845
rect 22192 21836 22244 21888
rect 23296 21879 23348 21888
rect 23296 21845 23305 21879
rect 23305 21845 23339 21879
rect 23339 21845 23348 21879
rect 23296 21836 23348 21845
rect 37924 21836 37976 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 2504 21632 2556 21684
rect 1952 21564 2004 21616
rect 2044 21564 2096 21616
rect 4160 21564 4212 21616
rect 6736 21607 6788 21616
rect 6736 21573 6745 21607
rect 6745 21573 6779 21607
rect 6779 21573 6788 21607
rect 6736 21564 6788 21573
rect 12440 21632 12492 21684
rect 13176 21632 13228 21684
rect 13452 21632 13504 21684
rect 13544 21632 13596 21684
rect 16304 21632 16356 21684
rect 23204 21632 23256 21684
rect 8944 21564 8996 21616
rect 9680 21564 9732 21616
rect 9956 21607 10008 21616
rect 9956 21573 9965 21607
rect 9965 21573 9999 21607
rect 9999 21573 10008 21607
rect 9956 21564 10008 21573
rect 15016 21564 15068 21616
rect 15660 21564 15712 21616
rect 15936 21564 15988 21616
rect 17500 21607 17552 21616
rect 17500 21573 17509 21607
rect 17509 21573 17543 21607
rect 17543 21573 17552 21607
rect 17500 21564 17552 21573
rect 17592 21607 17644 21616
rect 17592 21573 17601 21607
rect 17601 21573 17635 21607
rect 17635 21573 17644 21607
rect 17592 21564 17644 21573
rect 21548 21564 21600 21616
rect 23112 21607 23164 21616
rect 23112 21573 23121 21607
rect 23121 21573 23155 21607
rect 23155 21573 23164 21607
rect 23112 21564 23164 21573
rect 6368 21496 6420 21548
rect 2228 21428 2280 21480
rect 2412 21471 2464 21480
rect 2412 21437 2421 21471
rect 2421 21437 2455 21471
rect 2455 21437 2464 21471
rect 2412 21428 2464 21437
rect 3608 21471 3660 21480
rect 3608 21437 3617 21471
rect 3617 21437 3651 21471
rect 3651 21437 3660 21471
rect 3608 21428 3660 21437
rect 2872 21360 2924 21412
rect 4804 21428 4856 21480
rect 4252 21360 4304 21412
rect 5080 21403 5132 21412
rect 5080 21369 5089 21403
rect 5089 21369 5123 21403
rect 5123 21369 5132 21403
rect 5080 21360 5132 21369
rect 6460 21428 6512 21480
rect 6828 21428 6880 21480
rect 8116 21428 8168 21480
rect 8208 21360 8260 21412
rect 10968 21539 11020 21548
rect 10968 21505 10977 21539
rect 10977 21505 11011 21539
rect 11011 21505 11020 21539
rect 10968 21496 11020 21505
rect 11336 21496 11388 21548
rect 12440 21539 12492 21548
rect 12440 21505 12449 21539
rect 12449 21505 12483 21539
rect 12483 21505 12492 21539
rect 12440 21496 12492 21505
rect 13176 21496 13228 21548
rect 13728 21539 13780 21548
rect 13728 21505 13737 21539
rect 13737 21505 13771 21539
rect 13771 21505 13780 21539
rect 13728 21496 13780 21505
rect 15844 21539 15896 21548
rect 15844 21505 15853 21539
rect 15853 21505 15887 21539
rect 15887 21505 15896 21539
rect 15844 21496 15896 21505
rect 23020 21496 23072 21548
rect 27068 21496 27120 21548
rect 27988 21539 28040 21548
rect 27988 21505 27997 21539
rect 27997 21505 28031 21539
rect 28031 21505 28040 21539
rect 27988 21496 28040 21505
rect 37372 21564 37424 21616
rect 31392 21496 31444 21548
rect 8852 21428 8904 21480
rect 13636 21428 13688 21480
rect 8944 21360 8996 21412
rect 4804 21292 4856 21344
rect 5816 21292 5868 21344
rect 8760 21292 8812 21344
rect 9588 21360 9640 21412
rect 12256 21360 12308 21412
rect 17316 21428 17368 21480
rect 17684 21428 17736 21480
rect 18052 21428 18104 21480
rect 18880 21428 18932 21480
rect 23756 21428 23808 21480
rect 15016 21360 15068 21412
rect 20168 21360 20220 21412
rect 11704 21292 11756 21344
rect 12532 21335 12584 21344
rect 12532 21301 12541 21335
rect 12541 21301 12575 21335
rect 12575 21301 12584 21335
rect 12532 21292 12584 21301
rect 13728 21292 13780 21344
rect 13912 21292 13964 21344
rect 14004 21292 14056 21344
rect 16304 21292 16356 21344
rect 18696 21292 18748 21344
rect 23112 21292 23164 21344
rect 24492 21335 24544 21344
rect 24492 21301 24501 21335
rect 24501 21301 24535 21335
rect 24535 21301 24544 21335
rect 24492 21292 24544 21301
rect 27804 21335 27856 21344
rect 27804 21301 27813 21335
rect 27813 21301 27847 21335
rect 27847 21301 27856 21335
rect 27804 21292 27856 21301
rect 38200 21335 38252 21344
rect 38200 21301 38209 21335
rect 38209 21301 38243 21335
rect 38243 21301 38252 21335
rect 38200 21292 38252 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1768 21131 1820 21140
rect 1768 21097 1777 21131
rect 1777 21097 1811 21131
rect 1811 21097 1820 21131
rect 1768 21088 1820 21097
rect 3884 21088 3936 21140
rect 8760 21088 8812 21140
rect 9312 21088 9364 21140
rect 15844 21088 15896 21140
rect 17592 21088 17644 21140
rect 3608 21020 3660 21072
rect 3056 20952 3108 21004
rect 4252 20952 4304 21004
rect 4712 20952 4764 21004
rect 5264 20995 5316 21004
rect 5264 20961 5273 20995
rect 5273 20961 5307 20995
rect 5307 20961 5316 20995
rect 5264 20952 5316 20961
rect 5724 21020 5776 21072
rect 6828 21020 6880 21072
rect 13544 21020 13596 21072
rect 13636 21020 13688 21072
rect 7196 20995 7248 21004
rect 7196 20961 7205 20995
rect 7205 20961 7239 20995
rect 7239 20961 7248 20995
rect 7196 20952 7248 20961
rect 9404 20952 9456 21004
rect 9680 20952 9732 21004
rect 10784 20952 10836 21004
rect 12164 20952 12216 21004
rect 12624 20995 12676 21004
rect 12624 20961 12633 20995
rect 12633 20961 12667 20995
rect 12667 20961 12676 20995
rect 12624 20952 12676 20961
rect 13820 20952 13872 21004
rect 15476 21020 15528 21072
rect 16580 21020 16632 21072
rect 21456 21088 21508 21140
rect 31392 21131 31444 21140
rect 31392 21097 31401 21131
rect 31401 21097 31435 21131
rect 31435 21097 31444 21131
rect 31392 21088 31444 21097
rect 38476 21088 38528 21140
rect 23204 21020 23256 21072
rect 6828 20884 6880 20936
rect 9128 20884 9180 20936
rect 13728 20927 13780 20936
rect 13728 20893 13737 20927
rect 13737 20893 13771 20927
rect 13771 20893 13780 20927
rect 13728 20884 13780 20893
rect 14280 20927 14332 20936
rect 14280 20893 14289 20927
rect 14289 20893 14323 20927
rect 14323 20893 14332 20927
rect 14280 20884 14332 20893
rect 14648 20884 14700 20936
rect 14924 20927 14976 20936
rect 14924 20893 14933 20927
rect 14933 20893 14967 20927
rect 14967 20893 14976 20927
rect 14924 20884 14976 20893
rect 15476 20884 15528 20936
rect 2596 20816 2648 20868
rect 2412 20748 2464 20800
rect 4252 20816 4304 20868
rect 4804 20816 4856 20868
rect 5356 20859 5408 20868
rect 5356 20825 5365 20859
rect 5365 20825 5399 20859
rect 5399 20825 5408 20859
rect 5356 20816 5408 20825
rect 7564 20816 7616 20868
rect 8944 20816 8996 20868
rect 3976 20748 4028 20800
rect 6092 20748 6144 20800
rect 6368 20748 6420 20800
rect 9220 20748 9272 20800
rect 9404 20748 9456 20800
rect 10140 20816 10192 20868
rect 11796 20859 11848 20868
rect 11796 20825 11805 20859
rect 11805 20825 11839 20859
rect 11839 20825 11848 20859
rect 11796 20816 11848 20825
rect 13360 20816 13412 20868
rect 20720 20995 20772 21004
rect 20720 20961 20729 20995
rect 20729 20961 20763 20995
rect 20763 20961 20772 20995
rect 20720 20952 20772 20961
rect 16580 20927 16632 20936
rect 16580 20893 16589 20927
rect 16589 20893 16623 20927
rect 16623 20893 16632 20927
rect 16580 20884 16632 20893
rect 16948 20884 17000 20936
rect 19340 20884 19392 20936
rect 20904 20927 20956 20936
rect 20904 20893 20913 20927
rect 20913 20893 20947 20927
rect 20947 20893 20956 20927
rect 20904 20884 20956 20893
rect 13544 20791 13596 20800
rect 13544 20757 13553 20791
rect 13553 20757 13587 20791
rect 13587 20757 13596 20791
rect 13544 20748 13596 20757
rect 15384 20748 15436 20800
rect 16672 20791 16724 20800
rect 16672 20757 16681 20791
rect 16681 20757 16715 20791
rect 16715 20757 16724 20791
rect 16672 20748 16724 20757
rect 17960 20816 18012 20868
rect 22376 20927 22428 20936
rect 22376 20893 22385 20927
rect 22385 20893 22419 20927
rect 22419 20893 22428 20927
rect 22376 20884 22428 20893
rect 21456 20748 21508 20800
rect 38384 20952 38436 21004
rect 26240 20884 26292 20936
rect 37372 20884 37424 20936
rect 38016 20927 38068 20936
rect 38016 20893 38025 20927
rect 38025 20893 38059 20927
rect 38059 20893 38068 20927
rect 38016 20884 38068 20893
rect 35348 20816 35400 20868
rect 24492 20748 24544 20800
rect 24676 20748 24728 20800
rect 38200 20791 38252 20800
rect 38200 20757 38209 20791
rect 38209 20757 38243 20791
rect 38243 20757 38252 20791
rect 38200 20748 38252 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 1584 20544 1636 20596
rect 3700 20544 3752 20596
rect 7104 20544 7156 20596
rect 8024 20544 8076 20596
rect 14004 20544 14056 20596
rect 14648 20544 14700 20596
rect 3332 20519 3384 20528
rect 3332 20485 3341 20519
rect 3341 20485 3375 20519
rect 3375 20485 3384 20519
rect 3332 20476 3384 20485
rect 4804 20476 4856 20528
rect 5172 20476 5224 20528
rect 6000 20519 6052 20528
rect 6000 20485 6009 20519
rect 6009 20485 6043 20519
rect 6043 20485 6052 20519
rect 6000 20476 6052 20485
rect 7012 20519 7064 20528
rect 7012 20485 7021 20519
rect 7021 20485 7055 20519
rect 7055 20485 7064 20519
rect 7012 20476 7064 20485
rect 4160 20408 4212 20460
rect 3056 20340 3108 20392
rect 3332 20340 3384 20392
rect 3700 20204 3752 20256
rect 6184 20272 6236 20324
rect 7104 20340 7156 20392
rect 7748 20476 7800 20528
rect 8208 20519 8260 20528
rect 8208 20485 8217 20519
rect 8217 20485 8251 20519
rect 8251 20485 8260 20519
rect 8208 20476 8260 20485
rect 8392 20476 8444 20528
rect 10324 20519 10376 20528
rect 10324 20485 10333 20519
rect 10333 20485 10367 20519
rect 10367 20485 10376 20519
rect 10324 20476 10376 20485
rect 11888 20519 11940 20528
rect 11888 20485 11897 20519
rect 11897 20485 11931 20519
rect 11931 20485 11940 20519
rect 11888 20476 11940 20485
rect 12532 20476 12584 20528
rect 12992 20476 13044 20528
rect 15200 20519 15252 20528
rect 15200 20485 15209 20519
rect 15209 20485 15243 20519
rect 15243 20485 15252 20519
rect 15200 20476 15252 20485
rect 15936 20544 15988 20596
rect 8760 20451 8812 20460
rect 8760 20417 8769 20451
rect 8769 20417 8803 20451
rect 8803 20417 8812 20451
rect 8760 20408 8812 20417
rect 7932 20340 7984 20392
rect 7748 20272 7800 20324
rect 8852 20340 8904 20392
rect 10784 20408 10836 20460
rect 12808 20408 12860 20460
rect 13268 20408 13320 20460
rect 13544 20408 13596 20460
rect 16304 20476 16356 20528
rect 16396 20476 16448 20528
rect 19524 20519 19576 20528
rect 19524 20485 19533 20519
rect 19533 20485 19567 20519
rect 19567 20485 19576 20519
rect 19524 20476 19576 20485
rect 20904 20544 20956 20596
rect 22376 20544 22428 20596
rect 37740 20587 37792 20596
rect 37740 20553 37749 20587
rect 37749 20553 37783 20587
rect 37783 20553 37792 20587
rect 37740 20544 37792 20553
rect 9312 20383 9364 20392
rect 9312 20349 9321 20383
rect 9321 20349 9355 20383
rect 9355 20349 9364 20383
rect 9312 20340 9364 20349
rect 9680 20340 9732 20392
rect 9496 20204 9548 20256
rect 13912 20340 13964 20392
rect 12716 20272 12768 20324
rect 13360 20272 13412 20324
rect 16672 20272 16724 20324
rect 18696 20408 18748 20460
rect 19340 20408 19392 20460
rect 17316 20383 17368 20392
rect 17316 20349 17325 20383
rect 17325 20349 17359 20383
rect 17359 20349 17368 20383
rect 17316 20340 17368 20349
rect 18144 20383 18196 20392
rect 18144 20349 18153 20383
rect 18153 20349 18187 20383
rect 18187 20349 18196 20383
rect 18144 20340 18196 20349
rect 17408 20272 17460 20324
rect 17592 20272 17644 20324
rect 22192 20451 22244 20460
rect 22192 20417 22201 20451
rect 22201 20417 22235 20451
rect 22235 20417 22244 20451
rect 22192 20408 22244 20417
rect 27804 20451 27856 20460
rect 27804 20417 27813 20451
rect 27813 20417 27847 20451
rect 27847 20417 27856 20451
rect 27804 20408 27856 20417
rect 35348 20451 35400 20460
rect 35348 20417 35357 20451
rect 35357 20417 35391 20451
rect 35391 20417 35400 20451
rect 38108 20476 38160 20528
rect 35348 20408 35400 20417
rect 36820 20408 36872 20460
rect 22376 20340 22428 20392
rect 19708 20272 19760 20324
rect 31116 20272 31168 20324
rect 16856 20204 16908 20256
rect 17224 20204 17276 20256
rect 22560 20204 22612 20256
rect 26792 20204 26844 20256
rect 34796 20204 34848 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2872 20000 2924 20052
rect 3976 20000 4028 20052
rect 4068 20000 4120 20052
rect 4528 20000 4580 20052
rect 7196 20000 7248 20052
rect 7748 20000 7800 20052
rect 8208 20000 8260 20052
rect 11888 20000 11940 20052
rect 17224 20000 17276 20052
rect 17408 20000 17460 20052
rect 18880 20000 18932 20052
rect 38016 20000 38068 20052
rect 8760 19932 8812 19984
rect 12992 19932 13044 19984
rect 2136 19864 2188 19916
rect 3608 19864 3660 19916
rect 4160 19864 4212 19916
rect 6736 19907 6788 19916
rect 6736 19873 6745 19907
rect 6745 19873 6779 19907
rect 6779 19873 6788 19907
rect 6736 19864 6788 19873
rect 7564 19864 7616 19916
rect 9864 19907 9916 19916
rect 9864 19873 9873 19907
rect 9873 19873 9907 19907
rect 9907 19873 9916 19907
rect 9864 19864 9916 19873
rect 20444 19932 20496 19984
rect 20628 19932 20680 19984
rect 13268 19907 13320 19916
rect 13268 19873 13277 19907
rect 13277 19873 13311 19907
rect 13311 19873 13320 19907
rect 13268 19864 13320 19873
rect 14004 19864 14056 19916
rect 1860 19771 1912 19780
rect 1860 19737 1869 19771
rect 1869 19737 1903 19771
rect 1903 19737 1912 19771
rect 1860 19728 1912 19737
rect 3608 19728 3660 19780
rect 5724 19796 5776 19848
rect 6184 19796 6236 19848
rect 9128 19839 9180 19848
rect 9128 19805 9137 19839
rect 9137 19805 9171 19839
rect 9171 19805 9180 19839
rect 9128 19796 9180 19805
rect 16212 19796 16264 19848
rect 18696 19864 18748 19916
rect 20812 19864 20864 19916
rect 22468 19907 22520 19916
rect 22468 19873 22477 19907
rect 22477 19873 22511 19907
rect 22511 19873 22520 19907
rect 22468 19864 22520 19873
rect 22652 19907 22704 19916
rect 22652 19873 22661 19907
rect 22661 19873 22695 19907
rect 22695 19873 22704 19907
rect 22652 19864 22704 19873
rect 24952 19907 25004 19916
rect 24952 19873 24961 19907
rect 24961 19873 24995 19907
rect 24995 19873 25004 19907
rect 24952 19864 25004 19873
rect 26792 19907 26844 19916
rect 26792 19873 26801 19907
rect 26801 19873 26835 19907
rect 26835 19873 26844 19907
rect 26792 19864 26844 19873
rect 20168 19839 20220 19848
rect 20168 19805 20177 19839
rect 20177 19805 20211 19839
rect 20211 19805 20220 19839
rect 20168 19796 20220 19805
rect 34520 19796 34572 19848
rect 4068 19728 4120 19780
rect 4896 19728 4948 19780
rect 5080 19771 5132 19780
rect 5080 19737 5089 19771
rect 5089 19737 5123 19771
rect 5123 19737 5132 19771
rect 5080 19728 5132 19737
rect 5356 19728 5408 19780
rect 6460 19728 6512 19780
rect 5264 19660 5316 19712
rect 7748 19728 7800 19780
rect 8024 19771 8076 19780
rect 8024 19737 8033 19771
rect 8033 19737 8067 19771
rect 8067 19737 8076 19771
rect 8024 19728 8076 19737
rect 9680 19728 9732 19780
rect 9220 19660 9272 19712
rect 10968 19728 11020 19780
rect 9864 19660 9916 19712
rect 10876 19660 10928 19712
rect 12256 19728 12308 19780
rect 12532 19728 12584 19780
rect 13360 19728 13412 19780
rect 14372 19771 14424 19780
rect 14372 19737 14381 19771
rect 14381 19737 14415 19771
rect 14415 19737 14424 19771
rect 14372 19728 14424 19737
rect 15016 19771 15068 19780
rect 13820 19660 13872 19712
rect 15016 19737 15025 19771
rect 15025 19737 15059 19771
rect 15059 19737 15068 19771
rect 15016 19728 15068 19737
rect 15108 19728 15160 19780
rect 15292 19660 15344 19712
rect 15568 19703 15620 19712
rect 15568 19669 15577 19703
rect 15577 19669 15611 19703
rect 15611 19669 15620 19703
rect 15568 19660 15620 19669
rect 16488 19728 16540 19780
rect 16580 19728 16632 19780
rect 19984 19728 20036 19780
rect 16764 19660 16816 19712
rect 17040 19660 17092 19712
rect 21088 19771 21140 19780
rect 21088 19737 21097 19771
rect 21097 19737 21131 19771
rect 21131 19737 21140 19771
rect 21088 19728 21140 19737
rect 24400 19728 24452 19780
rect 24676 19771 24728 19780
rect 24676 19737 24685 19771
rect 24685 19737 24719 19771
rect 24719 19737 24728 19771
rect 24676 19728 24728 19737
rect 24768 19771 24820 19780
rect 24768 19737 24777 19771
rect 24777 19737 24811 19771
rect 24811 19737 24820 19771
rect 24768 19728 24820 19737
rect 22560 19660 22612 19712
rect 23940 19660 23992 19712
rect 24584 19660 24636 19712
rect 27252 19703 27304 19712
rect 27252 19669 27261 19703
rect 27261 19669 27295 19703
rect 27295 19669 27304 19703
rect 27252 19660 27304 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 3056 19456 3108 19508
rect 2780 19388 2832 19440
rect 3148 19388 3200 19440
rect 7012 19456 7064 19508
rect 5172 19388 5224 19440
rect 5448 19431 5500 19440
rect 5448 19397 5457 19431
rect 5457 19397 5491 19431
rect 5491 19397 5500 19431
rect 5448 19388 5500 19397
rect 6000 19431 6052 19440
rect 6000 19397 6009 19431
rect 6009 19397 6043 19431
rect 6043 19397 6052 19431
rect 6000 19388 6052 19397
rect 6460 19388 6512 19440
rect 4896 19320 4948 19372
rect 10416 19456 10468 19508
rect 7380 19431 7432 19440
rect 7380 19397 7389 19431
rect 7389 19397 7423 19431
rect 7423 19397 7432 19431
rect 7380 19388 7432 19397
rect 9036 19431 9088 19440
rect 9036 19397 9045 19431
rect 9045 19397 9079 19431
rect 9079 19397 9088 19431
rect 9036 19388 9088 19397
rect 9496 19388 9548 19440
rect 13360 19456 13412 19508
rect 11060 19363 11112 19372
rect 11060 19329 11069 19363
rect 11069 19329 11103 19363
rect 11103 19329 11112 19363
rect 11060 19320 11112 19329
rect 2964 19252 3016 19304
rect 3884 19252 3936 19304
rect 5080 19252 5132 19304
rect 5356 19295 5408 19304
rect 5356 19261 5365 19295
rect 5365 19261 5399 19295
rect 5399 19261 5408 19295
rect 5356 19252 5408 19261
rect 5724 19252 5776 19304
rect 6828 19252 6880 19304
rect 7472 19252 7524 19304
rect 8760 19295 8812 19304
rect 8760 19261 8769 19295
rect 8769 19261 8803 19295
rect 8803 19261 8812 19295
rect 8760 19252 8812 19261
rect 2228 19184 2280 19236
rect 3976 19184 4028 19236
rect 10324 19252 10376 19304
rect 10692 19252 10744 19304
rect 11980 19388 12032 19440
rect 12072 19388 12124 19440
rect 14280 19456 14332 19508
rect 13084 19320 13136 19372
rect 13452 19320 13504 19372
rect 12072 19252 12124 19304
rect 12808 19252 12860 19304
rect 17408 19456 17460 19508
rect 15568 19431 15620 19440
rect 13912 19295 13964 19304
rect 13912 19261 13921 19295
rect 13921 19261 13955 19295
rect 13955 19261 13964 19295
rect 13912 19252 13964 19261
rect 14372 19295 14424 19304
rect 14372 19261 14381 19295
rect 14381 19261 14415 19295
rect 14415 19261 14424 19295
rect 14372 19252 14424 19261
rect 12348 19184 12400 19236
rect 15200 19252 15252 19304
rect 15568 19397 15577 19431
rect 15577 19397 15611 19431
rect 15611 19397 15620 19431
rect 15568 19388 15620 19397
rect 17040 19431 17092 19440
rect 17040 19397 17049 19431
rect 17049 19397 17083 19431
rect 17083 19397 17092 19431
rect 17040 19388 17092 19397
rect 20352 19456 20404 19508
rect 20444 19456 20496 19508
rect 23112 19456 23164 19508
rect 36820 19499 36872 19508
rect 16672 19320 16724 19372
rect 20444 19320 20496 19372
rect 24124 19363 24176 19372
rect 24124 19329 24133 19363
rect 24133 19329 24167 19363
rect 24167 19329 24176 19363
rect 24124 19320 24176 19329
rect 17316 19295 17368 19304
rect 14832 19184 14884 19236
rect 17316 19261 17325 19295
rect 17325 19261 17359 19295
rect 17359 19261 17368 19295
rect 17316 19252 17368 19261
rect 20352 19252 20404 19304
rect 20628 19252 20680 19304
rect 24676 19252 24728 19304
rect 36820 19465 36829 19499
rect 36829 19465 36863 19499
rect 36863 19465 36872 19499
rect 36820 19456 36872 19465
rect 37832 19499 37884 19508
rect 37832 19465 37841 19499
rect 37841 19465 37875 19499
rect 37875 19465 37884 19499
rect 37832 19456 37884 19465
rect 27712 19320 27764 19372
rect 38016 19363 38068 19372
rect 38016 19329 38025 19363
rect 38025 19329 38059 19363
rect 38059 19329 38068 19363
rect 38016 19320 38068 19329
rect 16856 19184 16908 19236
rect 23204 19184 23256 19236
rect 26240 19184 26292 19236
rect 4068 19116 4120 19168
rect 6552 19116 6604 19168
rect 6644 19116 6696 19168
rect 10232 19116 10284 19168
rect 10508 19159 10560 19168
rect 10508 19125 10517 19159
rect 10517 19125 10551 19159
rect 10551 19125 10560 19159
rect 10508 19116 10560 19125
rect 10968 19116 11020 19168
rect 17224 19116 17276 19168
rect 17960 19116 18012 19168
rect 18420 19116 18472 19168
rect 19248 19116 19300 19168
rect 23480 19116 23532 19168
rect 24860 19116 24912 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 5356 18912 5408 18964
rect 5448 18912 5500 18964
rect 7288 18912 7340 18964
rect 7748 18912 7800 18964
rect 2964 18844 3016 18896
rect 3240 18776 3292 18828
rect 5172 18776 5224 18828
rect 6000 18776 6052 18828
rect 6552 18844 6604 18896
rect 7196 18844 7248 18896
rect 7472 18844 7524 18896
rect 10048 18912 10100 18964
rect 10140 18912 10192 18964
rect 11428 18912 11480 18964
rect 11888 18912 11940 18964
rect 12256 18912 12308 18964
rect 17684 18912 17736 18964
rect 21548 18955 21600 18964
rect 21548 18921 21557 18955
rect 21557 18921 21591 18955
rect 21591 18921 21600 18955
rect 21548 18912 21600 18921
rect 4252 18751 4304 18760
rect 4252 18717 4261 18751
rect 4261 18717 4295 18751
rect 4295 18717 4304 18751
rect 4252 18708 4304 18717
rect 6368 18708 6420 18760
rect 2320 18683 2372 18692
rect 2320 18649 2329 18683
rect 2329 18649 2363 18683
rect 2363 18649 2372 18683
rect 2320 18640 2372 18649
rect 4160 18640 4212 18692
rect 1492 18572 1544 18624
rect 5080 18683 5132 18692
rect 5080 18649 5089 18683
rect 5089 18649 5123 18683
rect 5123 18649 5132 18683
rect 8576 18776 8628 18828
rect 13176 18844 13228 18896
rect 14740 18844 14792 18896
rect 26240 18912 26292 18964
rect 23940 18844 23992 18896
rect 38568 18912 38620 18964
rect 38200 18844 38252 18896
rect 11520 18819 11572 18828
rect 11520 18785 11529 18819
rect 11529 18785 11563 18819
rect 11563 18785 11572 18819
rect 11520 18776 11572 18785
rect 12256 18776 12308 18828
rect 12532 18776 12584 18828
rect 12992 18776 13044 18828
rect 13084 18776 13136 18828
rect 13544 18819 13596 18828
rect 13544 18785 13553 18819
rect 13553 18785 13587 18819
rect 13587 18785 13596 18819
rect 13544 18776 13596 18785
rect 15844 18776 15896 18828
rect 21548 18776 21600 18828
rect 24676 18819 24728 18828
rect 24676 18785 24685 18819
rect 24685 18785 24719 18819
rect 24719 18785 24728 18819
rect 24676 18776 24728 18785
rect 5080 18640 5132 18649
rect 7012 18640 7064 18692
rect 7288 18640 7340 18692
rect 7472 18640 7524 18692
rect 8024 18640 8076 18692
rect 8852 18708 8904 18760
rect 12348 18708 12400 18760
rect 13912 18708 13964 18760
rect 16212 18708 16264 18760
rect 16672 18708 16724 18760
rect 16948 18751 17000 18760
rect 16948 18717 16957 18751
rect 16957 18717 16991 18751
rect 16991 18717 17000 18751
rect 16948 18708 17000 18717
rect 9404 18640 9456 18692
rect 9864 18640 9916 18692
rect 12808 18683 12860 18692
rect 12808 18649 12817 18683
rect 12817 18649 12851 18683
rect 12851 18649 12860 18683
rect 12808 18640 12860 18649
rect 13636 18640 13688 18692
rect 15384 18683 15436 18692
rect 8300 18572 8352 18624
rect 10048 18572 10100 18624
rect 10324 18572 10376 18624
rect 10876 18572 10928 18624
rect 11428 18572 11480 18624
rect 11520 18572 11572 18624
rect 12256 18572 12308 18624
rect 14464 18615 14516 18624
rect 14464 18581 14473 18615
rect 14473 18581 14507 18615
rect 14507 18581 14516 18615
rect 14464 18572 14516 18581
rect 15384 18649 15393 18683
rect 15393 18649 15427 18683
rect 15427 18649 15436 18683
rect 15384 18640 15436 18649
rect 15476 18683 15528 18692
rect 15476 18649 15485 18683
rect 15485 18649 15519 18683
rect 15519 18649 15528 18683
rect 17960 18708 18012 18760
rect 18144 18708 18196 18760
rect 18420 18708 18472 18760
rect 20260 18708 20312 18760
rect 26240 18708 26292 18760
rect 27988 18708 28040 18760
rect 37464 18708 37516 18760
rect 38292 18751 38344 18760
rect 38292 18717 38301 18751
rect 38301 18717 38335 18751
rect 38335 18717 38344 18751
rect 38292 18708 38344 18717
rect 15476 18640 15528 18649
rect 17224 18640 17276 18692
rect 23480 18683 23532 18692
rect 23480 18649 23489 18683
rect 23489 18649 23523 18683
rect 23523 18649 23532 18683
rect 23480 18640 23532 18649
rect 17040 18615 17092 18624
rect 17040 18581 17049 18615
rect 17049 18581 17083 18615
rect 17083 18581 17092 18615
rect 17040 18572 17092 18581
rect 17408 18572 17460 18624
rect 18420 18572 18472 18624
rect 23940 18572 23992 18624
rect 24860 18640 24912 18692
rect 34520 18640 34572 18692
rect 27344 18572 27396 18624
rect 38108 18615 38160 18624
rect 38108 18581 38117 18615
rect 38117 18581 38151 18615
rect 38151 18581 38160 18615
rect 38108 18572 38160 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 1676 18368 1728 18420
rect 4712 18368 4764 18420
rect 5264 18368 5316 18420
rect 3976 18300 4028 18352
rect 5172 18300 5224 18352
rect 1860 18275 1912 18284
rect 1860 18241 1869 18275
rect 1869 18241 1903 18275
rect 1903 18241 1912 18275
rect 1860 18232 1912 18241
rect 5080 18275 5132 18284
rect 5080 18241 5089 18275
rect 5089 18241 5123 18275
rect 5123 18241 5132 18275
rect 5080 18232 5132 18241
rect 3332 18164 3384 18216
rect 2964 18096 3016 18148
rect 4068 18164 4120 18216
rect 5724 18164 5776 18216
rect 6920 18368 6972 18420
rect 8760 18368 8812 18420
rect 15476 18368 15528 18420
rect 19984 18368 20036 18420
rect 10876 18300 10928 18352
rect 11888 18343 11940 18352
rect 11888 18309 11897 18343
rect 11897 18309 11931 18343
rect 11931 18309 11940 18343
rect 11888 18300 11940 18309
rect 12992 18300 13044 18352
rect 13544 18343 13596 18352
rect 13544 18309 13553 18343
rect 13553 18309 13587 18343
rect 13587 18309 13596 18343
rect 13544 18300 13596 18309
rect 13636 18300 13688 18352
rect 10324 18232 10376 18284
rect 15200 18275 15252 18284
rect 6644 18207 6696 18216
rect 6644 18173 6653 18207
rect 6653 18173 6687 18207
rect 6687 18173 6696 18207
rect 6644 18164 6696 18173
rect 1768 18028 1820 18080
rect 6552 18096 6604 18148
rect 4160 18028 4212 18080
rect 4804 18028 4856 18080
rect 7748 18096 7800 18148
rect 8668 18164 8720 18216
rect 10048 18164 10100 18216
rect 13084 18164 13136 18216
rect 14372 18207 14424 18216
rect 9680 18096 9732 18148
rect 10968 18096 11020 18148
rect 11428 18096 11480 18148
rect 11612 18096 11664 18148
rect 13360 18096 13412 18148
rect 14372 18173 14381 18207
rect 14381 18173 14415 18207
rect 14415 18173 14424 18207
rect 14372 18164 14424 18173
rect 14832 18164 14884 18216
rect 15200 18241 15209 18275
rect 15209 18241 15243 18275
rect 15243 18241 15252 18275
rect 15200 18232 15252 18241
rect 16212 18300 16264 18352
rect 17040 18300 17092 18352
rect 36360 18368 36412 18420
rect 38016 18368 38068 18420
rect 16488 18232 16540 18284
rect 16580 18232 16632 18284
rect 22284 18300 22336 18352
rect 20076 18232 20128 18284
rect 22100 18207 22152 18216
rect 22100 18173 22109 18207
rect 22109 18173 22143 18207
rect 22143 18173 22152 18207
rect 22100 18164 22152 18173
rect 21456 18096 21508 18148
rect 23204 18300 23256 18352
rect 27252 18300 27304 18352
rect 25136 18232 25188 18284
rect 27344 18275 27396 18284
rect 27344 18241 27353 18275
rect 27353 18241 27387 18275
rect 27387 18241 27396 18275
rect 27344 18232 27396 18241
rect 38108 18232 38160 18284
rect 38292 18275 38344 18284
rect 38292 18241 38301 18275
rect 38301 18241 38335 18275
rect 38335 18241 38344 18275
rect 38292 18232 38344 18241
rect 23756 18207 23808 18216
rect 23756 18173 23765 18207
rect 23765 18173 23799 18207
rect 23799 18173 23808 18207
rect 23756 18164 23808 18173
rect 7472 18028 7524 18080
rect 12164 18028 12216 18080
rect 13544 18028 13596 18080
rect 17684 18028 17736 18080
rect 24952 18164 25004 18216
rect 27160 18207 27212 18216
rect 27160 18173 27169 18207
rect 27169 18173 27203 18207
rect 27203 18173 27212 18207
rect 27160 18164 27212 18173
rect 26240 18028 26292 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 4620 17824 4672 17876
rect 4988 17824 5040 17876
rect 11428 17824 11480 17876
rect 8760 17756 8812 17808
rect 10876 17756 10928 17808
rect 12532 17824 12584 17876
rect 12624 17824 12676 17876
rect 1584 17663 1636 17672
rect 1584 17629 1593 17663
rect 1593 17629 1627 17663
rect 1627 17629 1636 17663
rect 1584 17620 1636 17629
rect 7104 17688 7156 17740
rect 12164 17688 12216 17740
rect 12532 17688 12584 17740
rect 14096 17756 14148 17808
rect 16120 17756 16172 17808
rect 20996 17824 21048 17876
rect 21180 17824 21232 17876
rect 24124 17824 24176 17876
rect 13820 17688 13872 17740
rect 14556 17688 14608 17740
rect 20812 17688 20864 17740
rect 22376 17756 22428 17808
rect 6828 17663 6880 17672
rect 1860 17595 1912 17604
rect 1860 17561 1869 17595
rect 1869 17561 1903 17595
rect 1903 17561 1912 17595
rect 1860 17552 1912 17561
rect 4252 17595 4304 17604
rect 4252 17561 4261 17595
rect 4261 17561 4295 17595
rect 4295 17561 4304 17595
rect 4252 17552 4304 17561
rect 4712 17552 4764 17604
rect 6000 17552 6052 17604
rect 6828 17629 6837 17663
rect 6837 17629 6871 17663
rect 6871 17629 6880 17663
rect 6828 17620 6880 17629
rect 8852 17620 8904 17672
rect 10876 17620 10928 17672
rect 11152 17620 11204 17672
rect 11796 17663 11848 17672
rect 11796 17629 11805 17663
rect 11805 17629 11839 17663
rect 11839 17629 11848 17663
rect 11796 17620 11848 17629
rect 14280 17663 14332 17672
rect 14280 17629 14289 17663
rect 14289 17629 14323 17663
rect 14323 17629 14332 17663
rect 17316 17663 17368 17672
rect 14280 17620 14332 17629
rect 17316 17629 17325 17663
rect 17325 17629 17359 17663
rect 17359 17629 17368 17663
rect 17316 17620 17368 17629
rect 17500 17620 17552 17672
rect 22008 17663 22060 17672
rect 22008 17629 22017 17663
rect 22017 17629 22051 17663
rect 22051 17629 22060 17663
rect 22008 17620 22060 17629
rect 6736 17552 6788 17604
rect 4068 17484 4120 17536
rect 7564 17552 7616 17604
rect 10048 17552 10100 17604
rect 12348 17552 12400 17604
rect 13360 17552 13412 17604
rect 15016 17595 15068 17604
rect 15016 17561 15025 17595
rect 15025 17561 15059 17595
rect 15059 17561 15068 17595
rect 15016 17552 15068 17561
rect 16212 17595 16264 17604
rect 10692 17484 10744 17536
rect 11152 17484 11204 17536
rect 13084 17484 13136 17536
rect 13636 17484 13688 17536
rect 16212 17561 16221 17595
rect 16221 17561 16255 17595
rect 16255 17561 16264 17595
rect 16212 17552 16264 17561
rect 16304 17595 16356 17604
rect 16304 17561 16313 17595
rect 16313 17561 16347 17595
rect 16347 17561 16356 17595
rect 16304 17552 16356 17561
rect 17132 17552 17184 17604
rect 17684 17552 17736 17604
rect 19892 17552 19944 17604
rect 19984 17595 20036 17604
rect 19984 17561 19993 17595
rect 19993 17561 20027 17595
rect 20027 17561 20036 17595
rect 19984 17552 20036 17561
rect 20168 17552 20220 17604
rect 20628 17552 20680 17604
rect 22928 17663 22980 17672
rect 22928 17629 22937 17663
rect 22937 17629 22971 17663
rect 22971 17629 22980 17663
rect 22928 17620 22980 17629
rect 28264 17620 28316 17672
rect 30564 17595 30616 17604
rect 30564 17561 30573 17595
rect 30573 17561 30607 17595
rect 30607 17561 30616 17595
rect 30564 17552 30616 17561
rect 27344 17484 27396 17536
rect 37832 17484 37884 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 1952 17280 2004 17332
rect 3700 17323 3752 17332
rect 2872 17212 2924 17264
rect 3700 17289 3709 17323
rect 3709 17289 3743 17323
rect 3743 17289 3752 17323
rect 3700 17280 3752 17289
rect 8484 17280 8536 17332
rect 8668 17280 8720 17332
rect 10048 17280 10100 17332
rect 12164 17280 12216 17332
rect 16212 17280 16264 17332
rect 16488 17280 16540 17332
rect 16672 17280 16724 17332
rect 19984 17280 20036 17332
rect 4620 17212 4672 17264
rect 5540 17212 5592 17264
rect 7840 17212 7892 17264
rect 11060 17212 11112 17264
rect 11152 17212 11204 17264
rect 12256 17212 12308 17264
rect 13820 17212 13872 17264
rect 14556 17255 14608 17264
rect 14556 17221 14565 17255
rect 14565 17221 14599 17255
rect 14599 17221 14608 17255
rect 14556 17212 14608 17221
rect 16856 17212 16908 17264
rect 6552 17187 6604 17196
rect 6552 17153 6561 17187
rect 6561 17153 6595 17187
rect 6595 17153 6604 17187
rect 6552 17144 6604 17153
rect 10600 17144 10652 17196
rect 11796 17144 11848 17196
rect 1584 17076 1636 17128
rect 4068 17076 4120 17128
rect 3976 17008 4028 17060
rect 6920 17076 6972 17128
rect 8852 17119 8904 17128
rect 8852 17085 8861 17119
rect 8861 17085 8895 17119
rect 8895 17085 8904 17119
rect 8852 17076 8904 17085
rect 10140 17076 10192 17128
rect 10232 17008 10284 17060
rect 10692 17008 10744 17060
rect 17776 17212 17828 17264
rect 17500 17144 17552 17196
rect 13728 17119 13780 17128
rect 13728 17085 13737 17119
rect 13737 17085 13771 17119
rect 13771 17085 13780 17119
rect 13728 17076 13780 17085
rect 14556 17076 14608 17128
rect 17316 17076 17368 17128
rect 6276 16940 6328 16992
rect 6920 16940 6972 16992
rect 7472 16940 7524 16992
rect 8484 16940 8536 16992
rect 14280 16940 14332 16992
rect 15660 17008 15712 17060
rect 16948 17008 17000 17060
rect 16120 16940 16172 16992
rect 16488 16940 16540 16992
rect 19432 17212 19484 17264
rect 20536 17212 20588 17264
rect 22928 17212 22980 17264
rect 19708 17144 19760 17196
rect 19524 17008 19576 17060
rect 19340 16940 19392 16992
rect 20168 17008 20220 17060
rect 19708 16940 19760 16992
rect 22376 17119 22428 17128
rect 22376 17085 22385 17119
rect 22385 17085 22419 17119
rect 22419 17085 22428 17119
rect 22376 17076 22428 17085
rect 27160 17280 27212 17332
rect 28264 17323 28316 17332
rect 28264 17289 28273 17323
rect 28273 17289 28307 17323
rect 28307 17289 28316 17323
rect 28264 17280 28316 17289
rect 27344 17187 27396 17196
rect 27344 17153 27353 17187
rect 27353 17153 27387 17187
rect 27387 17153 27396 17187
rect 27344 17144 27396 17153
rect 28448 17187 28500 17196
rect 28448 17153 28457 17187
rect 28457 17153 28491 17187
rect 28491 17153 28500 17187
rect 28448 17144 28500 17153
rect 27252 17076 27304 17128
rect 24400 16940 24452 16992
rect 27620 16983 27672 16992
rect 27620 16949 27629 16983
rect 27629 16949 27663 16983
rect 27663 16949 27672 16983
rect 27620 16940 27672 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 3240 16736 3292 16788
rect 3976 16736 4028 16788
rect 4988 16736 5040 16788
rect 7748 16736 7800 16788
rect 8668 16736 8720 16788
rect 3424 16600 3476 16652
rect 4252 16600 4304 16652
rect 6552 16600 6604 16652
rect 9220 16668 9272 16720
rect 9404 16668 9456 16720
rect 10692 16668 10744 16720
rect 12072 16668 12124 16720
rect 13176 16736 13228 16788
rect 13728 16736 13780 16788
rect 15016 16736 15068 16788
rect 15660 16736 15712 16788
rect 16304 16736 16356 16788
rect 8852 16600 8904 16652
rect 11336 16600 11388 16652
rect 14096 16668 14148 16720
rect 17868 16668 17920 16720
rect 22376 16736 22428 16788
rect 18972 16668 19024 16720
rect 1584 16575 1636 16584
rect 1584 16541 1593 16575
rect 1593 16541 1627 16575
rect 1627 16541 1636 16575
rect 1584 16532 1636 16541
rect 4528 16532 4580 16584
rect 6828 16575 6880 16584
rect 6828 16541 6837 16575
rect 6837 16541 6871 16575
rect 6871 16541 6880 16575
rect 6828 16532 6880 16541
rect 9312 16532 9364 16584
rect 3792 16464 3844 16516
rect 4620 16464 4672 16516
rect 5632 16464 5684 16516
rect 4068 16439 4120 16448
rect 4068 16405 4077 16439
rect 4077 16405 4111 16439
rect 4111 16405 4120 16439
rect 4068 16396 4120 16405
rect 5080 16396 5132 16448
rect 6368 16439 6420 16448
rect 6368 16405 6377 16439
rect 6377 16405 6411 16439
rect 6411 16405 6420 16439
rect 6368 16396 6420 16405
rect 7656 16464 7708 16516
rect 9680 16464 9732 16516
rect 10600 16532 10652 16584
rect 12440 16532 12492 16584
rect 14556 16600 14608 16652
rect 15752 16600 15804 16652
rect 15936 16600 15988 16652
rect 20076 16600 20128 16652
rect 20168 16600 20220 16652
rect 20444 16600 20496 16652
rect 20720 16600 20772 16652
rect 22008 16600 22060 16652
rect 24584 16643 24636 16652
rect 14280 16575 14332 16584
rect 14280 16541 14289 16575
rect 14289 16541 14323 16575
rect 14323 16541 14332 16575
rect 14280 16532 14332 16541
rect 16212 16532 16264 16584
rect 16672 16532 16724 16584
rect 16948 16575 17000 16584
rect 16948 16541 16957 16575
rect 16957 16541 16991 16575
rect 16991 16541 17000 16575
rect 17500 16575 17552 16584
rect 16948 16532 17000 16541
rect 17500 16541 17509 16575
rect 17509 16541 17543 16575
rect 17543 16541 17552 16575
rect 17500 16532 17552 16541
rect 18604 16532 18656 16584
rect 19340 16532 19392 16584
rect 24584 16609 24593 16643
rect 24593 16609 24627 16643
rect 24627 16609 24636 16643
rect 24584 16600 24636 16609
rect 26148 16600 26200 16652
rect 27620 16532 27672 16584
rect 38016 16575 38068 16584
rect 38016 16541 38025 16575
rect 38025 16541 38059 16575
rect 38059 16541 38068 16575
rect 38016 16532 38068 16541
rect 10968 16464 11020 16516
rect 12256 16464 12308 16516
rect 12808 16464 12860 16516
rect 14648 16464 14700 16516
rect 16304 16464 16356 16516
rect 19708 16464 19760 16516
rect 20444 16464 20496 16516
rect 8576 16439 8628 16448
rect 8576 16405 8585 16439
rect 8585 16405 8619 16439
rect 8619 16405 8628 16439
rect 8576 16396 8628 16405
rect 11060 16396 11112 16448
rect 11152 16396 11204 16448
rect 11980 16396 12032 16448
rect 12532 16396 12584 16448
rect 15936 16396 15988 16448
rect 18696 16396 18748 16448
rect 19524 16396 19576 16448
rect 28632 16464 28684 16516
rect 22560 16439 22612 16448
rect 22560 16405 22569 16439
rect 22569 16405 22603 16439
rect 22603 16405 22612 16439
rect 22560 16396 22612 16405
rect 38200 16439 38252 16448
rect 38200 16405 38209 16439
rect 38209 16405 38243 16439
rect 38243 16405 38252 16439
rect 38200 16396 38252 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 1124 16192 1176 16244
rect 4620 16124 4672 16176
rect 5540 16192 5592 16244
rect 6092 16192 6144 16244
rect 6368 16192 6420 16244
rect 8392 16192 8444 16244
rect 11612 16192 11664 16244
rect 13360 16192 13412 16244
rect 4252 16099 4304 16108
rect 1584 15988 1636 16040
rect 2872 15988 2924 16040
rect 4252 16065 4261 16099
rect 4261 16065 4295 16099
rect 4295 16065 4304 16099
rect 4252 16056 4304 16065
rect 3332 15852 3384 15904
rect 3608 15852 3660 15904
rect 4988 15988 5040 16040
rect 5172 15988 5224 16040
rect 6000 15988 6052 16040
rect 6644 16056 6696 16108
rect 8760 16056 8812 16108
rect 10140 16056 10192 16108
rect 10968 16099 11020 16108
rect 10968 16065 10977 16099
rect 10977 16065 11011 16099
rect 11011 16065 11020 16099
rect 10968 16056 11020 16065
rect 11060 16056 11112 16108
rect 13820 16167 13872 16176
rect 13820 16133 13829 16167
rect 13829 16133 13863 16167
rect 13863 16133 13872 16167
rect 13820 16124 13872 16133
rect 14464 16124 14516 16176
rect 16396 16192 16448 16244
rect 20076 16192 20128 16244
rect 21088 16192 21140 16244
rect 12808 16056 12860 16108
rect 7104 15988 7156 16040
rect 8668 15988 8720 16040
rect 8852 15988 8904 16040
rect 9956 15988 10008 16040
rect 10600 15988 10652 16040
rect 14280 15988 14332 16040
rect 17316 16056 17368 16108
rect 18972 16056 19024 16108
rect 19984 16099 20036 16108
rect 19984 16065 19993 16099
rect 19993 16065 20027 16099
rect 20027 16065 20036 16099
rect 19984 16056 20036 16065
rect 20812 16056 20864 16108
rect 18512 16031 18564 16040
rect 13268 15920 13320 15972
rect 15108 15920 15160 15972
rect 16580 15920 16632 15972
rect 10968 15852 11020 15904
rect 15016 15852 15068 15904
rect 15292 15895 15344 15904
rect 15292 15861 15301 15895
rect 15301 15861 15335 15895
rect 15335 15861 15344 15895
rect 15292 15852 15344 15861
rect 18512 15997 18521 16031
rect 18521 15997 18555 16031
rect 18555 15997 18564 16031
rect 18512 15988 18564 15997
rect 18696 15988 18748 16040
rect 21640 16124 21692 16176
rect 22468 16124 22520 16176
rect 23112 16167 23164 16176
rect 23112 16133 23121 16167
rect 23121 16133 23155 16167
rect 23155 16133 23164 16167
rect 23112 16124 23164 16133
rect 26148 16192 26200 16244
rect 28448 16124 28500 16176
rect 28540 16124 28592 16176
rect 27620 16056 27672 16108
rect 28724 16099 28776 16108
rect 28724 16065 28733 16099
rect 28733 16065 28767 16099
rect 28767 16065 28776 16099
rect 28724 16056 28776 16065
rect 37280 16056 37332 16108
rect 38292 16099 38344 16108
rect 38292 16065 38301 16099
rect 38301 16065 38335 16099
rect 38335 16065 38344 16099
rect 38292 16056 38344 16065
rect 22284 15920 22336 15972
rect 30380 15988 30432 16040
rect 26240 15920 26292 15972
rect 38016 15988 38068 16040
rect 20168 15852 20220 15904
rect 29736 15852 29788 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 3608 15648 3660 15700
rect 9128 15691 9180 15700
rect 3516 15580 3568 15632
rect 1584 15487 1636 15496
rect 1584 15453 1593 15487
rect 1593 15453 1627 15487
rect 1627 15453 1636 15487
rect 1584 15444 1636 15453
rect 3792 15512 3844 15564
rect 4068 15512 4120 15564
rect 5632 15580 5684 15632
rect 6736 15580 6788 15632
rect 4804 15512 4856 15564
rect 3976 15444 4028 15496
rect 6276 15512 6328 15564
rect 9128 15657 9137 15691
rect 9137 15657 9171 15691
rect 9171 15657 9180 15691
rect 9128 15648 9180 15657
rect 8852 15580 8904 15632
rect 10416 15580 10468 15632
rect 12532 15648 12584 15700
rect 12992 15691 13044 15700
rect 12992 15657 13001 15691
rect 13001 15657 13035 15691
rect 13035 15657 13044 15691
rect 12992 15648 13044 15657
rect 7104 15512 7156 15564
rect 10140 15512 10192 15564
rect 12440 15580 12492 15632
rect 19156 15648 19208 15700
rect 20444 15648 20496 15700
rect 21640 15648 21692 15700
rect 12072 15512 12124 15564
rect 12348 15555 12400 15564
rect 12348 15521 12357 15555
rect 12357 15521 12391 15555
rect 12391 15521 12400 15555
rect 12348 15512 12400 15521
rect 12808 15512 12860 15564
rect 6736 15487 6788 15496
rect 6736 15453 6745 15487
rect 6745 15453 6779 15487
rect 6779 15453 6788 15487
rect 6736 15444 6788 15453
rect 9312 15487 9364 15496
rect 9312 15453 9321 15487
rect 9321 15453 9355 15487
rect 9355 15453 9364 15487
rect 9312 15444 9364 15453
rect 9864 15444 9916 15496
rect 10600 15487 10652 15496
rect 10600 15453 10609 15487
rect 10609 15453 10643 15487
rect 10643 15453 10652 15487
rect 10600 15444 10652 15453
rect 13268 15444 13320 15496
rect 2136 15376 2188 15428
rect 7472 15376 7524 15428
rect 12624 15376 12676 15428
rect 7196 15308 7248 15360
rect 9956 15308 10008 15360
rect 10876 15308 10928 15360
rect 15476 15580 15528 15632
rect 16304 15580 16356 15632
rect 19248 15580 19300 15632
rect 20076 15580 20128 15632
rect 16396 15512 16448 15564
rect 16580 15512 16632 15564
rect 18972 15512 19024 15564
rect 19064 15512 19116 15564
rect 20628 15512 20680 15564
rect 24860 15512 24912 15564
rect 28540 15512 28592 15564
rect 14556 15444 14608 15496
rect 17316 15444 17368 15496
rect 18052 15444 18104 15496
rect 12992 15308 13044 15360
rect 14464 15308 14516 15360
rect 14740 15308 14792 15360
rect 15292 15419 15344 15428
rect 15292 15385 15301 15419
rect 15301 15385 15335 15419
rect 15335 15385 15344 15419
rect 15292 15376 15344 15385
rect 16672 15376 16724 15428
rect 16948 15376 17000 15428
rect 18236 15419 18288 15428
rect 18236 15385 18245 15419
rect 18245 15385 18279 15419
rect 18279 15385 18288 15419
rect 18236 15376 18288 15385
rect 18144 15308 18196 15360
rect 18972 15376 19024 15428
rect 19892 15444 19944 15496
rect 20260 15444 20312 15496
rect 21180 15444 21232 15496
rect 27068 15444 27120 15496
rect 29736 15487 29788 15496
rect 29736 15453 29745 15487
rect 29745 15453 29779 15487
rect 29779 15453 29788 15487
rect 29736 15444 29788 15453
rect 23388 15308 23440 15360
rect 27988 15308 28040 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 2688 15104 2740 15156
rect 3332 15147 3384 15156
rect 3332 15113 3341 15147
rect 3341 15113 3375 15147
rect 3375 15113 3384 15147
rect 3332 15104 3384 15113
rect 5540 15147 5592 15156
rect 5540 15113 5549 15147
rect 5549 15113 5583 15147
rect 5583 15113 5592 15147
rect 5540 15104 5592 15113
rect 6092 15104 6144 15156
rect 9036 15104 9088 15156
rect 9496 15104 9548 15156
rect 4068 15079 4120 15088
rect 4068 15045 4077 15079
rect 4077 15045 4111 15079
rect 4111 15045 4120 15079
rect 4068 15036 4120 15045
rect 9404 15036 9456 15088
rect 11888 15036 11940 15088
rect 12532 15036 12584 15088
rect 15292 15104 15344 15156
rect 18880 15104 18932 15156
rect 19156 15104 19208 15156
rect 19340 15147 19392 15156
rect 19340 15113 19349 15147
rect 19349 15113 19383 15147
rect 19383 15113 19392 15147
rect 19340 15104 19392 15113
rect 6184 14968 6236 15020
rect 8208 14968 8260 15020
rect 12072 14968 12124 15020
rect 13544 14968 13596 15020
rect 13728 14968 13780 15020
rect 15844 14968 15896 15020
rect 1584 14943 1636 14952
rect 1584 14909 1593 14943
rect 1593 14909 1627 14943
rect 1627 14909 1636 14943
rect 1584 14900 1636 14909
rect 1860 14943 1912 14952
rect 1216 14832 1268 14884
rect 1860 14909 1869 14943
rect 1869 14909 1903 14943
rect 1903 14909 1912 14943
rect 1860 14900 1912 14909
rect 3792 14943 3844 14952
rect 3792 14909 3801 14943
rect 3801 14909 3835 14943
rect 3835 14909 3844 14943
rect 3792 14900 3844 14909
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 7656 14900 7708 14952
rect 9036 14943 9088 14952
rect 9036 14909 9045 14943
rect 9045 14909 9079 14943
rect 9079 14909 9088 14943
rect 9036 14900 9088 14909
rect 9404 14900 9456 14952
rect 8484 14832 8536 14884
rect 10508 14900 10560 14952
rect 14188 14832 14240 14884
rect 14372 14832 14424 14884
rect 15108 14832 15160 14884
rect 17592 14900 17644 14952
rect 18052 14968 18104 15020
rect 18880 14968 18932 15020
rect 19340 14968 19392 15020
rect 17868 14943 17920 14952
rect 17868 14909 17877 14943
rect 17877 14909 17911 14943
rect 17911 14909 17920 14943
rect 18604 14943 18656 14952
rect 17868 14900 17920 14909
rect 18604 14909 18613 14943
rect 18613 14909 18647 14943
rect 18647 14909 18656 14943
rect 18604 14900 18656 14909
rect 18696 14900 18748 14952
rect 20444 14968 20496 15020
rect 21272 14968 21324 15020
rect 27988 15011 28040 15020
rect 27988 14977 27997 15011
rect 27997 14977 28031 15011
rect 28031 14977 28040 15011
rect 27988 14968 28040 14977
rect 25964 14900 26016 14952
rect 18420 14832 18472 14884
rect 9404 14764 9456 14816
rect 10692 14764 10744 14816
rect 11796 14764 11848 14816
rect 12072 14764 12124 14816
rect 12532 14764 12584 14816
rect 13176 14764 13228 14816
rect 13728 14764 13780 14816
rect 14464 14764 14516 14816
rect 17776 14764 17828 14816
rect 18788 14764 18840 14816
rect 19616 14764 19668 14816
rect 22100 14764 22152 14816
rect 26148 14764 26200 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 3424 14560 3476 14612
rect 4804 14560 4856 14612
rect 5172 14560 5224 14612
rect 5540 14603 5592 14612
rect 5540 14569 5549 14603
rect 5549 14569 5583 14603
rect 5583 14569 5592 14603
rect 5540 14560 5592 14569
rect 6184 14603 6236 14612
rect 6184 14569 6193 14603
rect 6193 14569 6227 14603
rect 6227 14569 6236 14603
rect 6184 14560 6236 14569
rect 12348 14560 12400 14612
rect 13084 14560 13136 14612
rect 14924 14560 14976 14612
rect 16028 14603 16080 14612
rect 16028 14569 16037 14603
rect 16037 14569 16071 14603
rect 16071 14569 16080 14603
rect 16028 14560 16080 14569
rect 17868 14560 17920 14612
rect 26056 14560 26108 14612
rect 4620 14492 4672 14544
rect 11428 14535 11480 14544
rect 1584 14467 1636 14476
rect 1584 14433 1593 14467
rect 1593 14433 1627 14467
rect 1627 14433 1636 14467
rect 1584 14424 1636 14433
rect 2872 14424 2924 14476
rect 3792 14424 3844 14476
rect 4068 14356 4120 14408
rect 5080 14356 5132 14408
rect 5172 14356 5224 14408
rect 11428 14501 11437 14535
rect 11437 14501 11471 14535
rect 11471 14501 11480 14535
rect 11428 14492 11480 14501
rect 6644 14424 6696 14476
rect 7104 14424 7156 14476
rect 9036 14424 9088 14476
rect 10600 14424 10652 14476
rect 12164 14492 12216 14544
rect 1952 14288 2004 14340
rect 3516 14288 3568 14340
rect 5264 14220 5316 14272
rect 11336 14399 11388 14408
rect 11336 14365 11345 14399
rect 11345 14365 11379 14399
rect 11379 14365 11388 14399
rect 11336 14356 11388 14365
rect 11980 14399 12032 14408
rect 11980 14365 11989 14399
rect 11989 14365 12023 14399
rect 12023 14365 12032 14399
rect 13268 14492 13320 14544
rect 12532 14424 12584 14476
rect 18696 14492 18748 14544
rect 21364 14492 21416 14544
rect 25964 14467 26016 14476
rect 25964 14433 25973 14467
rect 25973 14433 26007 14467
rect 26007 14433 26016 14467
rect 25964 14424 26016 14433
rect 26148 14467 26200 14476
rect 26148 14433 26157 14467
rect 26157 14433 26191 14467
rect 26191 14433 26200 14467
rect 26148 14424 26200 14433
rect 37280 14424 37332 14476
rect 11980 14356 12032 14365
rect 12348 14356 12400 14408
rect 7288 14288 7340 14340
rect 7472 14288 7524 14340
rect 8300 14288 8352 14340
rect 7656 14220 7708 14272
rect 13084 14288 13136 14340
rect 11612 14220 11664 14272
rect 13636 14263 13688 14272
rect 13636 14229 13645 14263
rect 13645 14229 13679 14263
rect 13679 14229 13688 14263
rect 13636 14220 13688 14229
rect 19616 14399 19668 14408
rect 14556 14288 14608 14340
rect 15016 14288 15068 14340
rect 19616 14365 19625 14399
rect 19625 14365 19659 14399
rect 19659 14365 19668 14399
rect 19616 14356 19668 14365
rect 21272 14399 21324 14408
rect 21272 14365 21281 14399
rect 21281 14365 21315 14399
rect 21315 14365 21324 14399
rect 21272 14356 21324 14365
rect 22100 14399 22152 14408
rect 22100 14365 22109 14399
rect 22109 14365 22143 14399
rect 22143 14365 22152 14399
rect 22100 14356 22152 14365
rect 22284 14356 22336 14408
rect 27068 14399 27120 14408
rect 17776 14331 17828 14340
rect 17776 14297 17785 14331
rect 17785 14297 17819 14331
rect 17819 14297 17828 14331
rect 17776 14288 17828 14297
rect 18144 14288 18196 14340
rect 18972 14288 19024 14340
rect 21640 14288 21692 14340
rect 27068 14365 27077 14399
rect 27077 14365 27111 14399
rect 27111 14365 27120 14399
rect 27068 14356 27120 14365
rect 37924 14356 37976 14408
rect 16672 14220 16724 14272
rect 18052 14220 18104 14272
rect 20444 14220 20496 14272
rect 20720 14220 20772 14272
rect 38200 14263 38252 14272
rect 38200 14229 38209 14263
rect 38209 14229 38243 14263
rect 38243 14229 38252 14263
rect 38200 14220 38252 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 2780 14016 2832 14068
rect 4620 14059 4672 14068
rect 2228 13991 2280 14000
rect 2228 13957 2237 13991
rect 2237 13957 2271 13991
rect 2271 13957 2280 13991
rect 2228 13948 2280 13957
rect 2320 13948 2372 14000
rect 4620 14025 4629 14059
rect 4629 14025 4663 14059
rect 4663 14025 4672 14059
rect 4620 14016 4672 14025
rect 5816 14059 5868 14068
rect 5816 14025 5825 14059
rect 5825 14025 5859 14059
rect 5859 14025 5868 14059
rect 5816 14016 5868 14025
rect 7012 14016 7064 14068
rect 7380 14059 7432 14068
rect 7380 14025 7389 14059
rect 7389 14025 7423 14059
rect 7423 14025 7432 14059
rect 7380 14016 7432 14025
rect 4712 13948 4764 14000
rect 8852 13991 8904 14000
rect 8852 13957 8861 13991
rect 8861 13957 8895 13991
rect 8895 13957 8904 13991
rect 8852 13948 8904 13957
rect 10324 14059 10376 14068
rect 10324 14025 10333 14059
rect 10333 14025 10367 14059
rect 10367 14025 10376 14059
rect 10324 14016 10376 14025
rect 11520 14016 11572 14068
rect 13912 14016 13964 14068
rect 16948 14016 17000 14068
rect 2872 13923 2924 13932
rect 2872 13889 2881 13923
rect 2881 13889 2915 13923
rect 2915 13889 2924 13923
rect 2872 13880 2924 13889
rect 5080 13923 5132 13932
rect 5080 13889 5089 13923
rect 5089 13889 5123 13923
rect 5123 13889 5132 13923
rect 5080 13880 5132 13889
rect 5908 13812 5960 13864
rect 6092 13880 6144 13932
rect 6736 13880 6788 13932
rect 7656 13880 7708 13932
rect 9956 13880 10008 13932
rect 6828 13812 6880 13864
rect 8852 13812 8904 13864
rect 13636 13948 13688 14000
rect 14740 13991 14792 14000
rect 14740 13957 14749 13991
rect 14749 13957 14783 13991
rect 14783 13957 14792 13991
rect 14740 13948 14792 13957
rect 15108 13948 15160 14000
rect 10692 13880 10744 13932
rect 11704 13880 11756 13932
rect 16856 13948 16908 14000
rect 7748 13744 7800 13796
rect 8024 13744 8076 13796
rect 12716 13812 12768 13864
rect 13452 13812 13504 13864
rect 14372 13812 14424 13864
rect 15200 13812 15252 13864
rect 15936 13812 15988 13864
rect 16672 13880 16724 13932
rect 18604 14016 18656 14068
rect 17684 13991 17736 14000
rect 17684 13957 17693 13991
rect 17693 13957 17727 13991
rect 17727 13957 17736 13991
rect 17684 13948 17736 13957
rect 18880 13880 18932 13932
rect 18972 13880 19024 13932
rect 19156 13880 19208 13932
rect 20628 14016 20680 14068
rect 20444 13991 20496 14000
rect 20444 13957 20453 13991
rect 20453 13957 20487 13991
rect 20487 13957 20496 13991
rect 20444 13948 20496 13957
rect 20904 13948 20956 14000
rect 21456 13991 21508 14000
rect 21456 13957 21465 13991
rect 21465 13957 21499 13991
rect 21499 13957 21508 13991
rect 21456 13948 21508 13957
rect 8576 13676 8628 13728
rect 11980 13744 12032 13796
rect 10232 13676 10284 13728
rect 16120 13744 16172 13796
rect 16212 13787 16264 13796
rect 16212 13753 16221 13787
rect 16221 13753 16255 13787
rect 16255 13753 16264 13787
rect 17776 13812 17828 13864
rect 21272 13812 21324 13864
rect 16212 13744 16264 13753
rect 18236 13744 18288 13796
rect 18696 13744 18748 13796
rect 13636 13676 13688 13728
rect 14648 13676 14700 13728
rect 16028 13676 16080 13728
rect 20628 13676 20680 13728
rect 20996 13676 21048 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 1308 13472 1360 13524
rect 3700 13472 3752 13524
rect 6368 13472 6420 13524
rect 7932 13472 7984 13524
rect 3976 13404 4028 13456
rect 3516 13336 3568 13388
rect 6276 13404 6328 13456
rect 11244 13447 11296 13456
rect 11244 13413 11253 13447
rect 11253 13413 11287 13447
rect 11287 13413 11296 13447
rect 11244 13404 11296 13413
rect 9772 13336 9824 13388
rect 11980 13472 12032 13524
rect 12348 13336 12400 13388
rect 1584 13311 1636 13320
rect 1584 13277 1593 13311
rect 1593 13277 1627 13311
rect 1627 13277 1636 13311
rect 1584 13268 1636 13277
rect 3792 13268 3844 13320
rect 6368 13311 6420 13320
rect 6368 13277 6377 13311
rect 6377 13277 6411 13311
rect 6411 13277 6420 13311
rect 6368 13268 6420 13277
rect 11244 13268 11296 13320
rect 16488 13472 16540 13524
rect 13268 13404 13320 13456
rect 14556 13336 14608 13388
rect 3976 13200 4028 13252
rect 4344 13243 4396 13252
rect 4344 13209 4353 13243
rect 4353 13209 4387 13243
rect 4387 13209 4396 13243
rect 4344 13200 4396 13209
rect 4804 13200 4856 13252
rect 6920 13200 6972 13252
rect 7104 13200 7156 13252
rect 940 13132 992 13184
rect 5632 13132 5684 13184
rect 6460 13132 6512 13184
rect 13544 13200 13596 13252
rect 13636 13200 13688 13252
rect 15476 13268 15528 13320
rect 16764 13268 16816 13320
rect 14372 13243 14424 13252
rect 14372 13209 14381 13243
rect 14381 13209 14415 13243
rect 14415 13209 14424 13243
rect 14372 13200 14424 13209
rect 14464 13243 14516 13252
rect 14464 13209 14473 13243
rect 14473 13209 14507 13243
rect 14507 13209 14516 13243
rect 14464 13200 14516 13209
rect 14832 13200 14884 13252
rect 16948 13268 17000 13320
rect 17316 13268 17368 13320
rect 20260 13404 20312 13456
rect 20628 13472 20680 13524
rect 22284 13472 22336 13524
rect 18788 13336 18840 13388
rect 19892 13336 19944 13388
rect 18696 13311 18748 13320
rect 18696 13277 18705 13311
rect 18705 13277 18739 13311
rect 18739 13277 18748 13311
rect 18696 13268 18748 13277
rect 22100 13311 22152 13320
rect 22100 13277 22109 13311
rect 22109 13277 22143 13311
rect 22143 13277 22152 13311
rect 37648 13472 37700 13524
rect 26424 13447 26476 13456
rect 26424 13413 26433 13447
rect 26433 13413 26467 13447
rect 26467 13413 26476 13447
rect 26424 13404 26476 13413
rect 26056 13379 26108 13388
rect 26056 13345 26065 13379
rect 26065 13345 26099 13379
rect 26099 13345 26108 13379
rect 26056 13336 26108 13345
rect 22100 13268 22152 13277
rect 27528 13268 27580 13320
rect 30380 13268 30432 13320
rect 37280 13268 37332 13320
rect 11060 13132 11112 13184
rect 19156 13200 19208 13252
rect 19524 13243 19576 13252
rect 19524 13209 19533 13243
rect 19533 13209 19567 13243
rect 19567 13209 19576 13243
rect 19524 13200 19576 13209
rect 16672 13132 16724 13184
rect 17960 13132 18012 13184
rect 18788 13132 18840 13184
rect 20444 13200 20496 13252
rect 20996 13200 21048 13252
rect 21272 13132 21324 13184
rect 27712 13132 27764 13184
rect 36912 13132 36964 13184
rect 38200 13175 38252 13184
rect 38200 13141 38209 13175
rect 38209 13141 38243 13175
rect 38243 13141 38252 13175
rect 38200 13132 38252 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 664 12928 716 12980
rect 4804 12928 4856 12980
rect 5908 12928 5960 12980
rect 2872 12860 2924 12912
rect 3424 12860 3476 12912
rect 6368 12860 6420 12912
rect 1584 12767 1636 12776
rect 1584 12733 1593 12767
rect 1593 12733 1627 12767
rect 1627 12733 1636 12767
rect 1584 12724 1636 12733
rect 3516 12724 3568 12776
rect 3240 12656 3292 12708
rect 5632 12792 5684 12844
rect 9772 12860 9824 12912
rect 12440 12928 12492 12980
rect 13084 12860 13136 12912
rect 9680 12792 9732 12844
rect 11060 12792 11112 12844
rect 11336 12792 11388 12844
rect 12624 12835 12676 12844
rect 12624 12801 12633 12835
rect 12633 12801 12667 12835
rect 12667 12801 12676 12835
rect 12624 12792 12676 12801
rect 12992 12792 13044 12844
rect 13452 12860 13504 12912
rect 15476 12860 15528 12912
rect 15660 12903 15712 12912
rect 15660 12869 15669 12903
rect 15669 12869 15703 12903
rect 15703 12869 15712 12903
rect 15660 12860 15712 12869
rect 17132 12860 17184 12912
rect 17316 12903 17368 12912
rect 17316 12869 17325 12903
rect 17325 12869 17359 12903
rect 17359 12869 17368 12903
rect 17316 12860 17368 12869
rect 3700 12724 3752 12776
rect 4252 12724 4304 12776
rect 5632 12699 5684 12708
rect 5632 12665 5641 12699
rect 5641 12665 5675 12699
rect 5675 12665 5684 12699
rect 5632 12656 5684 12665
rect 4620 12588 4672 12640
rect 5172 12588 5224 12640
rect 10324 12724 10376 12776
rect 10416 12724 10468 12776
rect 11980 12724 12032 12776
rect 14832 12792 14884 12844
rect 15292 12792 15344 12844
rect 16948 12835 17000 12844
rect 16948 12801 16957 12835
rect 16957 12801 16991 12835
rect 16991 12801 17000 12835
rect 16948 12792 17000 12801
rect 13636 12724 13688 12776
rect 16120 12724 16172 12776
rect 17316 12724 17368 12776
rect 10232 12588 10284 12640
rect 10324 12588 10376 12640
rect 11888 12656 11940 12708
rect 11796 12631 11848 12640
rect 11796 12597 11805 12631
rect 11805 12597 11839 12631
rect 11839 12597 11848 12631
rect 11796 12588 11848 12597
rect 11980 12588 12032 12640
rect 12624 12588 12676 12640
rect 13268 12588 13320 12640
rect 16212 12656 16264 12708
rect 20076 12928 20128 12980
rect 20904 12971 20956 12980
rect 17592 12860 17644 12912
rect 17776 12860 17828 12912
rect 18420 12860 18472 12912
rect 20904 12937 20913 12971
rect 20913 12937 20947 12971
rect 20947 12937 20956 12971
rect 20904 12928 20956 12937
rect 27528 12971 27580 12980
rect 27528 12937 27537 12971
rect 27537 12937 27571 12971
rect 27571 12937 27580 12971
rect 27528 12928 27580 12937
rect 22100 12860 22152 12912
rect 22836 12860 22888 12912
rect 18420 12767 18472 12776
rect 18420 12733 18429 12767
rect 18429 12733 18463 12767
rect 18463 12733 18472 12767
rect 18420 12724 18472 12733
rect 19524 12724 19576 12776
rect 20444 12724 20496 12776
rect 19892 12656 19944 12708
rect 20076 12656 20128 12708
rect 23572 12792 23624 12844
rect 28356 12835 28408 12844
rect 15936 12588 15988 12640
rect 18420 12588 18472 12640
rect 18604 12588 18656 12640
rect 22652 12656 22704 12708
rect 28356 12801 28365 12835
rect 28365 12801 28399 12835
rect 28399 12801 28408 12835
rect 28356 12792 28408 12801
rect 38108 12835 38160 12844
rect 38108 12801 38117 12835
rect 38117 12801 38151 12835
rect 38151 12801 38160 12835
rect 38108 12792 38160 12801
rect 38200 12631 38252 12640
rect 38200 12597 38209 12631
rect 38209 12597 38243 12631
rect 38243 12597 38252 12631
rect 38200 12588 38252 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 1032 12384 1084 12436
rect 3516 12384 3568 12436
rect 3240 12316 3292 12368
rect 3700 12384 3752 12436
rect 5172 12384 5224 12436
rect 7748 12384 7800 12436
rect 8944 12384 8996 12436
rect 9312 12384 9364 12436
rect 3976 12316 4028 12368
rect 7564 12316 7616 12368
rect 13544 12384 13596 12436
rect 16212 12384 16264 12436
rect 16580 12384 16632 12436
rect 16856 12384 16908 12436
rect 18604 12384 18656 12436
rect 19432 12384 19484 12436
rect 20444 12384 20496 12436
rect 15660 12316 15712 12368
rect 1400 12248 1452 12300
rect 3792 12248 3844 12300
rect 1584 12223 1636 12232
rect 1584 12189 1593 12223
rect 1593 12189 1627 12223
rect 1627 12189 1636 12223
rect 1584 12180 1636 12189
rect 4620 12180 4672 12232
rect 6276 12248 6328 12300
rect 11612 12248 11664 12300
rect 11704 12248 11756 12300
rect 12992 12248 13044 12300
rect 13452 12248 13504 12300
rect 14556 12248 14608 12300
rect 17040 12248 17092 12300
rect 19524 12291 19576 12300
rect 19524 12257 19533 12291
rect 19533 12257 19567 12291
rect 19567 12257 19576 12291
rect 19524 12248 19576 12257
rect 7840 12223 7892 12232
rect 7840 12189 7849 12223
rect 7849 12189 7883 12223
rect 7883 12189 7892 12223
rect 7840 12180 7892 12189
rect 8208 12180 8260 12232
rect 8668 12180 8720 12232
rect 9036 12180 9088 12232
rect 9680 12180 9732 12232
rect 19432 12223 19484 12232
rect 19432 12189 19441 12223
rect 19441 12189 19475 12223
rect 19475 12189 19484 12223
rect 19432 12180 19484 12189
rect 3148 12112 3200 12164
rect 4068 12112 4120 12164
rect 2780 12044 2832 12096
rect 3240 12044 3292 12096
rect 4160 12044 4212 12096
rect 4988 12044 5040 12096
rect 7748 12112 7800 12164
rect 9496 12112 9548 12164
rect 7932 12044 7984 12096
rect 9864 12044 9916 12096
rect 11796 12112 11848 12164
rect 12532 12112 12584 12164
rect 14556 12155 14608 12164
rect 14556 12121 14565 12155
rect 14565 12121 14599 12155
rect 14599 12121 14608 12155
rect 14556 12112 14608 12121
rect 16580 12112 16632 12164
rect 17224 12155 17276 12164
rect 10968 12044 11020 12096
rect 11520 12044 11572 12096
rect 13084 12044 13136 12096
rect 13268 12044 13320 12096
rect 15568 12044 15620 12096
rect 16120 12044 16172 12096
rect 17224 12121 17233 12155
rect 17233 12121 17267 12155
rect 17267 12121 17276 12155
rect 17224 12112 17276 12121
rect 17868 12155 17920 12164
rect 17868 12121 17877 12155
rect 17877 12121 17911 12155
rect 17911 12121 17920 12155
rect 18420 12155 18472 12164
rect 17868 12112 17920 12121
rect 18420 12121 18429 12155
rect 18429 12121 18463 12155
rect 18463 12121 18472 12155
rect 18420 12112 18472 12121
rect 18604 12112 18656 12164
rect 24492 12248 24544 12300
rect 22008 12180 22060 12232
rect 28356 12180 28408 12232
rect 19892 12112 19944 12164
rect 20628 12155 20680 12164
rect 20628 12121 20637 12155
rect 20637 12121 20671 12155
rect 20671 12121 20680 12155
rect 20628 12112 20680 12121
rect 22560 12112 22612 12164
rect 16764 12044 16816 12096
rect 21272 12044 21324 12096
rect 21824 12044 21876 12096
rect 26240 12044 26292 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 1584 11704 1636 11756
rect 3792 11840 3844 11892
rect 4804 11840 4856 11892
rect 7012 11840 7064 11892
rect 4620 11772 4672 11824
rect 6828 11772 6880 11824
rect 9956 11840 10008 11892
rect 9220 11772 9272 11824
rect 6460 11704 6512 11756
rect 6644 11704 6696 11756
rect 9680 11772 9732 11824
rect 10140 11772 10192 11824
rect 4160 11636 4212 11688
rect 5540 11636 5592 11688
rect 5816 11636 5868 11688
rect 6092 11636 6144 11688
rect 7104 11636 7156 11688
rect 12440 11840 12492 11892
rect 11612 11772 11664 11824
rect 11796 11704 11848 11756
rect 12164 11704 12216 11756
rect 13268 11840 13320 11892
rect 14832 11772 14884 11824
rect 12992 11747 13044 11756
rect 12992 11713 13001 11747
rect 13001 11713 13035 11747
rect 13035 11713 13044 11747
rect 12992 11704 13044 11713
rect 12716 11636 12768 11688
rect 15660 11772 15712 11824
rect 16028 11772 16080 11824
rect 16304 11815 16356 11824
rect 16304 11781 16313 11815
rect 16313 11781 16347 11815
rect 16347 11781 16356 11815
rect 16304 11772 16356 11781
rect 16580 11840 16632 11892
rect 16764 11772 16816 11824
rect 16948 11772 17000 11824
rect 17592 11815 17644 11824
rect 17592 11781 17601 11815
rect 17601 11781 17635 11815
rect 17635 11781 17644 11815
rect 17592 11772 17644 11781
rect 20444 11840 20496 11892
rect 23020 11840 23072 11892
rect 28724 11840 28776 11892
rect 21272 11772 21324 11824
rect 15660 11679 15712 11688
rect 15660 11645 15669 11679
rect 15669 11645 15703 11679
rect 15703 11645 15712 11679
rect 15660 11636 15712 11645
rect 16580 11636 16632 11688
rect 1860 11500 1912 11552
rect 6092 11500 6144 11552
rect 9404 11568 9456 11620
rect 12164 11568 12216 11620
rect 14648 11568 14700 11620
rect 17040 11636 17092 11688
rect 17868 11636 17920 11688
rect 18604 11636 18656 11688
rect 23572 11747 23624 11756
rect 18696 11568 18748 11620
rect 19248 11636 19300 11688
rect 23572 11713 23581 11747
rect 23581 11713 23615 11747
rect 23615 11713 23624 11747
rect 23572 11704 23624 11713
rect 24124 11704 24176 11756
rect 21180 11636 21232 11688
rect 22284 11636 22336 11688
rect 22376 11679 22428 11688
rect 22376 11645 22385 11679
rect 22385 11645 22419 11679
rect 22419 11645 22428 11679
rect 22376 11636 22428 11645
rect 20628 11568 20680 11620
rect 25964 11568 26016 11620
rect 8944 11543 8996 11552
rect 8944 11509 8953 11543
rect 8953 11509 8987 11543
rect 8987 11509 8996 11543
rect 8944 11500 8996 11509
rect 9496 11500 9548 11552
rect 18236 11500 18288 11552
rect 21272 11500 21324 11552
rect 21732 11500 21784 11552
rect 23204 11500 23256 11552
rect 23664 11543 23716 11552
rect 23664 11509 23673 11543
rect 23673 11509 23707 11543
rect 23707 11509 23716 11543
rect 23664 11500 23716 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 3424 11296 3476 11348
rect 6000 11296 6052 11348
rect 6644 11296 6696 11348
rect 8300 11296 8352 11348
rect 9220 11339 9272 11348
rect 9220 11305 9229 11339
rect 9229 11305 9263 11339
rect 9263 11305 9272 11339
rect 9220 11296 9272 11305
rect 1584 11203 1636 11212
rect 1584 11169 1593 11203
rect 1593 11169 1627 11203
rect 1627 11169 1636 11203
rect 1584 11160 1636 11169
rect 2320 11160 2372 11212
rect 4620 11160 4672 11212
rect 6276 11160 6328 11212
rect 6920 11160 6972 11212
rect 7288 11160 7340 11212
rect 8944 11228 8996 11280
rect 11612 11296 11664 11348
rect 12440 11296 12492 11348
rect 14188 11296 14240 11348
rect 9772 11228 9824 11280
rect 11520 11271 11572 11280
rect 11520 11237 11529 11271
rect 11529 11237 11563 11271
rect 11563 11237 11572 11271
rect 11520 11228 11572 11237
rect 14556 11296 14608 11348
rect 15568 11296 15620 11348
rect 15752 11228 15804 11280
rect 11980 11203 12032 11212
rect 11980 11169 11989 11203
rect 11989 11169 12023 11203
rect 12023 11169 12032 11203
rect 11980 11160 12032 11169
rect 12256 11160 12308 11212
rect 18236 11228 18288 11280
rect 18420 11228 18472 11280
rect 9772 11135 9824 11144
rect 9772 11101 9781 11135
rect 9781 11101 9815 11135
rect 9815 11101 9824 11135
rect 9772 11092 9824 11101
rect 14280 11135 14332 11144
rect 14280 11101 14289 11135
rect 14289 11101 14323 11135
rect 14323 11101 14332 11135
rect 14280 11092 14332 11101
rect 17960 11160 18012 11212
rect 17868 11092 17920 11144
rect 19340 11160 19392 11212
rect 19616 11160 19668 11212
rect 20720 11160 20772 11212
rect 4896 11024 4948 11076
rect 6000 11024 6052 11076
rect 9036 11024 9088 11076
rect 10048 11067 10100 11076
rect 5356 10956 5408 11008
rect 6736 10956 6788 11008
rect 10048 11033 10057 11067
rect 10057 11033 10091 11067
rect 10091 11033 10100 11067
rect 10048 11024 10100 11033
rect 12164 11024 12216 11076
rect 12348 11024 12400 11076
rect 13544 11024 13596 11076
rect 14188 11024 14240 11076
rect 19064 11092 19116 11144
rect 20168 11092 20220 11144
rect 20444 11092 20496 11144
rect 20628 11135 20680 11144
rect 20628 11101 20637 11135
rect 20637 11101 20671 11135
rect 20671 11101 20680 11135
rect 20628 11092 20680 11101
rect 21180 11296 21232 11348
rect 23112 11296 23164 11348
rect 23296 11339 23348 11348
rect 23296 11305 23305 11339
rect 23305 11305 23339 11339
rect 23339 11305 23348 11339
rect 23296 11296 23348 11305
rect 20996 11160 21048 11212
rect 21824 11160 21876 11212
rect 37372 11160 37424 11212
rect 21916 11135 21968 11144
rect 21916 11101 21925 11135
rect 21925 11101 21959 11135
rect 21959 11101 21968 11135
rect 21916 11092 21968 11101
rect 22836 11092 22888 11144
rect 23204 11135 23256 11144
rect 23204 11101 23213 11135
rect 23213 11101 23247 11135
rect 23247 11101 23256 11135
rect 23204 11092 23256 11101
rect 26240 11092 26292 11144
rect 37188 11092 37240 11144
rect 18696 11024 18748 11076
rect 11428 10956 11480 11008
rect 11612 10956 11664 11008
rect 12440 10956 12492 11008
rect 12900 10956 12952 11008
rect 14004 10956 14056 11008
rect 17040 10956 17092 11008
rect 18512 10956 18564 11008
rect 18880 10956 18932 11008
rect 19616 11067 19668 11076
rect 19616 11033 19625 11067
rect 19625 11033 19659 11067
rect 19659 11033 19668 11067
rect 19616 11024 19668 11033
rect 20260 11024 20312 11076
rect 26148 11067 26200 11076
rect 26148 11033 26157 11067
rect 26157 11033 26191 11067
rect 26191 11033 26200 11067
rect 26148 11024 26200 11033
rect 20628 10956 20680 11008
rect 20904 10956 20956 11008
rect 21364 10999 21416 11008
rect 21364 10965 21373 10999
rect 21373 10965 21407 10999
rect 21407 10965 21416 10999
rect 21364 10956 21416 10965
rect 22652 10999 22704 11008
rect 22652 10965 22661 10999
rect 22661 10965 22695 10999
rect 22695 10965 22704 10999
rect 22652 10956 22704 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 1768 10752 1820 10804
rect 2596 10795 2648 10804
rect 2596 10761 2605 10795
rect 2605 10761 2639 10795
rect 2639 10761 2648 10795
rect 2596 10752 2648 10761
rect 3056 10752 3108 10804
rect 5540 10795 5592 10804
rect 5540 10761 5549 10795
rect 5549 10761 5583 10795
rect 5583 10761 5592 10795
rect 5540 10752 5592 10761
rect 3608 10684 3660 10736
rect 5448 10684 5500 10736
rect 2596 10616 2648 10668
rect 3792 10659 3844 10668
rect 3792 10625 3801 10659
rect 3801 10625 3835 10659
rect 3835 10625 3844 10659
rect 3792 10616 3844 10625
rect 9772 10752 9824 10804
rect 12256 10752 12308 10804
rect 12532 10752 12584 10804
rect 6920 10684 6972 10736
rect 7288 10684 7340 10736
rect 9496 10684 9548 10736
rect 9588 10684 9640 10736
rect 10600 10684 10652 10736
rect 11060 10684 11112 10736
rect 12072 10684 12124 10736
rect 12716 10684 12768 10736
rect 8300 10616 8352 10668
rect 11336 10616 11388 10668
rect 11888 10616 11940 10668
rect 3700 10548 3752 10600
rect 5264 10548 5316 10600
rect 10692 10548 10744 10600
rect 5816 10412 5868 10464
rect 8300 10412 8352 10464
rect 9128 10480 9180 10532
rect 12624 10480 12676 10532
rect 11888 10412 11940 10464
rect 13176 10684 13228 10736
rect 15660 10684 15712 10736
rect 14372 10616 14424 10668
rect 13728 10548 13780 10600
rect 15016 10591 15068 10600
rect 15016 10557 15025 10591
rect 15025 10557 15059 10591
rect 15059 10557 15068 10591
rect 15016 10548 15068 10557
rect 16948 10616 17000 10668
rect 17960 10752 18012 10804
rect 21364 10752 21416 10804
rect 18420 10684 18472 10736
rect 20904 10727 20956 10736
rect 20904 10693 20913 10727
rect 20913 10693 20947 10727
rect 20947 10693 20956 10727
rect 20904 10684 20956 10693
rect 21180 10684 21232 10736
rect 23756 10752 23808 10804
rect 22192 10616 22244 10668
rect 23572 10684 23624 10736
rect 24676 10659 24728 10668
rect 24676 10625 24685 10659
rect 24685 10625 24719 10659
rect 24719 10625 24728 10659
rect 24676 10616 24728 10625
rect 15568 10480 15620 10532
rect 18328 10548 18380 10600
rect 19156 10548 19208 10600
rect 20168 10523 20220 10532
rect 13820 10412 13872 10464
rect 20168 10489 20177 10523
rect 20177 10489 20211 10523
rect 20211 10489 20220 10523
rect 20168 10480 20220 10489
rect 20996 10480 21048 10532
rect 21088 10480 21140 10532
rect 21364 10523 21416 10532
rect 21364 10489 21373 10523
rect 21373 10489 21407 10523
rect 21407 10489 21416 10523
rect 21364 10480 21416 10489
rect 21732 10548 21784 10600
rect 22744 10523 22796 10532
rect 16764 10412 16816 10464
rect 17224 10412 17276 10464
rect 19064 10412 19116 10464
rect 22744 10489 22753 10523
rect 22753 10489 22787 10523
rect 22787 10489 22796 10523
rect 22744 10480 22796 10489
rect 23664 10412 23716 10464
rect 26056 10412 26108 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2596 10251 2648 10260
rect 2596 10217 2605 10251
rect 2605 10217 2639 10251
rect 2639 10217 2648 10251
rect 2596 10208 2648 10217
rect 4712 10208 4764 10260
rect 6920 10208 6972 10260
rect 9680 10251 9732 10260
rect 9680 10217 9689 10251
rect 9689 10217 9723 10251
rect 9723 10217 9732 10251
rect 9680 10208 9732 10217
rect 11888 10208 11940 10260
rect 12164 10208 12216 10260
rect 2872 10140 2924 10192
rect 572 10004 624 10056
rect 3148 10004 3200 10056
rect 3700 10004 3752 10056
rect 6092 10140 6144 10192
rect 14372 10208 14424 10260
rect 22652 10208 22704 10260
rect 14188 10140 14240 10192
rect 15568 10140 15620 10192
rect 18972 10140 19024 10192
rect 19156 10140 19208 10192
rect 3976 10047 4028 10056
rect 3976 10013 3985 10047
rect 3985 10013 4019 10047
rect 4019 10013 4028 10047
rect 3976 10004 4028 10013
rect 8576 10072 8628 10124
rect 13820 10072 13872 10124
rect 14280 10115 14332 10124
rect 14280 10081 14289 10115
rect 14289 10081 14323 10115
rect 14323 10081 14332 10115
rect 14280 10072 14332 10081
rect 17592 10072 17644 10124
rect 20076 10072 20128 10124
rect 21456 10140 21508 10192
rect 21548 10140 21600 10192
rect 20628 10072 20680 10124
rect 4528 9936 4580 9988
rect 9864 10004 9916 10056
rect 4160 9868 4212 9920
rect 6184 9868 6236 9920
rect 6644 9936 6696 9988
rect 7196 9936 7248 9988
rect 9680 9936 9732 9988
rect 10784 10004 10836 10056
rect 12900 10047 12952 10056
rect 12900 10013 12909 10047
rect 12909 10013 12943 10047
rect 12943 10013 12952 10047
rect 12900 10004 12952 10013
rect 14004 10004 14056 10056
rect 16672 10004 16724 10056
rect 18052 10004 18104 10056
rect 22284 10047 22336 10056
rect 11152 9979 11204 9988
rect 11152 9945 11161 9979
rect 11161 9945 11195 9979
rect 11195 9945 11204 9979
rect 11152 9936 11204 9945
rect 12624 9936 12676 9988
rect 15292 9936 15344 9988
rect 15844 9936 15896 9988
rect 18420 9936 18472 9988
rect 19248 9936 19300 9988
rect 22284 10013 22293 10047
rect 22293 10013 22327 10047
rect 22327 10013 22336 10047
rect 22284 10004 22336 10013
rect 23204 10004 23256 10056
rect 19524 9936 19576 9988
rect 20352 9936 20404 9988
rect 21088 9979 21140 9988
rect 21088 9945 21097 9979
rect 21097 9945 21131 9979
rect 21131 9945 21140 9979
rect 21088 9936 21140 9945
rect 21732 9936 21784 9988
rect 21916 9936 21968 9988
rect 23020 9936 23072 9988
rect 36912 10004 36964 10056
rect 37740 9936 37792 9988
rect 6920 9868 6972 9920
rect 7472 9868 7524 9920
rect 7656 9868 7708 9920
rect 8116 9868 8168 9920
rect 13728 9868 13780 9920
rect 14372 9868 14424 9920
rect 14464 9868 14516 9920
rect 17224 9868 17276 9920
rect 22008 9868 22060 9920
rect 24952 9868 25004 9920
rect 38200 9911 38252 9920
rect 38200 9877 38209 9911
rect 38209 9877 38243 9911
rect 38243 9877 38252 9911
rect 38200 9868 38252 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 3792 9664 3844 9716
rect 5356 9664 5408 9716
rect 5540 9664 5592 9716
rect 3884 9596 3936 9648
rect 4988 9596 5040 9648
rect 6552 9664 6604 9716
rect 6644 9664 6696 9716
rect 13360 9664 13412 9716
rect 14188 9664 14240 9716
rect 17224 9664 17276 9716
rect 21916 9664 21968 9716
rect 22284 9664 22336 9716
rect 7104 9596 7156 9648
rect 8576 9596 8628 9648
rect 10784 9596 10836 9648
rect 11060 9596 11112 9648
rect 11704 9639 11756 9648
rect 11704 9605 11713 9639
rect 11713 9605 11747 9639
rect 11747 9605 11756 9639
rect 11704 9596 11756 9605
rect 11980 9596 12032 9648
rect 13268 9639 13320 9648
rect 13268 9605 13277 9639
rect 13277 9605 13311 9639
rect 13311 9605 13320 9639
rect 13268 9596 13320 9605
rect 15476 9596 15528 9648
rect 15844 9596 15896 9648
rect 1584 9503 1636 9512
rect 1584 9469 1593 9503
rect 1593 9469 1627 9503
rect 1627 9469 1636 9503
rect 1584 9460 1636 9469
rect 4160 9528 4212 9580
rect 7012 9528 7064 9580
rect 8944 9528 8996 9580
rect 12256 9528 12308 9580
rect 13820 9571 13872 9580
rect 13820 9537 13829 9571
rect 13829 9537 13863 9571
rect 13863 9537 13872 9571
rect 13820 9528 13872 9537
rect 16028 9528 16080 9580
rect 3976 9460 4028 9512
rect 1584 9324 1636 9376
rect 3424 9324 3476 9376
rect 5172 9460 5224 9512
rect 8208 9460 8260 9512
rect 8024 9392 8076 9444
rect 9680 9460 9732 9512
rect 10968 9392 11020 9444
rect 11888 9460 11940 9512
rect 14188 9460 14240 9512
rect 14464 9460 14516 9512
rect 16304 9571 16356 9580
rect 16304 9537 16313 9571
rect 16313 9537 16347 9571
rect 16347 9537 16356 9571
rect 16304 9528 16356 9537
rect 18144 9596 18196 9648
rect 20536 9596 20588 9648
rect 24952 9639 25004 9648
rect 24952 9605 24961 9639
rect 24961 9605 24995 9639
rect 24995 9605 25004 9639
rect 24952 9596 25004 9605
rect 25044 9639 25096 9648
rect 25044 9605 25053 9639
rect 25053 9605 25087 9639
rect 25087 9605 25096 9639
rect 25044 9596 25096 9605
rect 17408 9528 17460 9580
rect 19064 9528 19116 9580
rect 19156 9571 19208 9580
rect 19156 9537 19165 9571
rect 19165 9537 19199 9571
rect 19199 9537 19208 9571
rect 19156 9528 19208 9537
rect 19984 9528 20036 9580
rect 20628 9528 20680 9580
rect 21548 9528 21600 9580
rect 22008 9571 22060 9580
rect 22008 9537 22017 9571
rect 22017 9537 22051 9571
rect 22051 9537 22060 9571
rect 22008 9528 22060 9537
rect 22100 9571 22152 9580
rect 22100 9537 22109 9571
rect 22109 9537 22143 9571
rect 22143 9537 22152 9571
rect 22100 9528 22152 9537
rect 22284 9528 22336 9580
rect 22836 9528 22888 9580
rect 23388 9571 23440 9580
rect 23388 9537 23397 9571
rect 23397 9537 23431 9571
rect 23431 9537 23440 9571
rect 23388 9528 23440 9537
rect 23940 9528 23992 9580
rect 31392 9528 31444 9580
rect 20996 9460 21048 9512
rect 21088 9460 21140 9512
rect 4712 9324 4764 9376
rect 8116 9324 8168 9376
rect 12256 9324 12308 9376
rect 18052 9392 18104 9444
rect 18604 9392 18656 9444
rect 21732 9392 21784 9444
rect 22008 9392 22060 9444
rect 24032 9392 24084 9444
rect 24860 9392 24912 9444
rect 15568 9367 15620 9376
rect 15568 9333 15577 9367
rect 15577 9333 15611 9367
rect 15611 9333 15620 9367
rect 15568 9324 15620 9333
rect 16948 9324 17000 9376
rect 19340 9324 19392 9376
rect 20076 9324 20128 9376
rect 20168 9324 20220 9376
rect 22192 9324 22244 9376
rect 30012 9367 30064 9376
rect 30012 9333 30021 9367
rect 30021 9333 30055 9367
rect 30055 9333 30064 9367
rect 30012 9324 30064 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2044 9163 2096 9172
rect 2044 9129 2053 9163
rect 2053 9129 2087 9163
rect 2087 9129 2096 9163
rect 2044 9120 2096 9129
rect 2504 9120 2556 9172
rect 3332 9163 3384 9172
rect 3332 9129 3341 9163
rect 3341 9129 3375 9163
rect 3375 9129 3384 9163
rect 3332 9120 3384 9129
rect 7748 9120 7800 9172
rect 8944 9120 8996 9172
rect 9864 9120 9916 9172
rect 12256 9120 12308 9172
rect 12624 9163 12676 9172
rect 12624 9129 12633 9163
rect 12633 9129 12667 9163
rect 12667 9129 12676 9163
rect 12624 9120 12676 9129
rect 15292 9120 15344 9172
rect 16028 9120 16080 9172
rect 21548 9120 21600 9172
rect 21732 9120 21784 9172
rect 23480 9163 23532 9172
rect 7472 9052 7524 9104
rect 8392 9052 8444 9104
rect 4712 9027 4764 9036
rect 4712 8993 4721 9027
rect 4721 8993 4755 9027
rect 4755 8993 4764 9027
rect 4712 8984 4764 8993
rect 1952 8959 2004 8968
rect 1952 8925 1961 8959
rect 1961 8925 1995 8959
rect 1995 8925 2004 8959
rect 1952 8916 2004 8925
rect 2780 8959 2832 8968
rect 2780 8925 2789 8959
rect 2789 8925 2823 8959
rect 2823 8925 2832 8959
rect 2780 8916 2832 8925
rect 3516 8916 3568 8968
rect 4068 8916 4120 8968
rect 7012 8984 7064 9036
rect 9772 8984 9824 9036
rect 11888 9052 11940 9104
rect 12532 9052 12584 9104
rect 3700 8848 3752 8900
rect 6644 8916 6696 8968
rect 6920 8916 6972 8968
rect 8208 8916 8260 8968
rect 9864 8916 9916 8968
rect 13728 8984 13780 9036
rect 13820 8984 13872 9036
rect 15844 9052 15896 9104
rect 15568 8984 15620 9036
rect 16856 8984 16908 9036
rect 17224 9052 17276 9104
rect 23480 9129 23489 9163
rect 23489 9129 23523 9163
rect 23523 9129 23532 9163
rect 23480 9120 23532 9129
rect 17408 8984 17460 9036
rect 12348 8916 12400 8968
rect 13912 8916 13964 8968
rect 6736 8848 6788 8900
rect 7012 8848 7064 8900
rect 2780 8780 2832 8832
rect 3240 8780 3292 8832
rect 6092 8780 6144 8832
rect 9680 8848 9732 8900
rect 9956 8848 10008 8900
rect 12164 8848 12216 8900
rect 14464 8848 14516 8900
rect 14832 8848 14884 8900
rect 15844 8848 15896 8900
rect 20536 8916 20588 8968
rect 21640 8959 21692 8968
rect 21640 8925 21649 8959
rect 21649 8925 21683 8959
rect 21683 8925 21692 8959
rect 21640 8916 21692 8925
rect 22100 8959 22152 8968
rect 22100 8925 22109 8959
rect 22109 8925 22143 8959
rect 22143 8925 22152 8959
rect 22744 8959 22796 8968
rect 22100 8916 22152 8925
rect 22744 8925 22753 8959
rect 22753 8925 22787 8959
rect 22787 8925 22796 8959
rect 22744 8916 22796 8925
rect 17684 8848 17736 8900
rect 18144 8891 18196 8900
rect 18144 8857 18153 8891
rect 18153 8857 18187 8891
rect 18187 8857 18196 8891
rect 18144 8848 18196 8857
rect 10324 8780 10376 8832
rect 11060 8780 11112 8832
rect 12440 8780 12492 8832
rect 12532 8780 12584 8832
rect 17868 8780 17920 8832
rect 18512 8848 18564 8900
rect 19156 8848 19208 8900
rect 20996 8891 21048 8900
rect 20996 8857 21005 8891
rect 21005 8857 21039 8891
rect 21039 8857 21048 8891
rect 20996 8848 21048 8857
rect 20904 8780 20956 8832
rect 22836 8823 22888 8832
rect 22836 8789 22845 8823
rect 22845 8789 22879 8823
rect 22879 8789 22888 8823
rect 22836 8780 22888 8789
rect 25044 9052 25096 9104
rect 24584 8959 24636 8968
rect 24584 8925 24593 8959
rect 24593 8925 24627 8959
rect 24627 8925 24636 8959
rect 24584 8916 24636 8925
rect 25228 8848 25280 8900
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 1952 8576 2004 8628
rect 7104 8576 7156 8628
rect 2780 8508 2832 8560
rect 3516 8508 3568 8560
rect 3976 8508 4028 8560
rect 1676 8372 1728 8424
rect 4804 8440 4856 8492
rect 5356 8508 5408 8560
rect 11060 8576 11112 8628
rect 6736 8440 6788 8492
rect 10692 8508 10744 8560
rect 756 8304 808 8356
rect 4712 8372 4764 8424
rect 4896 8372 4948 8424
rect 5448 8304 5500 8356
rect 3976 8279 4028 8288
rect 3976 8245 3985 8279
rect 3985 8245 4019 8279
rect 4019 8245 4028 8279
rect 3976 8236 4028 8245
rect 4712 8236 4764 8288
rect 7840 8304 7892 8356
rect 11980 8508 12032 8560
rect 12624 8576 12676 8628
rect 13636 8576 13688 8628
rect 8208 8372 8260 8424
rect 10140 8372 10192 8424
rect 10232 8372 10284 8424
rect 17224 8576 17276 8628
rect 17408 8576 17460 8628
rect 15568 8508 15620 8560
rect 16304 8508 16356 8560
rect 17592 8551 17644 8560
rect 17592 8517 17601 8551
rect 17601 8517 17635 8551
rect 17635 8517 17644 8551
rect 17592 8508 17644 8517
rect 13820 8440 13872 8492
rect 15476 8440 15528 8492
rect 16396 8372 16448 8424
rect 18144 8576 18196 8628
rect 20444 8576 20496 8628
rect 20996 8576 21048 8628
rect 30012 8576 30064 8628
rect 17868 8508 17920 8560
rect 19340 8508 19392 8560
rect 22836 8508 22888 8560
rect 38384 8508 38436 8560
rect 18052 8483 18104 8492
rect 18052 8449 18061 8483
rect 18061 8449 18095 8483
rect 18095 8449 18104 8483
rect 18052 8440 18104 8449
rect 18696 8440 18748 8492
rect 18972 8440 19024 8492
rect 19340 8415 19392 8424
rect 10140 8236 10192 8288
rect 12532 8236 12584 8288
rect 16120 8304 16172 8356
rect 14280 8236 14332 8288
rect 14924 8236 14976 8288
rect 15200 8236 15252 8288
rect 16028 8236 16080 8288
rect 19340 8381 19349 8415
rect 19349 8381 19383 8415
rect 19383 8381 19392 8415
rect 19340 8372 19392 8381
rect 22376 8440 22428 8492
rect 22652 8483 22704 8492
rect 22652 8449 22661 8483
rect 22661 8449 22695 8483
rect 22695 8449 22704 8483
rect 22652 8440 22704 8449
rect 23296 8483 23348 8492
rect 23296 8449 23305 8483
rect 23305 8449 23339 8483
rect 23339 8449 23348 8483
rect 23296 8440 23348 8449
rect 23388 8440 23440 8492
rect 24032 8440 24084 8492
rect 25228 8483 25280 8492
rect 25228 8449 25237 8483
rect 25237 8449 25271 8483
rect 25271 8449 25280 8483
rect 25228 8440 25280 8449
rect 38108 8483 38160 8492
rect 38108 8449 38117 8483
rect 38117 8449 38151 8483
rect 38151 8449 38160 8483
rect 38108 8440 38160 8449
rect 20812 8372 20864 8424
rect 22008 8415 22060 8424
rect 22008 8381 22017 8415
rect 22017 8381 22051 8415
rect 22051 8381 22060 8415
rect 22008 8372 22060 8381
rect 22744 8415 22796 8424
rect 22744 8381 22753 8415
rect 22753 8381 22787 8415
rect 22787 8381 22796 8415
rect 22744 8372 22796 8381
rect 20628 8304 20680 8356
rect 20720 8304 20772 8356
rect 25320 8347 25372 8356
rect 25320 8313 25329 8347
rect 25329 8313 25363 8347
rect 25363 8313 25372 8347
rect 25320 8304 25372 8313
rect 18236 8236 18288 8288
rect 18696 8236 18748 8288
rect 21088 8236 21140 8288
rect 21180 8236 21232 8288
rect 21916 8236 21968 8288
rect 22836 8236 22888 8288
rect 24676 8279 24728 8288
rect 24676 8245 24685 8279
rect 24685 8245 24719 8279
rect 24719 8245 24728 8279
rect 24676 8236 24728 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 3424 8075 3476 8084
rect 1676 7939 1728 7948
rect 1676 7905 1685 7939
rect 1685 7905 1719 7939
rect 1719 7905 1728 7939
rect 1676 7896 1728 7905
rect 3424 8041 3433 8075
rect 3433 8041 3467 8075
rect 3467 8041 3476 8075
rect 3424 8032 3476 8041
rect 6000 8075 6052 8084
rect 6000 8041 6009 8075
rect 6009 8041 6043 8075
rect 6043 8041 6052 8075
rect 6000 8032 6052 8041
rect 7196 8032 7248 8084
rect 12072 8032 12124 8084
rect 12716 8032 12768 8084
rect 11612 7964 11664 8016
rect 16120 8032 16172 8084
rect 3976 7896 4028 7948
rect 11980 7939 12032 7948
rect 4712 7828 4764 7880
rect 3976 7760 4028 7812
rect 5540 7760 5592 7812
rect 6644 7828 6696 7880
rect 9036 7828 9088 7880
rect 6460 7760 6512 7812
rect 9772 7760 9824 7812
rect 10324 7760 10376 7812
rect 4160 7735 4212 7744
rect 4160 7701 4169 7735
rect 4169 7701 4203 7735
rect 4203 7701 4212 7735
rect 4160 7692 4212 7701
rect 5448 7692 5500 7744
rect 11612 7692 11664 7744
rect 11980 7905 11989 7939
rect 11989 7905 12023 7939
rect 12023 7905 12032 7939
rect 11980 7896 12032 7905
rect 14096 7896 14148 7948
rect 16396 7896 16448 7948
rect 18328 7964 18380 8016
rect 19248 7964 19300 8016
rect 19892 8032 19944 8084
rect 23940 8032 23992 8084
rect 23296 7964 23348 8016
rect 13728 7828 13780 7880
rect 19524 7939 19576 7948
rect 17868 7828 17920 7880
rect 14832 7760 14884 7812
rect 16396 7760 16448 7812
rect 16672 7803 16724 7812
rect 16672 7769 16681 7803
rect 16681 7769 16715 7803
rect 16715 7769 16724 7803
rect 16672 7760 16724 7769
rect 12900 7692 12952 7744
rect 14556 7692 14608 7744
rect 18236 7803 18288 7812
rect 18236 7769 18245 7803
rect 18245 7769 18279 7803
rect 18279 7769 18288 7803
rect 18236 7760 18288 7769
rect 19064 7760 19116 7812
rect 19524 7905 19533 7939
rect 19533 7905 19567 7939
rect 19567 7905 19576 7939
rect 19524 7896 19576 7905
rect 22008 7896 22060 7948
rect 22100 7896 22152 7948
rect 19432 7871 19484 7880
rect 19432 7837 19441 7871
rect 19441 7837 19475 7871
rect 19475 7837 19484 7871
rect 19432 7828 19484 7837
rect 19892 7760 19944 7812
rect 20260 7803 20312 7812
rect 20260 7769 20269 7803
rect 20269 7769 20303 7803
rect 20303 7769 20312 7803
rect 21180 7803 21232 7812
rect 20260 7760 20312 7769
rect 21180 7769 21189 7803
rect 21189 7769 21223 7803
rect 21223 7769 21232 7803
rect 21180 7760 21232 7769
rect 21272 7760 21324 7812
rect 22652 7760 22704 7812
rect 26240 7896 26292 7948
rect 37740 7939 37792 7948
rect 37740 7905 37749 7939
rect 37749 7905 37783 7939
rect 37783 7905 37792 7939
rect 37740 7896 37792 7905
rect 30748 7828 30800 7880
rect 37464 7871 37516 7880
rect 37464 7837 37473 7871
rect 37473 7837 37507 7871
rect 37507 7837 37516 7871
rect 37464 7828 37516 7837
rect 24676 7760 24728 7812
rect 22836 7692 22888 7744
rect 22928 7692 22980 7744
rect 23388 7692 23440 7744
rect 24584 7735 24636 7744
rect 24584 7701 24593 7735
rect 24593 7701 24627 7735
rect 24627 7701 24636 7735
rect 24584 7692 24636 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 5080 7488 5132 7540
rect 1400 7420 1452 7472
rect 1768 7352 1820 7404
rect 4160 7352 4212 7404
rect 6644 7488 6696 7540
rect 9956 7488 10008 7540
rect 9128 7463 9180 7472
rect 9128 7429 9137 7463
rect 9137 7429 9171 7463
rect 9171 7429 9180 7463
rect 9128 7420 9180 7429
rect 10968 7420 11020 7472
rect 17224 7488 17276 7540
rect 11980 7420 12032 7472
rect 13452 7420 13504 7472
rect 13820 7420 13872 7472
rect 20720 7488 20772 7540
rect 21272 7488 21324 7540
rect 25964 7488 26016 7540
rect 17684 7420 17736 7472
rect 18144 7420 18196 7472
rect 18696 7420 18748 7472
rect 18880 7463 18932 7472
rect 18880 7429 18889 7463
rect 18889 7429 18923 7463
rect 18923 7429 18932 7463
rect 18880 7420 18932 7429
rect 23388 7420 23440 7472
rect 3424 7284 3476 7336
rect 6552 7284 6604 7336
rect 8852 7327 8904 7336
rect 8852 7293 8861 7327
rect 8861 7293 8895 7327
rect 8895 7293 8904 7327
rect 8852 7284 8904 7293
rect 1860 7259 1912 7268
rect 1860 7225 1869 7259
rect 1869 7225 1903 7259
rect 1903 7225 1912 7259
rect 1860 7216 1912 7225
rect 8116 7148 8168 7200
rect 8576 7148 8628 7200
rect 12716 7284 12768 7336
rect 12992 7284 13044 7336
rect 13636 7284 13688 7336
rect 13728 7284 13780 7336
rect 14280 7327 14332 7336
rect 14280 7293 14289 7327
rect 14289 7293 14323 7327
rect 14323 7293 14332 7327
rect 14280 7284 14332 7293
rect 15752 7327 15804 7336
rect 15752 7293 15761 7327
rect 15761 7293 15795 7327
rect 15795 7293 15804 7327
rect 15752 7284 15804 7293
rect 17592 7284 17644 7336
rect 20168 7352 20220 7404
rect 20812 7395 20864 7404
rect 20812 7361 20821 7395
rect 20821 7361 20855 7395
rect 20855 7361 20864 7395
rect 20812 7352 20864 7361
rect 15568 7216 15620 7268
rect 17684 7216 17736 7268
rect 19432 7216 19484 7268
rect 21364 7352 21416 7404
rect 22192 7395 22244 7404
rect 22192 7361 22201 7395
rect 22201 7361 22235 7395
rect 22235 7361 22244 7395
rect 22192 7352 22244 7361
rect 16580 7148 16632 7200
rect 18512 7148 18564 7200
rect 19156 7148 19208 7200
rect 20904 7148 20956 7200
rect 22284 7284 22336 7336
rect 24584 7352 24636 7404
rect 27160 7395 27212 7404
rect 22468 7284 22520 7336
rect 27160 7361 27169 7395
rect 27169 7361 27203 7395
rect 27203 7361 27212 7395
rect 27160 7352 27212 7361
rect 30104 7284 30156 7336
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 6828 6944 6880 6996
rect 9680 6944 9732 6996
rect 9772 6944 9824 6996
rect 1768 6919 1820 6928
rect 1768 6885 1777 6919
rect 1777 6885 1811 6919
rect 1811 6885 1820 6919
rect 1768 6876 1820 6885
rect 3884 6808 3936 6860
rect 6552 6808 6604 6860
rect 1584 6783 1636 6792
rect 1584 6749 1593 6783
rect 1593 6749 1627 6783
rect 1627 6749 1636 6783
rect 1584 6740 1636 6749
rect 1952 6740 2004 6792
rect 3240 6740 3292 6792
rect 3608 6740 3660 6792
rect 6736 6808 6788 6860
rect 8944 6808 8996 6860
rect 9036 6808 9088 6860
rect 12716 6944 12768 6996
rect 13820 6944 13872 6996
rect 15936 6944 15988 6996
rect 16396 6944 16448 6996
rect 8208 6740 8260 6792
rect 9220 6783 9272 6792
rect 9220 6749 9229 6783
rect 9229 6749 9263 6783
rect 9263 6749 9272 6783
rect 9220 6740 9272 6749
rect 9312 6783 9364 6792
rect 9312 6749 9321 6783
rect 9321 6749 9355 6783
rect 9355 6749 9364 6783
rect 9312 6740 9364 6749
rect 9680 6740 9732 6792
rect 11152 6851 11204 6860
rect 11152 6817 11161 6851
rect 11161 6817 11195 6851
rect 11195 6817 11204 6851
rect 11152 6808 11204 6817
rect 13268 6876 13320 6928
rect 10508 6783 10560 6792
rect 10508 6749 10517 6783
rect 10517 6749 10551 6783
rect 10551 6749 10560 6783
rect 10508 6740 10560 6749
rect 13176 6740 13228 6792
rect 13544 6808 13596 6860
rect 16488 6876 16540 6928
rect 15568 6808 15620 6860
rect 17776 6851 17828 6860
rect 13728 6740 13780 6792
rect 10876 6672 10928 6724
rect 11428 6715 11480 6724
rect 2228 6604 2280 6656
rect 6828 6604 6880 6656
rect 7656 6647 7708 6656
rect 7656 6613 7665 6647
rect 7665 6613 7699 6647
rect 7699 6613 7708 6647
rect 7656 6604 7708 6613
rect 9680 6604 9732 6656
rect 10416 6604 10468 6656
rect 11060 6604 11112 6656
rect 11428 6681 11437 6715
rect 11437 6681 11471 6715
rect 11471 6681 11480 6715
rect 11428 6672 11480 6681
rect 16580 6715 16632 6724
rect 16580 6681 16589 6715
rect 16589 6681 16623 6715
rect 16623 6681 16632 6715
rect 16580 6672 16632 6681
rect 17776 6817 17785 6851
rect 17785 6817 17819 6851
rect 17819 6817 17828 6851
rect 17776 6808 17828 6817
rect 18236 6876 18288 6928
rect 19064 6876 19116 6928
rect 20904 6876 20956 6928
rect 21732 6876 21784 6928
rect 22284 6876 22336 6928
rect 23388 6876 23440 6928
rect 18512 6808 18564 6860
rect 19340 6808 19392 6860
rect 17408 6740 17460 6792
rect 20444 6740 20496 6792
rect 21548 6808 21600 6860
rect 19432 6604 19484 6656
rect 20904 6672 20956 6724
rect 22100 6740 22152 6792
rect 22652 6740 22704 6792
rect 23112 6740 23164 6792
rect 23296 6783 23348 6792
rect 23296 6749 23305 6783
rect 23305 6749 23339 6783
rect 23339 6749 23348 6783
rect 23296 6740 23348 6749
rect 22376 6672 22428 6724
rect 21272 6604 21324 6656
rect 21456 6604 21508 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 1952 6443 2004 6452
rect 1952 6409 1961 6443
rect 1961 6409 1995 6443
rect 1995 6409 2004 6443
rect 1952 6400 2004 6409
rect 4988 6400 5040 6452
rect 7012 6400 7064 6452
rect 2320 6264 2372 6316
rect 3424 6264 3476 6316
rect 5540 6264 5592 6316
rect 6920 6332 6972 6384
rect 8668 6332 8720 6384
rect 11060 6400 11112 6452
rect 13268 6400 13320 6452
rect 11336 6332 11388 6384
rect 11704 6375 11756 6384
rect 11704 6341 11713 6375
rect 11713 6341 11747 6375
rect 11747 6341 11756 6375
rect 11704 6332 11756 6341
rect 9036 6307 9088 6316
rect 9036 6273 9045 6307
rect 9045 6273 9079 6307
rect 9079 6273 9088 6307
rect 9036 6264 9088 6273
rect 4712 6196 4764 6248
rect 5264 6196 5316 6248
rect 5540 6128 5592 6180
rect 9864 6196 9916 6248
rect 11152 6264 11204 6316
rect 15752 6400 15804 6452
rect 13728 6332 13780 6384
rect 13820 6332 13872 6384
rect 13452 6239 13504 6248
rect 13452 6205 13461 6239
rect 13461 6205 13495 6239
rect 13495 6205 13504 6239
rect 13452 6196 13504 6205
rect 15200 6196 15252 6248
rect 10324 6128 10376 6180
rect 12256 6128 12308 6180
rect 15660 6239 15712 6248
rect 15660 6205 15669 6239
rect 15669 6205 15703 6239
rect 15703 6205 15712 6239
rect 15660 6196 15712 6205
rect 17132 6332 17184 6384
rect 17776 6375 17828 6384
rect 17776 6341 17785 6375
rect 17785 6341 17819 6375
rect 17819 6341 17828 6375
rect 17776 6332 17828 6341
rect 18052 6400 18104 6452
rect 19800 6400 19852 6452
rect 20352 6443 20404 6452
rect 20352 6409 20361 6443
rect 20361 6409 20395 6443
rect 20395 6409 20404 6443
rect 20352 6400 20404 6409
rect 20904 6400 20956 6452
rect 22744 6400 22796 6452
rect 21088 6332 21140 6384
rect 17316 6264 17368 6316
rect 20168 6264 20220 6316
rect 20628 6264 20680 6316
rect 20904 6307 20956 6316
rect 20904 6273 20913 6307
rect 20913 6273 20947 6307
rect 20947 6273 20956 6307
rect 20904 6264 20956 6273
rect 18144 6239 18196 6248
rect 2504 6103 2556 6112
rect 2504 6069 2513 6103
rect 2513 6069 2547 6103
rect 2547 6069 2556 6103
rect 2504 6060 2556 6069
rect 3056 6060 3108 6112
rect 5632 6060 5684 6112
rect 8392 6060 8444 6112
rect 8668 6103 8720 6112
rect 8668 6069 8677 6103
rect 8677 6069 8711 6103
rect 8711 6069 8720 6103
rect 8668 6060 8720 6069
rect 10048 6060 10100 6112
rect 12440 6060 12492 6112
rect 15384 6128 15436 6180
rect 17408 6128 17460 6180
rect 18144 6205 18153 6239
rect 18153 6205 18187 6239
rect 18187 6205 18196 6239
rect 18144 6196 18196 6205
rect 21088 6196 21140 6248
rect 38292 6307 38344 6316
rect 38292 6273 38301 6307
rect 38301 6273 38335 6307
rect 38335 6273 38344 6307
rect 38292 6264 38344 6273
rect 20628 6128 20680 6180
rect 23020 6196 23072 6248
rect 23204 6239 23256 6248
rect 23204 6205 23213 6239
rect 23213 6205 23247 6239
rect 23247 6205 23256 6239
rect 23204 6196 23256 6205
rect 23112 6128 23164 6180
rect 30656 6171 30708 6180
rect 30656 6137 30665 6171
rect 30665 6137 30699 6171
rect 30699 6137 30708 6171
rect 30656 6128 30708 6137
rect 15936 6060 15988 6112
rect 16304 6103 16356 6112
rect 16304 6069 16313 6103
rect 16313 6069 16347 6103
rect 16347 6069 16356 6103
rect 16304 6060 16356 6069
rect 18604 6060 18656 6112
rect 19524 6103 19576 6112
rect 19524 6069 19533 6103
rect 19533 6069 19567 6103
rect 19567 6069 19576 6103
rect 19524 6060 19576 6069
rect 19800 6060 19852 6112
rect 20904 6060 20956 6112
rect 21088 6060 21140 6112
rect 22928 6060 22980 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 1584 5856 1636 5908
rect 6920 5856 6972 5908
rect 7288 5856 7340 5908
rect 10324 5856 10376 5908
rect 12440 5856 12492 5908
rect 16304 5856 16356 5908
rect 19524 5856 19576 5908
rect 19616 5856 19668 5908
rect 4068 5788 4120 5840
rect 5264 5763 5316 5772
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 2872 5584 2924 5636
rect 3792 5584 3844 5636
rect 4896 5516 4948 5568
rect 5264 5729 5273 5763
rect 5273 5729 5307 5763
rect 5307 5729 5316 5763
rect 5264 5720 5316 5729
rect 6552 5720 6604 5772
rect 8484 5720 8536 5772
rect 6828 5652 6880 5704
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 8852 5720 8904 5772
rect 5632 5584 5684 5636
rect 7288 5627 7340 5636
rect 7288 5593 7297 5627
rect 7297 5593 7331 5627
rect 7331 5593 7340 5627
rect 7288 5584 7340 5593
rect 9036 5584 9088 5636
rect 9680 5584 9732 5636
rect 10600 5584 10652 5636
rect 11060 5516 11112 5568
rect 13452 5720 13504 5772
rect 16028 5720 16080 5772
rect 17408 5720 17460 5772
rect 17592 5763 17644 5772
rect 17592 5729 17601 5763
rect 17601 5729 17635 5763
rect 17635 5729 17644 5763
rect 17592 5720 17644 5729
rect 19248 5788 19300 5840
rect 20260 5856 20312 5908
rect 20628 5856 20680 5908
rect 22284 5856 22336 5908
rect 22376 5856 22428 5908
rect 24492 5856 24544 5908
rect 12256 5584 12308 5636
rect 13452 5584 13504 5636
rect 15660 5652 15712 5704
rect 14556 5627 14608 5636
rect 14556 5593 14565 5627
rect 14565 5593 14599 5627
rect 14599 5593 14608 5627
rect 14556 5584 14608 5593
rect 19156 5584 19208 5636
rect 13268 5559 13320 5568
rect 13268 5525 13277 5559
rect 13277 5525 13311 5559
rect 13311 5525 13320 5559
rect 13268 5516 13320 5525
rect 14096 5516 14148 5568
rect 19064 5516 19116 5568
rect 19616 5652 19668 5704
rect 19708 5627 19760 5636
rect 19708 5593 19717 5627
rect 19717 5593 19751 5627
rect 19751 5593 19760 5627
rect 19708 5584 19760 5593
rect 20260 5720 20312 5772
rect 22284 5763 22336 5772
rect 22284 5729 22293 5763
rect 22293 5729 22327 5763
rect 22327 5729 22336 5763
rect 22284 5720 22336 5729
rect 22652 5720 22704 5772
rect 20812 5652 20864 5704
rect 21272 5652 21324 5704
rect 21364 5652 21416 5704
rect 21824 5652 21876 5704
rect 23204 5720 23256 5772
rect 21180 5516 21232 5568
rect 25228 5516 25280 5568
rect 26424 5516 26476 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 3516 5312 3568 5364
rect 4620 5312 4672 5364
rect 11060 5312 11112 5364
rect 1400 5176 1452 5228
rect 7012 5244 7064 5296
rect 8852 5244 8904 5296
rect 11704 5244 11756 5296
rect 13360 5244 13412 5296
rect 13728 5244 13780 5296
rect 15752 5244 15804 5296
rect 3608 5176 3660 5228
rect 8300 5219 8352 5228
rect 3332 5040 3384 5092
rect 6736 5108 6788 5160
rect 5264 4972 5316 5024
rect 5540 4972 5592 5024
rect 8300 5185 8309 5219
rect 8309 5185 8343 5219
rect 8343 5185 8352 5219
rect 8300 5176 8352 5185
rect 8576 5151 8628 5160
rect 8576 5117 8585 5151
rect 8585 5117 8619 5151
rect 8619 5117 8628 5151
rect 8576 5108 8628 5117
rect 9864 5176 9916 5228
rect 10324 5176 10376 5228
rect 10968 5219 11020 5228
rect 10968 5185 10977 5219
rect 10977 5185 11011 5219
rect 11011 5185 11020 5219
rect 10968 5176 11020 5185
rect 11152 5176 11204 5228
rect 19984 5312 20036 5364
rect 20168 5312 20220 5364
rect 22284 5312 22336 5364
rect 22376 5312 22428 5364
rect 17040 5287 17092 5296
rect 17040 5253 17049 5287
rect 17049 5253 17083 5287
rect 17083 5253 17092 5287
rect 17040 5244 17092 5253
rect 17224 5244 17276 5296
rect 17960 5244 18012 5296
rect 19340 5244 19392 5296
rect 19524 5244 19576 5296
rect 20260 5244 20312 5296
rect 21548 5244 21600 5296
rect 21640 5244 21692 5296
rect 22192 5287 22244 5296
rect 22192 5253 22201 5287
rect 22201 5253 22235 5287
rect 22235 5253 22244 5287
rect 22192 5244 22244 5253
rect 22560 5244 22612 5296
rect 18236 5176 18288 5228
rect 19156 5176 19208 5228
rect 19708 5176 19760 5228
rect 21088 5219 21140 5228
rect 21088 5185 21097 5219
rect 21097 5185 21131 5219
rect 21131 5185 21140 5219
rect 21088 5176 21140 5185
rect 12164 5108 12216 5160
rect 14096 5108 14148 5160
rect 14188 5108 14240 5160
rect 15476 5108 15528 5160
rect 16488 5108 16540 5160
rect 17868 5151 17920 5160
rect 17868 5117 17877 5151
rect 17877 5117 17911 5151
rect 17911 5117 17920 5151
rect 17868 5108 17920 5117
rect 18604 5108 18656 5160
rect 19432 5108 19484 5160
rect 23112 5176 23164 5228
rect 26148 5244 26200 5296
rect 26424 5219 26476 5228
rect 23020 5108 23072 5160
rect 26424 5185 26433 5219
rect 26433 5185 26467 5219
rect 26467 5185 26476 5219
rect 26424 5176 26476 5185
rect 37924 5176 37976 5228
rect 38108 5108 38160 5160
rect 13176 5040 13228 5092
rect 15200 5083 15252 5092
rect 15200 5049 15209 5083
rect 15209 5049 15243 5083
rect 15243 5049 15252 5083
rect 15200 5040 15252 5049
rect 18144 5040 18196 5092
rect 20352 5040 20404 5092
rect 21548 5040 21600 5092
rect 21916 5040 21968 5092
rect 10416 4972 10468 5024
rect 14188 4972 14240 5024
rect 18236 4972 18288 5024
rect 18328 4972 18380 5024
rect 21732 4972 21784 5024
rect 29460 4972 29512 5024
rect 33048 4972 33100 5024
rect 38200 5015 38252 5024
rect 38200 4981 38209 5015
rect 38209 4981 38243 5015
rect 38243 4981 38252 5015
rect 38200 4972 38252 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 3148 4768 3200 4820
rect 3976 4768 4028 4820
rect 3700 4700 3752 4752
rect 7380 4768 7432 4820
rect 13268 4768 13320 4820
rect 13360 4700 13412 4752
rect 1584 4632 1636 4684
rect 3332 4632 3384 4684
rect 5264 4632 5316 4684
rect 7104 4632 7156 4684
rect 9404 4632 9456 4684
rect 11152 4632 11204 4684
rect 16028 4743 16080 4752
rect 16028 4709 16037 4743
rect 16037 4709 16071 4743
rect 16071 4709 16080 4743
rect 16028 4700 16080 4709
rect 3608 4564 3660 4616
rect 11060 4564 11112 4616
rect 14188 4632 14240 4684
rect 17040 4768 17092 4820
rect 23848 4811 23900 4820
rect 23848 4777 23857 4811
rect 23857 4777 23891 4811
rect 23891 4777 23900 4811
rect 23848 4768 23900 4777
rect 17224 4700 17276 4752
rect 17592 4700 17644 4752
rect 18236 4675 18288 4684
rect 13728 4564 13780 4616
rect 7932 4496 7984 4548
rect 8116 4539 8168 4548
rect 8116 4505 8125 4539
rect 8125 4505 8159 4539
rect 8159 4505 8168 4539
rect 8116 4496 8168 4505
rect 12164 4496 12216 4548
rect 13636 4496 13688 4548
rect 15568 4496 15620 4548
rect 3516 4428 3568 4480
rect 4620 4428 4672 4480
rect 6000 4428 6052 4480
rect 9680 4428 9732 4480
rect 9956 4428 10008 4480
rect 11428 4471 11480 4480
rect 11428 4437 11437 4471
rect 11437 4437 11471 4471
rect 11471 4437 11480 4471
rect 11428 4428 11480 4437
rect 13176 4428 13228 4480
rect 16580 4496 16632 4548
rect 18236 4641 18245 4675
rect 18245 4641 18279 4675
rect 18279 4641 18288 4675
rect 18236 4632 18288 4641
rect 18512 4675 18564 4684
rect 18512 4641 18521 4675
rect 18521 4641 18555 4675
rect 18555 4641 18564 4675
rect 18512 4632 18564 4641
rect 18880 4632 18932 4684
rect 18052 4428 18104 4480
rect 18328 4539 18380 4548
rect 18328 4505 18337 4539
rect 18337 4505 18371 4539
rect 18371 4505 18380 4539
rect 20352 4564 20404 4616
rect 20536 4607 20588 4616
rect 20536 4573 20545 4607
rect 20545 4573 20579 4607
rect 20579 4573 20588 4607
rect 20536 4564 20588 4573
rect 20812 4564 20864 4616
rect 21180 4607 21232 4616
rect 21180 4573 21189 4607
rect 21189 4573 21223 4607
rect 21223 4573 21232 4607
rect 21180 4564 21232 4573
rect 18328 4496 18380 4505
rect 19708 4496 19760 4548
rect 20168 4496 20220 4548
rect 20260 4496 20312 4548
rect 23112 4607 23164 4616
rect 23112 4573 23121 4607
rect 23121 4573 23155 4607
rect 23155 4573 23164 4607
rect 23112 4564 23164 4573
rect 23756 4607 23808 4616
rect 23756 4573 23765 4607
rect 23765 4573 23799 4607
rect 23799 4573 23808 4607
rect 23756 4564 23808 4573
rect 24400 4564 24452 4616
rect 27804 4564 27856 4616
rect 37740 4564 37792 4616
rect 23572 4496 23624 4548
rect 19800 4428 19852 4480
rect 20352 4428 20404 4480
rect 20720 4428 20772 4480
rect 22284 4428 22336 4480
rect 38016 4428 38068 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 1676 4199 1728 4208
rect 1676 4165 1685 4199
rect 1685 4165 1719 4199
rect 1719 4165 1728 4199
rect 1676 4156 1728 4165
rect 3516 4156 3568 4208
rect 4620 4156 4672 4208
rect 2044 4088 2096 4140
rect 3332 4131 3384 4140
rect 3332 4097 3341 4131
rect 3341 4097 3375 4131
rect 3375 4097 3384 4131
rect 3332 4088 3384 4097
rect 7104 4156 7156 4208
rect 6552 4131 6604 4140
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 6552 4088 6604 4097
rect 8300 4224 8352 4276
rect 9220 4224 9272 4276
rect 10508 4224 10560 4276
rect 11428 4224 11480 4276
rect 9588 4156 9640 4208
rect 9680 4156 9732 4208
rect 9404 4131 9456 4140
rect 9404 4097 9413 4131
rect 9413 4097 9447 4131
rect 9447 4097 9456 4131
rect 9404 4088 9456 4097
rect 11520 4088 11572 4140
rect 13452 4156 13504 4208
rect 13820 4156 13872 4208
rect 14004 4156 14056 4208
rect 16580 4156 16632 4208
rect 17408 4156 17460 4208
rect 19156 4224 19208 4276
rect 19616 4224 19668 4276
rect 23112 4224 23164 4276
rect 23664 4224 23716 4276
rect 24400 4224 24452 4276
rect 6460 4020 6512 4072
rect 8116 4020 8168 4072
rect 12532 4020 12584 4072
rect 5448 3952 5500 4004
rect 5908 3952 5960 4004
rect 11612 3952 11664 4004
rect 12072 3995 12124 4004
rect 3976 3884 4028 3936
rect 4620 3884 4672 3936
rect 5540 3884 5592 3936
rect 5632 3884 5684 3936
rect 7104 3884 7156 3936
rect 9864 3884 9916 3936
rect 11704 3884 11756 3936
rect 12072 3961 12081 3995
rect 12081 3961 12115 3995
rect 12115 3961 12124 3995
rect 12072 3952 12124 3961
rect 12164 3952 12216 4004
rect 14832 4088 14884 4140
rect 15200 4020 15252 4072
rect 15476 4088 15528 4140
rect 16212 4131 16264 4140
rect 16212 4097 16221 4131
rect 16221 4097 16255 4131
rect 16255 4097 16264 4131
rect 16212 4088 16264 4097
rect 16764 4088 16816 4140
rect 18236 4088 18288 4140
rect 20812 4156 20864 4208
rect 23204 4156 23256 4208
rect 16856 4063 16908 4072
rect 16856 4029 16865 4063
rect 16865 4029 16899 4063
rect 16899 4029 16908 4063
rect 16856 4020 16908 4029
rect 14556 3952 14608 4004
rect 16028 3952 16080 4004
rect 16120 3952 16172 4004
rect 18144 4020 18196 4072
rect 19984 4131 20036 4140
rect 19984 4097 19993 4131
rect 19993 4097 20027 4131
rect 20027 4097 20036 4131
rect 19984 4088 20036 4097
rect 20260 4088 20312 4140
rect 22008 4131 22060 4140
rect 22008 4097 22017 4131
rect 22017 4097 22051 4131
rect 22051 4097 22060 4131
rect 22008 4088 22060 4097
rect 22284 4088 22336 4140
rect 23572 4088 23624 4140
rect 24676 4131 24728 4140
rect 24676 4097 24685 4131
rect 24685 4097 24719 4131
rect 24719 4097 24728 4131
rect 24676 4088 24728 4097
rect 26056 4131 26108 4140
rect 20812 4020 20864 4072
rect 21548 4020 21600 4072
rect 22744 3995 22796 4004
rect 12624 3884 12676 3936
rect 12992 3884 13044 3936
rect 22744 3961 22753 3995
rect 22753 3961 22787 3995
rect 22787 3961 22796 3995
rect 22744 3952 22796 3961
rect 26056 4097 26065 4131
rect 26065 4097 26099 4131
rect 26099 4097 26108 4131
rect 26056 4088 26108 4097
rect 38292 4131 38344 4140
rect 38292 4097 38301 4131
rect 38301 4097 38335 4131
rect 38335 4097 38344 4131
rect 38292 4088 38344 4097
rect 20996 3884 21048 3936
rect 21088 3884 21140 3936
rect 22560 3884 22612 3936
rect 25780 3952 25832 4004
rect 31392 3952 31444 4004
rect 23388 3927 23440 3936
rect 23388 3893 23397 3927
rect 23397 3893 23431 3927
rect 23431 3893 23440 3927
rect 23388 3884 23440 3893
rect 25320 3927 25372 3936
rect 25320 3893 25329 3927
rect 25329 3893 25363 3927
rect 25363 3893 25372 3927
rect 25320 3884 25372 3893
rect 27436 3884 27488 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 6552 3680 6604 3732
rect 3884 3612 3936 3664
rect 11612 3680 11664 3732
rect 11704 3680 11756 3732
rect 13360 3680 13412 3732
rect 13452 3680 13504 3732
rect 16028 3723 16080 3732
rect 4068 3544 4120 3596
rect 5816 3544 5868 3596
rect 4620 3476 4672 3528
rect 4896 3519 4948 3528
rect 4896 3485 4905 3519
rect 4905 3485 4939 3519
rect 4939 3485 4948 3519
rect 4896 3476 4948 3485
rect 4160 3408 4212 3460
rect 4344 3451 4396 3460
rect 4344 3417 4353 3451
rect 4353 3417 4387 3451
rect 4387 3417 4396 3451
rect 4344 3408 4396 3417
rect 3148 3340 3200 3392
rect 4620 3340 4672 3392
rect 5172 3340 5224 3392
rect 5540 3383 5592 3392
rect 5540 3349 5549 3383
rect 5549 3349 5583 3383
rect 5583 3349 5592 3383
rect 5540 3340 5592 3349
rect 8116 3612 8168 3664
rect 8300 3544 8352 3596
rect 8392 3544 8444 3596
rect 8668 3544 8720 3596
rect 9772 3544 9824 3596
rect 10876 3544 10928 3596
rect 11152 3544 11204 3596
rect 12532 3612 12584 3664
rect 14188 3612 14240 3664
rect 16028 3689 16037 3723
rect 16037 3689 16071 3723
rect 16071 3689 16080 3723
rect 16028 3680 16080 3689
rect 17592 3680 17644 3732
rect 17776 3680 17828 3732
rect 18328 3680 18380 3732
rect 19064 3680 19116 3732
rect 19524 3680 19576 3732
rect 22192 3680 22244 3732
rect 22836 3723 22888 3732
rect 22836 3689 22845 3723
rect 22845 3689 22879 3723
rect 22879 3689 22888 3723
rect 22836 3680 22888 3689
rect 24584 3680 24636 3732
rect 25228 3680 25280 3732
rect 37464 3723 37516 3732
rect 37464 3689 37473 3723
rect 37473 3689 37507 3723
rect 37507 3689 37516 3723
rect 37464 3680 37516 3689
rect 38108 3723 38160 3732
rect 38108 3689 38117 3723
rect 38117 3689 38151 3723
rect 38151 3689 38160 3723
rect 38108 3680 38160 3689
rect 13636 3544 13688 3596
rect 13728 3544 13780 3596
rect 16856 3544 16908 3596
rect 9312 3519 9364 3528
rect 9312 3485 9321 3519
rect 9321 3485 9355 3519
rect 9355 3485 9364 3519
rect 9312 3476 9364 3485
rect 9864 3476 9916 3528
rect 13084 3476 13136 3528
rect 13360 3476 13412 3528
rect 18236 3612 18288 3664
rect 7104 3451 7156 3460
rect 7104 3417 7113 3451
rect 7113 3417 7147 3451
rect 7147 3417 7156 3451
rect 7104 3408 7156 3417
rect 9128 3408 9180 3460
rect 7012 3340 7064 3392
rect 7196 3340 7248 3392
rect 9680 3340 9732 3392
rect 9772 3340 9824 3392
rect 10140 3340 10192 3392
rect 10232 3340 10284 3392
rect 11152 3408 11204 3460
rect 11428 3408 11480 3460
rect 13544 3408 13596 3460
rect 14832 3408 14884 3460
rect 16396 3408 16448 3460
rect 16580 3451 16632 3460
rect 16580 3417 16589 3451
rect 16589 3417 16623 3451
rect 16623 3417 16632 3451
rect 16580 3408 16632 3417
rect 17776 3408 17828 3460
rect 21088 3544 21140 3596
rect 23388 3612 23440 3664
rect 27252 3612 27304 3664
rect 18696 3519 18748 3528
rect 18696 3485 18705 3519
rect 18705 3485 18739 3519
rect 18739 3485 18748 3519
rect 18696 3476 18748 3485
rect 18512 3408 18564 3460
rect 19524 3476 19576 3528
rect 20720 3476 20772 3528
rect 21456 3519 21508 3528
rect 21456 3485 21465 3519
rect 21465 3485 21499 3519
rect 21499 3485 21508 3519
rect 21456 3476 21508 3485
rect 22100 3519 22152 3528
rect 22100 3485 22109 3519
rect 22109 3485 22143 3519
rect 22143 3485 22152 3519
rect 22100 3476 22152 3485
rect 22652 3476 22704 3528
rect 23572 3476 23624 3528
rect 24676 3476 24728 3528
rect 25780 3476 25832 3528
rect 37648 3519 37700 3528
rect 37648 3485 37657 3519
rect 37657 3485 37691 3519
rect 37691 3485 37700 3519
rect 37648 3476 37700 3485
rect 38108 3476 38160 3528
rect 20628 3408 20680 3460
rect 22284 3408 22336 3460
rect 24032 3408 24084 3460
rect 26148 3408 26200 3460
rect 33600 3408 33652 3460
rect 20904 3383 20956 3392
rect 20904 3349 20913 3383
rect 20913 3349 20947 3383
rect 20947 3349 20956 3383
rect 21548 3383 21600 3392
rect 20904 3340 20956 3349
rect 21548 3349 21557 3383
rect 21557 3349 21591 3383
rect 21591 3349 21600 3383
rect 21548 3340 21600 3349
rect 21916 3340 21968 3392
rect 23572 3340 23624 3392
rect 24400 3340 24452 3392
rect 26240 3340 26292 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 3424 3179 3476 3188
rect 3424 3145 3433 3179
rect 3433 3145 3467 3179
rect 3467 3145 3476 3179
rect 3424 3136 3476 3145
rect 4712 3136 4764 3188
rect 5540 3136 5592 3188
rect 1952 3068 2004 3120
rect 3792 3068 3844 3120
rect 4160 3068 4212 3120
rect 5356 3068 5408 3120
rect 2504 3000 2556 3052
rect 3700 3000 3752 3052
rect 3976 3043 4028 3052
rect 3976 3009 3985 3043
rect 3985 3009 4019 3043
rect 4019 3009 4028 3043
rect 3976 3000 4028 3009
rect 4988 3000 5040 3052
rect 5172 3000 5224 3052
rect 8116 3068 8168 3120
rect 7564 3000 7616 3052
rect 7748 3043 7800 3052
rect 7748 3009 7757 3043
rect 7757 3009 7791 3043
rect 7791 3009 7800 3043
rect 7748 3000 7800 3009
rect 4068 2907 4120 2916
rect 4068 2873 4077 2907
rect 4077 2873 4111 2907
rect 4111 2873 4120 2907
rect 4068 2864 4120 2873
rect 6920 2932 6972 2984
rect 9496 3068 9548 3120
rect 9680 3068 9732 3120
rect 10692 3068 10744 3120
rect 8392 3000 8444 3052
rect 11152 3000 11204 3052
rect 11888 3000 11940 3052
rect 12164 3043 12216 3052
rect 12164 3009 12173 3043
rect 12173 3009 12207 3043
rect 12207 3009 12216 3043
rect 12164 3000 12216 3009
rect 13360 3068 13412 3120
rect 13452 3111 13504 3120
rect 13452 3077 13461 3111
rect 13461 3077 13495 3111
rect 13495 3077 13504 3111
rect 13452 3068 13504 3077
rect 15476 3068 15528 3120
rect 20812 3136 20864 3188
rect 16580 3068 16632 3120
rect 17684 3068 17736 3120
rect 19984 3068 20036 3120
rect 20076 3068 20128 3120
rect 20628 3068 20680 3120
rect 20720 3068 20772 3120
rect 22008 3136 22060 3188
rect 22652 3179 22704 3188
rect 22652 3145 22661 3179
rect 22661 3145 22695 3179
rect 22695 3145 22704 3179
rect 22652 3136 22704 3145
rect 16672 3000 16724 3052
rect 18052 3043 18104 3052
rect 18052 3009 18061 3043
rect 18061 3009 18095 3043
rect 18095 3009 18104 3043
rect 18052 3000 18104 3009
rect 8668 2932 8720 2984
rect 9956 2932 10008 2984
rect 664 2796 716 2848
rect 2688 2839 2740 2848
rect 2688 2805 2697 2839
rect 2697 2805 2731 2839
rect 2731 2805 2740 2839
rect 2688 2796 2740 2805
rect 6000 2796 6052 2848
rect 8484 2796 8536 2848
rect 14004 2932 14056 2984
rect 10324 2864 10376 2916
rect 11612 2796 11664 2848
rect 16304 2864 16356 2916
rect 18604 2932 18656 2984
rect 18788 2975 18840 2984
rect 18788 2941 18797 2975
rect 18797 2941 18831 2975
rect 18831 2941 18840 2975
rect 18788 2932 18840 2941
rect 18880 2932 18932 2984
rect 19248 2932 19300 2984
rect 22468 3000 22520 3052
rect 21916 2932 21968 2984
rect 23204 3000 23256 3052
rect 24584 3000 24636 3052
rect 25412 3043 25464 3052
rect 22928 2932 22980 2984
rect 25412 3009 25421 3043
rect 25421 3009 25455 3043
rect 25455 3009 25464 3043
rect 25412 3000 25464 3009
rect 27160 3136 27212 3188
rect 27252 3111 27304 3120
rect 27252 3077 27261 3111
rect 27261 3077 27295 3111
rect 27295 3077 27304 3111
rect 27252 3068 27304 3077
rect 36728 3068 36780 3120
rect 26240 3000 26292 3052
rect 33600 3043 33652 3052
rect 33600 3009 33609 3043
rect 33609 3009 33643 3043
rect 33643 3009 33652 3043
rect 33600 3000 33652 3009
rect 36912 3043 36964 3052
rect 36912 3009 36921 3043
rect 36921 3009 36955 3043
rect 36955 3009 36964 3043
rect 36912 3000 36964 3009
rect 38292 3043 38344 3052
rect 38292 3009 38301 3043
rect 38301 3009 38335 3043
rect 38335 3009 38344 3043
rect 38292 3000 38344 3009
rect 17592 2864 17644 2916
rect 20260 2864 20312 2916
rect 22652 2864 22704 2916
rect 22744 2864 22796 2916
rect 30748 2932 30800 2984
rect 25872 2864 25924 2916
rect 30564 2864 30616 2916
rect 15108 2796 15160 2848
rect 17960 2796 18012 2848
rect 21272 2796 21324 2848
rect 22100 2796 22152 2848
rect 23480 2796 23532 2848
rect 24492 2796 24544 2848
rect 33508 2796 33560 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 1492 2592 1544 2644
rect 9128 2592 9180 2644
rect 11244 2592 11296 2644
rect 11980 2592 12032 2644
rect 20 2524 72 2576
rect 7748 2524 7800 2576
rect 9312 2524 9364 2576
rect 11060 2524 11112 2576
rect 2228 2388 2280 2440
rect 3056 2431 3108 2440
rect 3056 2397 3065 2431
rect 3065 2397 3099 2431
rect 3099 2397 3108 2431
rect 3056 2388 3108 2397
rect 5632 2456 5684 2508
rect 6920 2456 6972 2508
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 7748 2431 7800 2440
rect 7748 2397 7757 2431
rect 7757 2397 7791 2431
rect 7791 2397 7800 2431
rect 7748 2388 7800 2397
rect 1676 2363 1728 2372
rect 1676 2329 1685 2363
rect 1685 2329 1719 2363
rect 1719 2329 1728 2363
rect 1676 2320 1728 2329
rect 9404 2320 9456 2372
rect 2504 2295 2556 2304
rect 2504 2261 2513 2295
rect 2513 2261 2547 2295
rect 2547 2261 2556 2295
rect 2504 2252 2556 2261
rect 3976 2295 4028 2304
rect 3976 2261 3985 2295
rect 3985 2261 4019 2295
rect 4019 2261 4028 2295
rect 3976 2252 4028 2261
rect 4712 2295 4764 2304
rect 4712 2261 4721 2295
rect 4721 2261 4755 2295
rect 4755 2261 4764 2295
rect 4712 2252 4764 2261
rect 5172 2252 5224 2304
rect 7840 2295 7892 2304
rect 7840 2261 7849 2295
rect 7849 2261 7883 2295
rect 7883 2261 7892 2295
rect 7840 2252 7892 2261
rect 8484 2295 8536 2304
rect 8484 2261 8493 2295
rect 8493 2261 8527 2295
rect 8527 2261 8536 2295
rect 8484 2252 8536 2261
rect 10140 2388 10192 2440
rect 10876 2431 10928 2440
rect 10876 2397 10885 2431
rect 10885 2397 10919 2431
rect 10919 2397 10928 2431
rect 10876 2388 10928 2397
rect 13912 2524 13964 2576
rect 13728 2456 13780 2508
rect 15936 2592 15988 2644
rect 16764 2592 16816 2644
rect 17316 2592 17368 2644
rect 17408 2592 17460 2644
rect 20168 2592 20220 2644
rect 21364 2592 21416 2644
rect 25228 2592 25280 2644
rect 27804 2635 27856 2644
rect 27804 2601 27813 2635
rect 27813 2601 27847 2635
rect 27847 2601 27856 2635
rect 27804 2592 27856 2601
rect 28632 2635 28684 2644
rect 28632 2601 28641 2635
rect 28641 2601 28675 2635
rect 28675 2601 28684 2635
rect 28632 2592 28684 2601
rect 30104 2592 30156 2644
rect 16120 2524 16172 2576
rect 16580 2456 16632 2508
rect 22744 2524 22796 2576
rect 23388 2567 23440 2576
rect 23388 2533 23397 2567
rect 23397 2533 23431 2567
rect 23431 2533 23440 2567
rect 23388 2524 23440 2533
rect 27436 2524 27488 2576
rect 13452 2431 13504 2440
rect 13452 2397 13461 2431
rect 13461 2397 13495 2431
rect 13495 2397 13504 2431
rect 13452 2388 13504 2397
rect 21548 2456 21600 2508
rect 18236 2431 18288 2440
rect 11520 2320 11572 2372
rect 11612 2320 11664 2372
rect 12164 2320 12216 2372
rect 10968 2252 11020 2304
rect 13544 2252 13596 2304
rect 14832 2252 14884 2304
rect 16764 2320 16816 2372
rect 18236 2397 18245 2431
rect 18245 2397 18279 2431
rect 18279 2397 18288 2431
rect 18236 2388 18288 2397
rect 17408 2252 17460 2304
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 20628 2388 20680 2440
rect 19340 2320 19392 2372
rect 22008 2388 22060 2440
rect 22652 2431 22704 2440
rect 22652 2397 22661 2431
rect 22661 2397 22695 2431
rect 22695 2397 22704 2431
rect 22652 2388 22704 2397
rect 24124 2456 24176 2508
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 25228 2431 25280 2440
rect 25228 2397 25237 2431
rect 25237 2397 25271 2431
rect 25271 2397 25280 2431
rect 25228 2388 25280 2397
rect 25872 2388 25924 2440
rect 27344 2431 27396 2440
rect 27344 2397 27353 2431
rect 27353 2397 27387 2431
rect 27387 2397 27396 2431
rect 27344 2388 27396 2397
rect 27068 2320 27120 2372
rect 29460 2388 29512 2440
rect 30288 2388 30340 2440
rect 31576 2388 31628 2440
rect 33048 2388 33100 2440
rect 34796 2388 34848 2440
rect 38016 2431 38068 2440
rect 38016 2397 38025 2431
rect 38025 2397 38059 2431
rect 38059 2397 38068 2431
rect 38016 2388 38068 2397
rect 28356 2320 28408 2372
rect 22192 2252 22244 2304
rect 22560 2252 22612 2304
rect 24676 2295 24728 2304
rect 24676 2261 24685 2295
rect 24685 2261 24719 2295
rect 24719 2261 24728 2295
rect 24676 2252 24728 2261
rect 25136 2252 25188 2304
rect 25780 2252 25832 2304
rect 27160 2295 27212 2304
rect 27160 2261 27169 2295
rect 27169 2261 27203 2295
rect 27203 2261 27212 2295
rect 27160 2252 27212 2261
rect 29644 2252 29696 2304
rect 32864 2252 32916 2304
rect 34796 2252 34848 2304
rect 36084 2252 36136 2304
rect 39304 2252 39356 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 3976 2048 4028 2100
rect 11980 2048 12032 2100
rect 18236 2048 18288 2100
rect 22376 2048 22428 2100
rect 7840 1980 7892 2032
rect 15568 1980 15620 2032
rect 16764 1980 16816 2032
rect 25320 1980 25372 2032
rect 4988 1912 5040 1964
rect 14464 1912 14516 1964
rect 15936 1912 15988 1964
rect 19156 1912 19208 1964
rect 8484 1844 8536 1896
rect 12532 1844 12584 1896
rect 10600 1776 10652 1828
rect 24676 1844 24728 1896
rect 14464 1708 14516 1760
rect 20076 1776 20128 1828
rect 18052 1708 18104 1760
rect 27344 1708 27396 1760
rect 12532 1640 12584 1692
rect 15660 1640 15712 1692
rect 16948 1640 17000 1692
rect 22652 1640 22704 1692
rect 23848 1640 23900 1692
rect 25412 1640 25464 1692
rect 13544 1572 13596 1624
rect 22928 1572 22980 1624
rect 7288 1504 7340 1556
rect 20444 1504 20496 1556
rect 4712 1436 4764 1488
rect 18788 1436 18840 1488
<< metal2 >>
rect 18 39200 74 39800
rect 1306 39200 1362 39800
rect 2594 39200 2650 39800
rect 3238 39200 3294 39800
rect 4526 39200 4582 39800
rect 5814 39200 5870 39800
rect 6458 39200 6514 39800
rect 7746 39200 7802 39800
rect 9034 39200 9090 39800
rect 9678 39200 9734 39800
rect 10966 39200 11022 39800
rect 12254 39200 12310 39800
rect 13542 39200 13598 39800
rect 14186 39200 14242 39800
rect 15474 39200 15530 39800
rect 16762 39200 16818 39800
rect 17406 39200 17462 39800
rect 18694 39200 18750 39800
rect 19982 39200 20038 39800
rect 21270 39200 21326 39800
rect 21914 39200 21970 39800
rect 23202 39200 23258 39800
rect 24490 39200 24546 39800
rect 25134 39200 25190 39800
rect 26422 39200 26478 39800
rect 27710 39200 27766 39800
rect 28354 39200 28410 39800
rect 29642 39200 29698 39800
rect 30930 39200 30986 39800
rect 32218 39200 32274 39800
rect 32862 39200 32918 39800
rect 34150 39200 34206 39800
rect 34256 39222 34468 39250
rect 32 36854 60 39200
rect 20 36848 72 36854
rect 20 36790 72 36796
rect 1320 36174 1348 39200
rect 1766 38856 1822 38865
rect 1766 38791 1822 38800
rect 1674 38176 1730 38185
rect 1674 38111 1730 38120
rect 1688 36922 1716 38111
rect 1780 37466 1808 38791
rect 1768 37460 1820 37466
rect 1768 37402 1820 37408
rect 2412 37256 2464 37262
rect 2412 37198 2464 37204
rect 2608 37210 2636 39200
rect 2780 37256 2832 37262
rect 2608 37204 2780 37210
rect 2608 37198 2832 37204
rect 1676 36916 1728 36922
rect 1676 36858 1728 36864
rect 2320 36576 2372 36582
rect 2320 36518 2372 36524
rect 1308 36168 1360 36174
rect 1308 36110 1360 36116
rect 1584 35624 1636 35630
rect 1584 35566 1636 35572
rect 1596 35465 1624 35566
rect 1582 35456 1638 35465
rect 1582 35391 1638 35400
rect 1768 35080 1820 35086
rect 1768 35022 1820 35028
rect 1860 35080 1912 35086
rect 1860 35022 1912 35028
rect 1780 34785 1808 35022
rect 1766 34776 1822 34785
rect 1766 34711 1822 34720
rect 1766 33416 1822 33425
rect 1766 33351 1768 33360
rect 1820 33351 1822 33360
rect 1768 33322 1820 33328
rect 1768 32224 1820 32230
rect 1768 32166 1820 32172
rect 1780 32065 1808 32166
rect 1766 32056 1822 32065
rect 1766 31991 1822 32000
rect 1872 31890 1900 35022
rect 2228 32224 2280 32230
rect 2228 32166 2280 32172
rect 2240 32026 2268 32166
rect 2228 32020 2280 32026
rect 2228 31962 2280 31968
rect 1860 31884 1912 31890
rect 1860 31826 1912 31832
rect 1584 31816 1636 31822
rect 1584 31758 1636 31764
rect 1596 31385 1624 31758
rect 1582 31376 1638 31385
rect 1582 31311 1638 31320
rect 2332 30734 2360 36518
rect 2424 33862 2452 37198
rect 2608 37182 2820 37198
rect 3252 37126 3280 39200
rect 4540 37754 4568 39200
rect 4540 37726 4660 37754
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4632 37262 4660 37726
rect 5828 37262 5856 39200
rect 6472 37262 6500 39200
rect 3976 37256 4028 37262
rect 3976 37198 4028 37204
rect 4620 37256 4672 37262
rect 4620 37198 4672 37204
rect 5816 37256 5868 37262
rect 5816 37198 5868 37204
rect 6460 37256 6512 37262
rect 6460 37198 6512 37204
rect 3240 37120 3292 37126
rect 3240 37062 3292 37068
rect 2502 36816 2558 36825
rect 2502 36751 2504 36760
rect 2556 36751 2558 36760
rect 2504 36722 2556 36728
rect 2596 36032 2648 36038
rect 2596 35974 2648 35980
rect 2412 33856 2464 33862
rect 2412 33798 2464 33804
rect 2608 30802 2636 35974
rect 3988 35290 4016 37198
rect 6828 37188 6880 37194
rect 6828 37130 6880 37136
rect 4712 37120 4764 37126
rect 4712 37062 4764 37068
rect 6368 37120 6420 37126
rect 6368 37062 6420 37068
rect 6552 37120 6604 37126
rect 6552 37062 6604 37068
rect 4068 36712 4120 36718
rect 4068 36654 4120 36660
rect 3976 35284 4028 35290
rect 3976 35226 4028 35232
rect 2688 34944 2740 34950
rect 2688 34886 2740 34892
rect 2596 30796 2648 30802
rect 2596 30738 2648 30744
rect 2320 30728 2372 30734
rect 2320 30670 2372 30676
rect 2700 30258 2728 34886
rect 4080 34746 4108 36654
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4068 34740 4120 34746
rect 4068 34682 4120 34688
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4724 33522 4752 37062
rect 5816 36576 5868 36582
rect 5816 36518 5868 36524
rect 5724 34604 5776 34610
rect 5724 34546 5776 34552
rect 4068 33516 4120 33522
rect 4068 33458 4120 33464
rect 4712 33516 4764 33522
rect 4712 33458 4764 33464
rect 2964 31884 3016 31890
rect 2964 31826 3016 31832
rect 2688 30252 2740 30258
rect 2688 30194 2740 30200
rect 1768 30048 1820 30054
rect 1766 30016 1768 30025
rect 1820 30016 1822 30025
rect 1766 29951 1822 29960
rect 1768 29640 1820 29646
rect 1768 29582 1820 29588
rect 1582 29064 1638 29073
rect 1582 28999 1584 29008
rect 1636 28999 1638 29008
rect 1584 28970 1636 28976
rect 1780 28665 1808 29582
rect 2780 29164 2832 29170
rect 2780 29106 2832 29112
rect 1766 28656 1822 28665
rect 756 28620 808 28626
rect 1766 28591 1822 28600
rect 756 28562 808 28568
rect 572 26988 624 26994
rect 572 26930 624 26936
rect 584 10062 612 26930
rect 664 26444 716 26450
rect 664 26386 716 26392
rect 676 12986 704 26386
rect 664 12980 716 12986
rect 664 12922 716 12928
rect 572 10056 624 10062
rect 572 9998 624 10004
rect 768 8362 796 28562
rect 1860 28552 1912 28558
rect 1860 28494 1912 28500
rect 1584 27940 1636 27946
rect 1584 27882 1636 27888
rect 1216 27056 1268 27062
rect 1216 26998 1268 27004
rect 848 26852 900 26858
rect 848 26794 900 26800
rect 860 17377 888 26794
rect 1124 26784 1176 26790
rect 1124 26726 1176 26732
rect 940 24608 992 24614
rect 940 24550 992 24556
rect 846 17368 902 17377
rect 846 17303 902 17312
rect 952 13190 980 24550
rect 1032 24132 1084 24138
rect 1032 24074 1084 24080
rect 940 13184 992 13190
rect 940 13126 992 13132
rect 1044 12442 1072 24074
rect 1136 16250 1164 26726
rect 1124 16244 1176 16250
rect 1124 16186 1176 16192
rect 1228 14890 1256 26998
rect 1400 25900 1452 25906
rect 1400 25842 1452 25848
rect 1308 25220 1360 25226
rect 1308 25162 1360 25168
rect 1216 14884 1268 14890
rect 1216 14826 1268 14832
rect 1320 13530 1348 25162
rect 1412 24993 1440 25842
rect 1398 24984 1454 24993
rect 1398 24919 1454 24928
rect 1596 20602 1624 27882
rect 1872 27713 1900 28494
rect 2320 28416 2372 28422
rect 2320 28358 2372 28364
rect 1952 28076 2004 28082
rect 1952 28018 2004 28024
rect 1858 27704 1914 27713
rect 1858 27639 1914 27648
rect 1860 27464 1912 27470
rect 1964 27452 1992 28018
rect 2044 27872 2096 27878
rect 2044 27814 2096 27820
rect 2056 27713 2084 27814
rect 2042 27704 2098 27713
rect 2042 27639 2098 27648
rect 1912 27424 1992 27452
rect 1860 27406 1912 27412
rect 1872 26994 1900 27406
rect 1952 27328 2004 27334
rect 1952 27270 2004 27276
rect 2136 27328 2188 27334
rect 2136 27270 2188 27276
rect 1860 26988 1912 26994
rect 1860 26930 1912 26936
rect 1964 26761 1992 27270
rect 1950 26752 2006 26761
rect 1950 26687 2006 26696
rect 1858 26480 1914 26489
rect 1858 26415 1914 26424
rect 1872 26382 1900 26415
rect 1860 26376 1912 26382
rect 1860 26318 1912 26324
rect 1952 26308 2004 26314
rect 1952 26250 2004 26256
rect 1766 25256 1822 25265
rect 1766 25191 1822 25200
rect 1780 25158 1808 25191
rect 1768 25152 1820 25158
rect 1768 25094 1820 25100
rect 1860 25152 1912 25158
rect 1860 25094 1912 25100
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1780 23905 1808 24006
rect 1766 23896 1822 23905
rect 1766 23831 1822 23840
rect 1676 23724 1728 23730
rect 1676 23666 1728 23672
rect 1688 23225 1716 23666
rect 1674 23216 1730 23225
rect 1674 23151 1730 23160
rect 1872 23050 1900 25094
rect 1860 23044 1912 23050
rect 1860 22986 1912 22992
rect 1676 22976 1728 22982
rect 1676 22918 1728 22924
rect 1584 20596 1636 20602
rect 1584 20538 1636 20544
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1308 13524 1360 13530
rect 1308 13466 1360 13472
rect 1320 12458 1348 13466
rect 1032 12436 1084 12442
rect 1320 12430 1440 12458
rect 1032 12378 1084 12384
rect 1412 12306 1440 12430
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 756 8356 808 8362
rect 756 8298 808 8304
rect 1398 7576 1454 7585
rect 1398 7511 1454 7520
rect 1412 7478 1440 7511
rect 1400 7472 1452 7478
rect 1400 7414 1452 7420
rect 1398 5536 1454 5545
rect 1398 5471 1454 5480
rect 1412 5234 1440 5471
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 664 2848 716 2854
rect 664 2790 716 2796
rect 20 2576 72 2582
rect 20 2518 72 2524
rect 32 800 60 2518
rect 676 800 704 2790
rect 1504 2650 1532 18566
rect 1688 18426 1716 22918
rect 1860 22772 1912 22778
rect 1860 22714 1912 22720
rect 1766 21856 1822 21865
rect 1766 21791 1822 21800
rect 1780 21146 1808 21791
rect 1768 21140 1820 21146
rect 1768 21082 1820 21088
rect 1872 19786 1900 22714
rect 1964 21622 1992 26250
rect 2044 25968 2096 25974
rect 2044 25910 2096 25916
rect 2056 24970 2084 25910
rect 2148 25140 2176 27270
rect 2332 25786 2360 28358
rect 2594 28112 2650 28121
rect 2594 28047 2596 28056
rect 2648 28047 2650 28056
rect 2596 28018 2648 28024
rect 2504 27464 2556 27470
rect 2504 27406 2556 27412
rect 2516 26897 2544 27406
rect 2502 26888 2558 26897
rect 2502 26823 2558 26832
rect 2504 26376 2556 26382
rect 2502 26344 2504 26353
rect 2556 26344 2558 26353
rect 2502 26279 2558 26288
rect 2688 26308 2740 26314
rect 2688 26250 2740 26256
rect 2700 25974 2728 26250
rect 2792 26217 2820 29106
rect 2872 28484 2924 28490
rect 2872 28426 2924 28432
rect 2778 26208 2834 26217
rect 2778 26143 2834 26152
rect 2884 26058 2912 28426
rect 2976 27130 3004 31826
rect 4080 29850 4108 33458
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 5356 30592 5408 30598
rect 5356 30534 5408 30540
rect 5172 30184 5224 30190
rect 5172 30126 5224 30132
rect 4988 30048 5040 30054
rect 4988 29990 5040 29996
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4068 29844 4120 29850
rect 4068 29786 4120 29792
rect 4712 29504 4764 29510
rect 4712 29446 4764 29452
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 3424 28076 3476 28082
rect 3424 28018 3476 28024
rect 4068 28076 4120 28082
rect 4068 28018 4120 28024
rect 3240 27872 3292 27878
rect 3238 27840 3240 27849
rect 3292 27840 3294 27849
rect 3238 27775 3294 27784
rect 3240 27464 3292 27470
rect 3240 27406 3292 27412
rect 2964 27124 3016 27130
rect 2964 27066 3016 27072
rect 2964 26988 3016 26994
rect 2964 26930 3016 26936
rect 2976 26382 3004 26930
rect 3056 26920 3108 26926
rect 3056 26862 3108 26868
rect 2964 26376 3016 26382
rect 2964 26318 3016 26324
rect 2792 26030 2912 26058
rect 2688 25968 2740 25974
rect 2688 25910 2740 25916
rect 2332 25758 2728 25786
rect 2596 25696 2648 25702
rect 2596 25638 2648 25644
rect 2228 25288 2280 25294
rect 2226 25256 2228 25265
rect 2280 25256 2282 25265
rect 2226 25191 2282 25200
rect 2148 25112 2360 25140
rect 2056 24942 2268 24970
rect 2044 24812 2096 24818
rect 2044 24754 2096 24760
rect 2056 22098 2084 24754
rect 2240 23746 2268 24942
rect 2148 23718 2268 23746
rect 2044 22092 2096 22098
rect 2044 22034 2096 22040
rect 1952 21616 2004 21622
rect 1952 21558 2004 21564
rect 2044 21616 2096 21622
rect 2044 21558 2096 21564
rect 1860 19780 1912 19786
rect 1860 19722 1912 19728
rect 1858 19272 1914 19281
rect 1858 19207 1914 19216
rect 1676 18420 1728 18426
rect 1676 18362 1728 18368
rect 1872 18290 1900 19207
rect 1860 18284 1912 18290
rect 1860 18226 1912 18232
rect 1768 18080 1820 18086
rect 1768 18022 1820 18028
rect 1584 17672 1636 17678
rect 1584 17614 1636 17620
rect 1596 17134 1624 17614
rect 1584 17128 1636 17134
rect 1584 17070 1636 17076
rect 1596 16590 1624 17070
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 1596 16046 1624 16526
rect 1584 16040 1636 16046
rect 1584 15982 1636 15988
rect 1596 15502 1624 15982
rect 1584 15496 1636 15502
rect 1584 15438 1636 15444
rect 1596 14958 1624 15438
rect 1584 14952 1636 14958
rect 1584 14894 1636 14900
rect 1596 14482 1624 14894
rect 1584 14476 1636 14482
rect 1584 14418 1636 14424
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 1596 12782 1624 13262
rect 1584 12776 1636 12782
rect 1584 12718 1636 12724
rect 1596 12238 1624 12718
rect 1584 12232 1636 12238
rect 1584 12174 1636 12180
rect 1596 11762 1624 12174
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 1596 11218 1624 11698
rect 1584 11212 1636 11218
rect 1584 11154 1636 11160
rect 1780 10810 1808 18022
rect 1860 17604 1912 17610
rect 1860 17546 1912 17552
rect 1872 17513 1900 17546
rect 1858 17504 1914 17513
rect 1858 17439 1914 17448
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 1860 14952 1912 14958
rect 1860 14894 1912 14900
rect 1872 11558 1900 14894
rect 1964 14346 1992 17274
rect 1952 14340 2004 14346
rect 1952 14282 2004 14288
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1596 9382 1624 9454
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 8786 1624 9318
rect 2056 9178 2084 21558
rect 2148 19922 2176 23718
rect 2228 22500 2280 22506
rect 2228 22442 2280 22448
rect 2240 21486 2268 22442
rect 2228 21480 2280 21486
rect 2228 21422 2280 21428
rect 2136 19916 2188 19922
rect 2136 19858 2188 19864
rect 2134 19272 2190 19281
rect 2134 19207 2190 19216
rect 2228 19236 2280 19242
rect 2148 15434 2176 19207
rect 2228 19178 2280 19184
rect 2240 16538 2268 19178
rect 2332 18698 2360 25112
rect 2412 24744 2464 24750
rect 2412 24686 2464 24692
rect 2424 22098 2452 24686
rect 2504 24064 2556 24070
rect 2502 24032 2504 24041
rect 2556 24032 2558 24041
rect 2502 23967 2558 23976
rect 2504 23520 2556 23526
rect 2504 23462 2556 23468
rect 2412 22092 2464 22098
rect 2412 22034 2464 22040
rect 2516 21962 2544 23462
rect 2504 21956 2556 21962
rect 2504 21898 2556 21904
rect 2504 21684 2556 21690
rect 2504 21626 2556 21632
rect 2412 21480 2464 21486
rect 2412 21422 2464 21428
rect 2424 20806 2452 21422
rect 2412 20800 2464 20806
rect 2412 20742 2464 20748
rect 2320 18692 2372 18698
rect 2320 18634 2372 18640
rect 2240 16510 2360 16538
rect 2226 16416 2282 16425
rect 2226 16351 2282 16360
rect 2136 15428 2188 15434
rect 2136 15370 2188 15376
rect 2240 15042 2268 16351
rect 2148 15014 2268 15042
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 1596 8758 1716 8786
rect 1582 8664 1638 8673
rect 1582 8599 1584 8608
rect 1636 8599 1638 8608
rect 1584 8570 1636 8576
rect 1688 8430 1716 8758
rect 1964 8634 1992 8910
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1688 7954 1716 8366
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1688 7426 1716 7890
rect 1688 7410 1808 7426
rect 1688 7404 1820 7410
rect 1688 7398 1768 7404
rect 1768 7346 1820 7352
rect 1858 7304 1914 7313
rect 1858 7239 1860 7248
rect 1912 7239 1914 7248
rect 1860 7210 1912 7216
rect 1768 6928 1820 6934
rect 1766 6896 1768 6905
rect 2148 6914 2176 15014
rect 2226 14920 2282 14929
rect 2226 14855 2282 14864
rect 2240 14006 2268 14855
rect 2332 14385 2360 16510
rect 2318 14376 2374 14385
rect 2318 14311 2374 14320
rect 2228 14000 2280 14006
rect 2228 13942 2280 13948
rect 2320 14000 2372 14006
rect 2320 13942 2372 13948
rect 2332 11218 2360 13942
rect 2320 11212 2372 11218
rect 2320 11154 2372 11160
rect 2424 6914 2452 20742
rect 2516 19122 2544 21626
rect 2608 20874 2636 25638
rect 2700 22710 2728 25758
rect 2688 22704 2740 22710
rect 2688 22646 2740 22652
rect 2686 22536 2742 22545
rect 2686 22471 2742 22480
rect 2596 20868 2648 20874
rect 2596 20810 2648 20816
rect 2700 19334 2728 22471
rect 2792 22094 2820 26030
rect 2872 25152 2924 25158
rect 2872 25094 2924 25100
rect 2884 22710 2912 25094
rect 2976 24750 3004 26318
rect 2964 24744 3016 24750
rect 2964 24686 3016 24692
rect 2964 24064 3016 24070
rect 2964 24006 3016 24012
rect 2976 22710 3004 24006
rect 2872 22704 2924 22710
rect 2872 22646 2924 22652
rect 2964 22704 3016 22710
rect 2964 22646 3016 22652
rect 2792 22066 3004 22094
rect 2872 21412 2924 21418
rect 2872 21354 2924 21360
rect 2884 20058 2912 21354
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 2780 19440 2832 19446
rect 2780 19382 2832 19388
rect 2608 19306 2728 19334
rect 2608 19224 2636 19306
rect 2608 19196 2728 19224
rect 2516 19094 2636 19122
rect 2502 19000 2558 19009
rect 2502 18935 2558 18944
rect 2516 9178 2544 18935
rect 2608 10810 2636 19094
rect 2700 15162 2728 19196
rect 2792 17105 2820 19382
rect 2976 19310 3004 22066
rect 3068 21010 3096 26862
rect 3148 26784 3200 26790
rect 3148 26726 3200 26732
rect 3056 21004 3108 21010
rect 3056 20946 3108 20952
rect 3056 20392 3108 20398
rect 3056 20334 3108 20340
rect 3068 19514 3096 20334
rect 3056 19508 3108 19514
rect 3056 19450 3108 19456
rect 3160 19446 3188 26726
rect 3148 19440 3200 19446
rect 3148 19382 3200 19388
rect 2964 19304 3016 19310
rect 2870 19272 2926 19281
rect 2964 19246 3016 19252
rect 2870 19207 2926 19216
rect 2884 17270 2912 19207
rect 2976 18902 3004 19246
rect 2964 18896 3016 18902
rect 2964 18838 3016 18844
rect 3252 18834 3280 27406
rect 3436 26625 3464 28018
rect 3884 27396 3936 27402
rect 3884 27338 3936 27344
rect 3700 27328 3752 27334
rect 3700 27270 3752 27276
rect 3422 26616 3478 26625
rect 3422 26551 3478 26560
rect 3332 25696 3384 25702
rect 3332 25638 3384 25644
rect 3344 20534 3372 25638
rect 3608 25288 3660 25294
rect 3608 25230 3660 25236
rect 3424 24608 3476 24614
rect 3424 24550 3476 24556
rect 3436 23497 3464 24550
rect 3516 24200 3568 24206
rect 3516 24142 3568 24148
rect 3422 23488 3478 23497
rect 3422 23423 3478 23432
rect 3528 23202 3556 24142
rect 3620 23730 3648 25230
rect 3608 23724 3660 23730
rect 3608 23666 3660 23672
rect 3620 23497 3648 23666
rect 3606 23488 3662 23497
rect 3606 23423 3662 23432
rect 3436 23174 3556 23202
rect 3332 20528 3384 20534
rect 3332 20470 3384 20476
rect 3332 20392 3384 20398
rect 3330 20360 3332 20369
rect 3384 20360 3386 20369
rect 3330 20295 3386 20304
rect 3240 18828 3292 18834
rect 3240 18770 3292 18776
rect 3054 18456 3110 18465
rect 3054 18391 3110 18400
rect 2964 18148 3016 18154
rect 2964 18090 3016 18096
rect 2872 17264 2924 17270
rect 2872 17206 2924 17212
rect 2778 17096 2834 17105
rect 2778 17031 2834 17040
rect 2870 16416 2926 16425
rect 2870 16351 2926 16360
rect 2884 16046 2912 16351
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2778 15736 2834 15745
rect 2778 15671 2834 15680
rect 2688 15156 2740 15162
rect 2688 15098 2740 15104
rect 2792 14074 2820 15671
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2884 13938 2912 14418
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2778 13696 2834 13705
rect 2778 13631 2834 13640
rect 2792 12102 2820 13631
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2778 11656 2834 11665
rect 2778 11591 2834 11600
rect 2596 10804 2648 10810
rect 2596 10746 2648 10752
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2608 10266 2636 10610
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2792 8974 2820 11591
rect 2884 10198 2912 12854
rect 2976 11234 3004 18090
rect 3068 11336 3096 18391
rect 3344 18222 3372 20295
rect 3332 18216 3384 18222
rect 3332 18158 3384 18164
rect 3240 16788 3292 16794
rect 3240 16730 3292 16736
rect 3146 16688 3202 16697
rect 3146 16623 3202 16632
rect 3160 12594 3188 16623
rect 3252 12714 3280 16730
rect 3436 16658 3464 23174
rect 3516 23112 3568 23118
rect 3516 23054 3568 23060
rect 3424 16652 3476 16658
rect 3424 16594 3476 16600
rect 3330 16008 3386 16017
rect 3330 15943 3386 15952
rect 3344 15910 3372 15943
rect 3332 15904 3384 15910
rect 3332 15846 3384 15852
rect 3344 15162 3372 15846
rect 3332 15156 3384 15162
rect 3332 15098 3384 15104
rect 3436 14618 3464 16594
rect 3528 16289 3556 23054
rect 3608 23044 3660 23050
rect 3608 22986 3660 22992
rect 3620 22574 3648 22986
rect 3608 22568 3660 22574
rect 3608 22510 3660 22516
rect 3620 22234 3648 22510
rect 3608 22228 3660 22234
rect 3608 22170 3660 22176
rect 3608 21956 3660 21962
rect 3608 21898 3660 21904
rect 3620 21486 3648 21898
rect 3608 21480 3660 21486
rect 3608 21422 3660 21428
rect 3620 21078 3648 21422
rect 3608 21072 3660 21078
rect 3608 21014 3660 21020
rect 3620 19922 3648 21014
rect 3712 20602 3740 27270
rect 3792 25696 3844 25702
rect 3792 25638 3844 25644
rect 3700 20596 3752 20602
rect 3700 20538 3752 20544
rect 3698 20496 3754 20505
rect 3698 20431 3754 20440
rect 3712 20262 3740 20431
rect 3700 20256 3752 20262
rect 3700 20198 3752 20204
rect 3608 19916 3660 19922
rect 3608 19858 3660 19864
rect 3608 19780 3660 19786
rect 3608 19722 3660 19728
rect 3514 16280 3570 16289
rect 3514 16215 3570 16224
rect 3528 15638 3556 16215
rect 3620 15994 3648 19722
rect 3698 19408 3754 19417
rect 3698 19343 3754 19352
rect 3712 17338 3740 19343
rect 3700 17332 3752 17338
rect 3700 17274 3752 17280
rect 3712 16096 3740 17274
rect 3804 16522 3832 25638
rect 3896 24993 3924 27338
rect 4080 27305 4108 28018
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4066 27296 4122 27305
rect 4066 27231 4122 27240
rect 4620 26784 4672 26790
rect 4620 26726 4672 26732
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4632 26353 4660 26726
rect 4618 26344 4674 26353
rect 4618 26279 4674 26288
rect 3976 25900 4028 25906
rect 3976 25842 4028 25848
rect 3882 24984 3938 24993
rect 3882 24919 3938 24928
rect 3884 24812 3936 24818
rect 3884 24754 3936 24760
rect 3896 24188 3924 24754
rect 3988 24342 4016 25842
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 3976 24336 4028 24342
rect 3976 24278 4028 24284
rect 3976 24200 4028 24206
rect 3896 24168 3976 24188
rect 4028 24168 4030 24177
rect 3896 24160 3974 24168
rect 4724 24154 4752 29446
rect 4804 25900 4856 25906
rect 4804 25842 4856 25848
rect 4816 24954 4844 25842
rect 4896 25152 4948 25158
rect 4896 25094 4948 25100
rect 4804 24948 4856 24954
rect 4804 24890 4856 24896
rect 4816 24857 4844 24890
rect 4802 24848 4858 24857
rect 4802 24783 4858 24792
rect 4804 24200 4856 24206
rect 3974 24103 4030 24112
rect 4632 24126 4752 24154
rect 4802 24168 4804 24177
rect 4856 24168 4858 24177
rect 3882 23896 3938 23905
rect 3882 23831 3884 23840
rect 3936 23831 3938 23840
rect 3884 23802 3936 23808
rect 3884 23520 3936 23526
rect 3884 23462 3936 23468
rect 3896 21146 3924 23462
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23118 4660 24126
rect 4802 24103 4858 24112
rect 4712 23724 4764 23730
rect 4712 23666 4764 23672
rect 4724 23633 4752 23666
rect 4710 23624 4766 23633
rect 4710 23559 4766 23568
rect 4712 23520 4764 23526
rect 4712 23462 4764 23468
rect 4620 23112 4672 23118
rect 4620 23054 4672 23060
rect 3976 23044 4028 23050
rect 3976 22986 4028 22992
rect 3884 21140 3936 21146
rect 3884 21082 3936 21088
rect 3988 20806 4016 22986
rect 4068 22976 4120 22982
rect 4068 22918 4120 22924
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 3976 20800 4028 20806
rect 3976 20742 4028 20748
rect 3988 20505 4016 20742
rect 3974 20496 4030 20505
rect 3974 20431 4030 20440
rect 4080 20346 4108 22918
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4632 22098 4660 22918
rect 4620 22092 4672 22098
rect 4620 22034 4672 22040
rect 4160 22024 4212 22030
rect 4160 21966 4212 21972
rect 4172 21622 4200 21966
rect 4252 21888 4304 21894
rect 4252 21830 4304 21836
rect 4344 21888 4396 21894
rect 4344 21830 4396 21836
rect 4160 21616 4212 21622
rect 4160 21558 4212 21564
rect 4264 21418 4292 21830
rect 4356 21729 4384 21830
rect 4342 21720 4398 21729
rect 4342 21655 4398 21664
rect 4252 21412 4304 21418
rect 4252 21354 4304 21360
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4158 21040 4214 21049
rect 4724 21010 4752 23462
rect 4804 22024 4856 22030
rect 4804 21966 4856 21972
rect 4816 21486 4844 21966
rect 4804 21480 4856 21486
rect 4804 21422 4856 21428
rect 4804 21344 4856 21350
rect 4804 21286 4856 21292
rect 4158 20975 4214 20984
rect 4252 21004 4304 21010
rect 4172 20466 4200 20975
rect 4252 20946 4304 20952
rect 4712 21004 4764 21010
rect 4712 20946 4764 20952
rect 4264 20874 4292 20946
rect 4816 20874 4844 21286
rect 4252 20868 4304 20874
rect 4252 20810 4304 20816
rect 4804 20868 4856 20874
rect 4804 20810 4856 20816
rect 4710 20768 4766 20777
rect 4710 20703 4766 20712
rect 4160 20460 4212 20466
rect 4160 20402 4212 20408
rect 3896 20318 4108 20346
rect 3896 19310 3924 20318
rect 4172 20244 4200 20402
rect 4080 20216 4200 20244
rect 4080 20058 4108 20216
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3976 20052 4028 20058
rect 3976 19994 4028 20000
rect 4068 20052 4120 20058
rect 4068 19994 4120 20000
rect 4528 20052 4580 20058
rect 4528 19994 4580 20000
rect 3884 19304 3936 19310
rect 3884 19246 3936 19252
rect 3988 19242 4016 19994
rect 4160 19916 4212 19922
rect 4160 19858 4212 19864
rect 4172 19802 4200 19858
rect 4080 19786 4200 19802
rect 4068 19780 4200 19786
rect 4120 19774 4200 19780
rect 4068 19722 4120 19728
rect 4540 19281 4568 19994
rect 4618 19952 4674 19961
rect 4618 19887 4674 19896
rect 4526 19272 4582 19281
rect 3976 19236 4028 19242
rect 4526 19207 4582 19216
rect 3976 19178 4028 19184
rect 3988 18358 4016 19178
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 3976 18352 4028 18358
rect 3976 18294 4028 18300
rect 4080 18222 4108 19110
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4250 18864 4306 18873
rect 4250 18799 4306 18808
rect 4264 18766 4292 18799
rect 4252 18760 4304 18766
rect 4252 18702 4304 18708
rect 4160 18692 4212 18698
rect 4160 18634 4212 18640
rect 4068 18216 4120 18222
rect 4068 18158 4120 18164
rect 4172 18086 4200 18634
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17882 4660 19887
rect 4724 18426 4752 20703
rect 4816 20641 4844 20810
rect 4802 20632 4858 20641
rect 4802 20567 4858 20576
rect 4816 20534 4844 20567
rect 4804 20528 4856 20534
rect 4804 20470 4856 20476
rect 4802 20224 4858 20233
rect 4802 20159 4858 20168
rect 4712 18420 4764 18426
rect 4712 18362 4764 18368
rect 4816 18086 4844 20159
rect 4908 19786 4936 25094
rect 5000 22098 5028 29990
rect 5080 27872 5132 27878
rect 5080 27814 5132 27820
rect 5092 22642 5120 27814
rect 5184 27130 5212 30126
rect 5172 27124 5224 27130
rect 5172 27066 5224 27072
rect 5264 26920 5316 26926
rect 5264 26862 5316 26868
rect 5172 26376 5224 26382
rect 5172 26318 5224 26324
rect 5184 24993 5212 26318
rect 5170 24984 5226 24993
rect 5170 24919 5226 24928
rect 5170 24848 5226 24857
rect 5170 24783 5226 24792
rect 5184 23730 5212 24783
rect 5172 23724 5224 23730
rect 5172 23666 5224 23672
rect 5276 23610 5304 26862
rect 5184 23582 5304 23610
rect 5080 22636 5132 22642
rect 5080 22578 5132 22584
rect 5184 22522 5212 23582
rect 5264 23520 5316 23526
rect 5264 23462 5316 23468
rect 5276 22545 5304 23462
rect 5092 22494 5212 22522
rect 5262 22536 5318 22545
rect 4988 22092 5040 22098
rect 4988 22034 5040 22040
rect 4986 21992 5042 22001
rect 4986 21927 5042 21936
rect 4896 19780 4948 19786
rect 4896 19722 4948 19728
rect 4894 19680 4950 19689
rect 4894 19615 4950 19624
rect 4908 19378 4936 19615
rect 4896 19372 4948 19378
rect 4896 19314 4948 19320
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 3974 17640 4030 17649
rect 3974 17575 4030 17584
rect 4250 17640 4306 17649
rect 4250 17575 4252 17584
rect 3988 17066 4016 17575
rect 4304 17575 4306 17584
rect 4526 17640 4582 17649
rect 4526 17575 4582 17584
rect 4252 17546 4304 17552
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 4080 17134 4108 17478
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 4540 17082 4568 17575
rect 4632 17270 4660 17818
rect 4710 17776 4766 17785
rect 4710 17711 4766 17720
rect 4724 17610 4752 17711
rect 4712 17604 4764 17610
rect 4712 17546 4764 17552
rect 4908 17490 4936 19314
rect 5000 17882 5028 21927
rect 5092 21865 5120 22494
rect 5262 22471 5318 22480
rect 5172 22432 5224 22438
rect 5172 22374 5224 22380
rect 5078 21856 5134 21865
rect 5078 21791 5134 21800
rect 5080 21412 5132 21418
rect 5080 21354 5132 21360
rect 5092 20233 5120 21354
rect 5184 20534 5212 22374
rect 5368 22094 5396 30534
rect 5736 29306 5764 34546
rect 5828 30734 5856 36518
rect 6380 30734 6408 37062
rect 6564 32910 6592 37062
rect 6552 32904 6604 32910
rect 6552 32846 6604 32852
rect 5816 30728 5868 30734
rect 5816 30670 5868 30676
rect 6368 30728 6420 30734
rect 6368 30670 6420 30676
rect 6552 30592 6604 30598
rect 6552 30534 6604 30540
rect 5816 29640 5868 29646
rect 5816 29582 5868 29588
rect 5724 29300 5776 29306
rect 5724 29242 5776 29248
rect 5828 28218 5856 29582
rect 5816 28212 5868 28218
rect 5816 28154 5868 28160
rect 6460 28076 6512 28082
rect 6460 28018 6512 28024
rect 5448 26376 5500 26382
rect 5448 26318 5500 26324
rect 6092 26376 6144 26382
rect 6092 26318 6144 26324
rect 5276 22066 5396 22094
rect 5276 21010 5304 22066
rect 5264 21004 5316 21010
rect 5264 20946 5316 20952
rect 5356 20868 5408 20874
rect 5356 20810 5408 20816
rect 5172 20528 5224 20534
rect 5172 20470 5224 20476
rect 5078 20224 5134 20233
rect 5078 20159 5134 20168
rect 5368 20097 5396 20810
rect 5354 20088 5410 20097
rect 5354 20023 5410 20032
rect 5080 19780 5132 19786
rect 5080 19722 5132 19728
rect 5356 19780 5408 19786
rect 5356 19722 5408 19728
rect 5092 19553 5120 19722
rect 5264 19712 5316 19718
rect 5170 19680 5226 19689
rect 5264 19654 5316 19660
rect 5170 19615 5226 19624
rect 5078 19544 5134 19553
rect 5078 19479 5134 19488
rect 5184 19446 5212 19615
rect 5172 19440 5224 19446
rect 5172 19382 5224 19388
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 5092 18698 5120 19246
rect 5184 18834 5212 19382
rect 5172 18828 5224 18834
rect 5172 18770 5224 18776
rect 5080 18692 5132 18698
rect 5080 18634 5132 18640
rect 5276 18426 5304 19654
rect 5368 19310 5396 19722
rect 5460 19446 5488 26318
rect 6000 25968 6052 25974
rect 6000 25910 6052 25916
rect 5632 25900 5684 25906
rect 5632 25842 5684 25848
rect 5644 25294 5672 25842
rect 5724 25832 5776 25838
rect 5724 25774 5776 25780
rect 5632 25288 5684 25294
rect 5632 25230 5684 25236
rect 5540 24812 5592 24818
rect 5540 24754 5592 24760
rect 5448 19440 5500 19446
rect 5448 19382 5500 19388
rect 5356 19304 5408 19310
rect 5356 19246 5408 19252
rect 5368 18970 5396 19246
rect 5356 18964 5408 18970
rect 5356 18906 5408 18912
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5264 18420 5316 18426
rect 5264 18362 5316 18368
rect 5172 18352 5224 18358
rect 5172 18294 5224 18300
rect 5080 18284 5132 18290
rect 5080 18226 5132 18232
rect 4988 17876 5040 17882
rect 4988 17818 5040 17824
rect 4724 17462 4936 17490
rect 4620 17264 4672 17270
rect 4620 17206 4672 17212
rect 3976 17060 4028 17066
rect 3976 17002 4028 17008
rect 3988 16794 4016 17002
rect 3976 16788 4028 16794
rect 3976 16730 4028 16736
rect 4080 16640 4108 17070
rect 4540 17054 4660 17082
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4252 16652 4304 16658
rect 4080 16612 4252 16640
rect 4252 16594 4304 16600
rect 3792 16516 3844 16522
rect 3792 16458 3844 16464
rect 4068 16448 4120 16454
rect 4066 16416 4068 16425
rect 4120 16416 4122 16425
rect 4066 16351 4122 16360
rect 4264 16114 4292 16594
rect 4528 16584 4580 16590
rect 4528 16526 4580 16532
rect 4252 16108 4304 16114
rect 3712 16068 3832 16096
rect 3620 15966 3740 15994
rect 3608 15904 3660 15910
rect 3608 15846 3660 15852
rect 3620 15706 3648 15846
rect 3608 15700 3660 15706
rect 3608 15642 3660 15648
rect 3516 15632 3568 15638
rect 3516 15574 3568 15580
rect 3514 15056 3570 15065
rect 3514 14991 3570 15000
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 3528 14346 3556 14991
rect 3516 14340 3568 14346
rect 3516 14282 3568 14288
rect 3516 13388 3568 13394
rect 3516 13330 3568 13336
rect 3424 12912 3476 12918
rect 3424 12854 3476 12860
rect 3240 12708 3292 12714
rect 3240 12650 3292 12656
rect 3160 12566 3280 12594
rect 3252 12374 3280 12566
rect 3436 12434 3464 12854
rect 3528 12782 3556 13330
rect 3516 12776 3568 12782
rect 3516 12718 3568 12724
rect 3344 12406 3464 12434
rect 3516 12436 3568 12442
rect 3240 12368 3292 12374
rect 3146 12336 3202 12345
rect 3240 12310 3292 12316
rect 3146 12271 3202 12280
rect 3160 12170 3188 12271
rect 3148 12164 3200 12170
rect 3148 12106 3200 12112
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 3068 11308 3188 11336
rect 2976 11206 3096 11234
rect 3068 10810 3096 11206
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 2872 10192 2924 10198
rect 2872 10134 2924 10140
rect 3160 10062 3188 11308
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 3252 8838 3280 12038
rect 3344 9178 3372 12406
rect 3516 12378 3568 12384
rect 3422 11656 3478 11665
rect 3422 11591 3478 11600
rect 3436 11354 3464 11591
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3422 9480 3478 9489
rect 3422 9415 3478 9424
rect 3436 9382 3464 9415
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 2792 8566 2820 8774
rect 2780 8560 2832 8566
rect 2780 8502 2832 8508
rect 3436 8242 3464 9318
rect 3528 8974 3556 12378
rect 3620 10742 3648 15642
rect 3712 13841 3740 15966
rect 3804 15570 3832 16068
rect 4080 16068 4252 16096
rect 3974 15600 4030 15609
rect 3792 15564 3844 15570
rect 4080 15570 4108 16068
rect 4252 16050 4304 16056
rect 4540 16028 4568 16526
rect 4632 16522 4660 17054
rect 4620 16516 4672 16522
rect 4620 16458 4672 16464
rect 4620 16176 4672 16182
rect 4724 16164 4752 17462
rect 4802 17368 4858 17377
rect 4802 17303 4858 17312
rect 4672 16136 4752 16164
rect 4620 16118 4672 16124
rect 4540 16000 4660 16028
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 3974 15535 4030 15544
rect 4068 15564 4120 15570
rect 3792 15506 3844 15512
rect 3988 15502 4016 15535
rect 4068 15506 4120 15512
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 4066 15328 4122 15337
rect 4066 15263 4122 15272
rect 4080 15094 4108 15263
rect 4068 15088 4120 15094
rect 3896 15048 4068 15076
rect 3792 14952 3844 14958
rect 3792 14894 3844 14900
rect 3804 14482 3832 14894
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 3698 13832 3754 13841
rect 3698 13767 3754 13776
rect 3700 13524 3752 13530
rect 3700 13466 3752 13472
rect 3712 12782 3740 13466
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 3700 12776 3752 12782
rect 3700 12718 3752 12724
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 3712 12209 3740 12378
rect 3804 12306 3832 13262
rect 3792 12300 3844 12306
rect 3792 12242 3844 12248
rect 3698 12200 3754 12209
rect 3698 12135 3754 12144
rect 3804 11898 3832 12242
rect 3792 11892 3844 11898
rect 3792 11834 3844 11840
rect 3608 10736 3660 10742
rect 3608 10678 3660 10684
rect 3804 10674 3832 11834
rect 3896 11642 3924 15048
rect 4068 15030 4120 15036
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4632 14550 4660 16000
rect 4724 14793 4752 16136
rect 4816 15570 4844 17303
rect 5000 16794 5028 17818
rect 4988 16788 5040 16794
rect 4988 16730 5040 16736
rect 5092 16454 5120 18226
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 4988 16040 5040 16046
rect 4988 15982 5040 15988
rect 4804 15564 4856 15570
rect 4804 15506 4856 15512
rect 4710 14784 4766 14793
rect 4710 14719 4766 14728
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4620 14544 4672 14550
rect 4620 14486 4672 14492
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 3974 13968 4030 13977
rect 3974 13903 4030 13912
rect 3988 13462 4016 13903
rect 3976 13456 4028 13462
rect 3976 13398 4028 13404
rect 3974 13288 4030 13297
rect 3974 13223 3976 13232
rect 4028 13223 4030 13232
rect 3976 13194 4028 13200
rect 3974 12744 4030 12753
rect 3974 12679 4030 12688
rect 3988 12374 4016 12679
rect 3976 12368 4028 12374
rect 3976 12310 4028 12316
rect 4080 12170 4108 14350
rect 4618 14104 4674 14113
rect 4618 14039 4620 14048
rect 4672 14039 4674 14048
rect 4620 14010 4672 14016
rect 4712 14000 4764 14006
rect 4712 13942 4764 13948
rect 4816 13954 4844 14554
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4342 13424 4398 13433
rect 4342 13359 4398 13368
rect 4356 13258 4384 13359
rect 4344 13252 4396 13258
rect 4344 13194 4396 13200
rect 4252 12776 4304 12782
rect 4250 12744 4252 12753
rect 4304 12744 4306 12753
rect 4250 12679 4306 12688
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 12238 4660 12582
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4068 12164 4120 12170
rect 4068 12106 4120 12112
rect 3896 11614 4016 11642
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3700 10600 3752 10606
rect 3988 10554 4016 11614
rect 3752 10548 4016 10554
rect 3700 10542 4016 10548
rect 3712 10526 4016 10542
rect 3790 10296 3846 10305
rect 3790 10231 3846 10240
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3516 8968 3568 8974
rect 3516 8910 3568 8916
rect 3528 8650 3556 8910
rect 3712 8906 3740 9998
rect 3804 9722 3832 10231
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3884 9648 3936 9654
rect 3884 9590 3936 9596
rect 3700 8900 3752 8906
rect 3700 8842 3752 8848
rect 3528 8622 3648 8650
rect 3516 8560 3568 8566
rect 3516 8502 3568 8508
rect 1820 6896 1822 6905
rect 1766 6831 1822 6840
rect 2056 6886 2176 6914
rect 2332 6886 2452 6914
rect 3160 8214 3464 8242
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 1596 5914 1624 6734
rect 1964 6458 1992 6734
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1596 4690 1624 5646
rect 1584 4684 1636 4690
rect 1584 4626 1636 4632
rect 1676 4208 1728 4214
rect 1674 4176 1676 4185
rect 1728 4176 1730 4185
rect 2056 4146 2084 6886
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 1674 4111 1730 4120
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 1492 2644 1544 2650
rect 1492 2586 1544 2592
rect 1676 2372 1728 2378
rect 1676 2314 1728 2320
rect 18 200 74 800
rect 662 200 718 800
rect 1688 785 1716 2314
rect 1964 800 1992 3062
rect 2240 2446 2268 6598
rect 2332 6322 2360 6886
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2504 6112 2556 6118
rect 2504 6054 2556 6060
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 2516 3058 2544 6054
rect 2872 5636 2924 5642
rect 2872 5578 2924 5584
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 2688 2848 2740 2854
rect 2688 2790 2740 2796
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 2516 2145 2544 2246
rect 2502 2136 2558 2145
rect 2502 2071 2558 2080
rect 2700 2009 2728 2790
rect 2686 2000 2742 2009
rect 2686 1935 2742 1944
rect 2884 1873 2912 5578
rect 3068 2446 3096 6054
rect 3160 4826 3188 8214
rect 3422 8120 3478 8129
rect 3422 8055 3424 8064
rect 3476 8055 3478 8064
rect 3424 8026 3476 8032
rect 3436 7342 3464 8026
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3148 3392 3200 3398
rect 3146 3360 3148 3369
rect 3200 3360 3202 3369
rect 3146 3295 3202 3304
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 2870 1864 2926 1873
rect 2870 1799 2926 1808
rect 3252 800 3280 6734
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 3344 4690 3372 5034
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3344 4146 3372 4626
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3436 3194 3464 6258
rect 3528 5370 3556 8502
rect 3620 6798 3648 8622
rect 3896 6866 3924 9590
rect 3988 9518 4016 9998
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 4080 8974 4108 12106
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 4172 11694 4200 12038
rect 4632 11830 4660 12174
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 11218 4660 11766
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4618 11112 4674 11121
rect 4618 11047 4674 11056
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 4160 9920 4212 9926
rect 4540 9897 4568 9930
rect 4160 9862 4212 9868
rect 4526 9888 4582 9897
rect 4172 9586 4200 9862
rect 4526 9823 4582 9832
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4068 8968 4120 8974
rect 3974 8936 4030 8945
rect 4068 8910 4120 8916
rect 3974 8871 4030 8880
rect 3988 8566 4016 8871
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3988 7954 4016 8230
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3976 7948 4028 7954
rect 3976 7890 4028 7896
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 3608 6792 3660 6798
rect 3608 6734 3660 6740
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3620 5234 3648 6734
rect 3792 5636 3844 5642
rect 3792 5578 3844 5584
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3620 4622 3648 5170
rect 3700 4752 3752 4758
rect 3700 4694 3752 4700
rect 3608 4616 3660 4622
rect 3608 4558 3660 4564
rect 3516 4480 3568 4486
rect 3516 4422 3568 4428
rect 3528 4214 3556 4422
rect 3516 4208 3568 4214
rect 3516 4150 3568 4156
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 3712 3058 3740 4694
rect 3804 3126 3832 5578
rect 3988 4826 4016 7754
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 4172 7410 4200 7686
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4068 5840 4120 5846
rect 4066 5808 4068 5817
rect 4120 5808 4122 5817
rect 4066 5743 4122 5752
rect 4632 5370 4660 11047
rect 4724 10266 4752 13942
rect 4816 13926 4936 13954
rect 4804 13252 4856 13258
rect 4804 13194 4856 13200
rect 4816 12986 4844 13194
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4724 9042 4752 9318
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4816 8498 4844 11834
rect 4908 11257 4936 13926
rect 5000 12481 5028 15982
rect 5092 14414 5120 16390
rect 5184 16153 5212 18294
rect 5262 18184 5318 18193
rect 5262 18119 5318 18128
rect 5170 16144 5226 16153
rect 5170 16079 5226 16088
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 5184 14618 5212 15982
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 5080 14408 5132 14414
rect 5080 14350 5132 14356
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5078 14240 5134 14249
rect 5078 14175 5134 14184
rect 5092 13938 5120 14175
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 5184 13138 5212 14350
rect 5276 14278 5304 18119
rect 5460 15609 5488 18906
rect 5552 17270 5580 24754
rect 5632 24132 5684 24138
rect 5632 24074 5684 24080
rect 5540 17264 5592 17270
rect 5540 17206 5592 17212
rect 5644 16522 5672 24074
rect 5736 21894 5764 25774
rect 5816 24064 5868 24070
rect 5816 24006 5868 24012
rect 5828 23594 5856 24006
rect 5816 23588 5868 23594
rect 5816 23530 5868 23536
rect 5816 22432 5868 22438
rect 5816 22374 5868 22380
rect 5828 22098 5856 22374
rect 5816 22092 5868 22098
rect 5816 22034 5868 22040
rect 5816 21956 5868 21962
rect 5816 21898 5868 21904
rect 5724 21888 5776 21894
rect 5724 21830 5776 21836
rect 5828 21350 5856 21898
rect 5816 21344 5868 21350
rect 5816 21286 5868 21292
rect 5724 21072 5776 21078
rect 5724 21014 5776 21020
rect 5736 19854 5764 21014
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 5724 19304 5776 19310
rect 5828 19292 5856 21286
rect 6012 20618 6040 25910
rect 6104 24188 6132 26318
rect 6184 25696 6236 25702
rect 6184 25638 6236 25644
rect 6276 25696 6328 25702
rect 6276 25638 6328 25644
rect 6196 25362 6224 25638
rect 6184 25356 6236 25362
rect 6184 25298 6236 25304
rect 6288 25294 6316 25638
rect 6276 25288 6328 25294
rect 6276 25230 6328 25236
rect 6368 25288 6420 25294
rect 6368 25230 6420 25236
rect 6104 24160 6224 24188
rect 6092 23792 6144 23798
rect 6092 23734 6144 23740
rect 6104 20806 6132 23734
rect 6092 20800 6144 20806
rect 6092 20742 6144 20748
rect 6012 20590 6132 20618
rect 6000 20528 6052 20534
rect 6000 20470 6052 20476
rect 5906 20224 5962 20233
rect 5906 20159 5962 20168
rect 5776 19264 5856 19292
rect 5724 19246 5776 19252
rect 5736 18222 5764 19246
rect 5724 18216 5776 18222
rect 5724 18158 5776 18164
rect 5632 16516 5684 16522
rect 5632 16458 5684 16464
rect 5538 16280 5594 16289
rect 5538 16215 5540 16224
rect 5592 16215 5594 16224
rect 5540 16186 5592 16192
rect 5814 16144 5870 16153
rect 5814 16079 5870 16088
rect 5632 15632 5684 15638
rect 5446 15600 5502 15609
rect 5632 15574 5684 15580
rect 5446 15535 5502 15544
rect 5538 15192 5594 15201
rect 5538 15127 5540 15136
rect 5592 15127 5594 15136
rect 5540 15098 5592 15104
rect 5538 14648 5594 14657
rect 5538 14583 5540 14592
rect 5592 14583 5594 14592
rect 5540 14554 5592 14560
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5644 13954 5672 15574
rect 5828 14074 5856 16079
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5920 13954 5948 20159
rect 6012 19446 6040 20470
rect 6000 19440 6052 19446
rect 6000 19382 6052 19388
rect 6012 18834 6040 19382
rect 6000 18828 6052 18834
rect 6000 18770 6052 18776
rect 6000 17604 6052 17610
rect 6000 17546 6052 17552
rect 6012 16046 6040 17546
rect 6104 16250 6132 20590
rect 6196 20330 6224 24160
rect 6288 23322 6316 25230
rect 6276 23316 6328 23322
rect 6276 23258 6328 23264
rect 6276 22500 6328 22506
rect 6276 22442 6328 22448
rect 6184 20324 6236 20330
rect 6184 20266 6236 20272
rect 6184 19848 6236 19854
rect 6184 19790 6236 19796
rect 6196 17513 6224 19790
rect 6182 17504 6238 17513
rect 6182 17439 6238 17448
rect 6092 16244 6144 16250
rect 6092 16186 6144 16192
rect 6000 16040 6052 16046
rect 6000 15982 6052 15988
rect 6196 15858 6224 17439
rect 6288 16998 6316 22442
rect 6380 22001 6408 25230
rect 6472 24732 6500 28018
rect 6564 27538 6592 30534
rect 6840 29646 6868 37130
rect 7760 37126 7788 39200
rect 7840 37256 7892 37262
rect 7840 37198 7892 37204
rect 7748 37120 7800 37126
rect 7748 37062 7800 37068
rect 7852 36854 7880 37198
rect 9048 36922 9076 39200
rect 9496 37188 9548 37194
rect 9496 37130 9548 37136
rect 9036 36916 9088 36922
rect 9036 36858 9088 36864
rect 7840 36848 7892 36854
rect 7840 36790 7892 36796
rect 9128 36780 9180 36786
rect 9128 36722 9180 36728
rect 7472 35624 7524 35630
rect 7472 35566 7524 35572
rect 6828 29640 6880 29646
rect 6828 29582 6880 29588
rect 6552 27532 6604 27538
rect 6552 27474 6604 27480
rect 6564 24857 6592 27474
rect 6828 26988 6880 26994
rect 6828 26930 6880 26936
rect 6840 26042 6868 26930
rect 7288 26784 7340 26790
rect 7288 26726 7340 26732
rect 6920 26376 6972 26382
rect 6920 26318 6972 26324
rect 6828 26036 6880 26042
rect 6828 25978 6880 25984
rect 6932 25906 6960 26318
rect 6920 25900 6972 25906
rect 6920 25842 6972 25848
rect 7012 25764 7064 25770
rect 7012 25706 7064 25712
rect 6736 25152 6788 25158
rect 6736 25094 6788 25100
rect 6550 24848 6606 24857
rect 6550 24783 6606 24792
rect 6472 24704 6592 24732
rect 6460 24404 6512 24410
rect 6460 24346 6512 24352
rect 6472 23730 6500 24346
rect 6460 23724 6512 23730
rect 6460 23666 6512 23672
rect 6564 23610 6592 24704
rect 6644 24132 6696 24138
rect 6644 24074 6696 24080
rect 6656 23866 6684 24074
rect 6644 23860 6696 23866
rect 6644 23802 6696 23808
rect 6472 23582 6592 23610
rect 6472 22710 6500 23582
rect 6644 23520 6696 23526
rect 6644 23462 6696 23468
rect 6656 23186 6684 23462
rect 6644 23180 6696 23186
rect 6644 23122 6696 23128
rect 6552 23112 6604 23118
rect 6552 23054 6604 23060
rect 6460 22704 6512 22710
rect 6460 22646 6512 22652
rect 6472 22506 6500 22646
rect 6460 22500 6512 22506
rect 6460 22442 6512 22448
rect 6460 22092 6512 22098
rect 6564 22094 6592 23054
rect 6748 22778 6776 25094
rect 7024 24993 7052 25706
rect 7196 25492 7248 25498
rect 7196 25434 7248 25440
rect 7208 25129 7236 25434
rect 7194 25120 7250 25129
rect 7194 25055 7250 25064
rect 7010 24984 7066 24993
rect 7010 24919 7066 24928
rect 6828 24744 6880 24750
rect 6828 24686 6880 24692
rect 7012 24744 7064 24750
rect 7012 24686 7064 24692
rect 6840 24342 6868 24686
rect 6828 24336 6880 24342
rect 6828 24278 6880 24284
rect 7024 24274 7052 24686
rect 7012 24268 7064 24274
rect 7012 24210 7064 24216
rect 6828 24200 6880 24206
rect 6828 24142 6880 24148
rect 6840 23866 6868 24142
rect 7196 24132 7248 24138
rect 7116 24092 7196 24120
rect 6828 23860 6880 23866
rect 6828 23802 6880 23808
rect 7012 23792 7064 23798
rect 7012 23734 7064 23740
rect 7024 23118 7052 23734
rect 7012 23112 7064 23118
rect 7012 23054 7064 23060
rect 6736 22772 6788 22778
rect 6736 22714 6788 22720
rect 6736 22636 6788 22642
rect 6736 22578 6788 22584
rect 6644 22432 6696 22438
rect 6748 22409 6776 22578
rect 6644 22374 6696 22380
rect 6734 22400 6790 22409
rect 6656 22250 6684 22374
rect 6734 22335 6790 22344
rect 6656 22222 6776 22250
rect 6564 22066 6684 22094
rect 6460 22034 6512 22040
rect 6366 21992 6422 22001
rect 6366 21927 6422 21936
rect 6366 21584 6422 21593
rect 6366 21519 6368 21528
rect 6420 21519 6422 21528
rect 6368 21490 6420 21496
rect 6472 21486 6500 22034
rect 6460 21480 6512 21486
rect 6460 21422 6512 21428
rect 6368 20800 6420 20806
rect 6368 20742 6420 20748
rect 6380 18766 6408 20742
rect 6458 20496 6514 20505
rect 6458 20431 6514 20440
rect 6472 19786 6500 20431
rect 6460 19780 6512 19786
rect 6460 19722 6512 19728
rect 6460 19440 6512 19446
rect 6656 19417 6684 22066
rect 6748 21622 6776 22222
rect 6736 21616 6788 21622
rect 6736 21558 6788 21564
rect 6828 21480 6880 21486
rect 6828 21422 6880 21428
rect 6840 21078 6868 21422
rect 6828 21072 6880 21078
rect 6828 21014 6880 21020
rect 6828 20936 6880 20942
rect 6828 20878 6880 20884
rect 6734 20224 6790 20233
rect 6734 20159 6790 20168
rect 6748 19922 6776 20159
rect 6840 19938 6868 20878
rect 7116 20602 7144 24092
rect 7196 24074 7248 24080
rect 7300 24018 7328 26726
rect 7380 24336 7432 24342
rect 7380 24278 7432 24284
rect 7208 23990 7328 24018
rect 7208 23050 7236 23990
rect 7288 23724 7340 23730
rect 7288 23666 7340 23672
rect 7196 23044 7248 23050
rect 7196 22986 7248 22992
rect 7208 21010 7236 22986
rect 7196 21004 7248 21010
rect 7196 20946 7248 20952
rect 7104 20596 7156 20602
rect 7104 20538 7156 20544
rect 7012 20528 7064 20534
rect 7012 20470 7064 20476
rect 6736 19916 6788 19922
rect 6840 19910 6960 19938
rect 6736 19858 6788 19864
rect 6826 19816 6882 19825
rect 6826 19751 6882 19760
rect 6460 19382 6512 19388
rect 6642 19408 6698 19417
rect 6368 18760 6420 18766
rect 6366 18728 6368 18737
rect 6420 18728 6422 18737
rect 6366 18663 6422 18672
rect 6276 16992 6328 16998
rect 6276 16934 6328 16940
rect 5552 13926 5672 13954
rect 5828 13926 5948 13954
rect 6012 15830 6224 15858
rect 5262 13696 5318 13705
rect 5262 13631 5318 13640
rect 5092 13110 5212 13138
rect 4986 12472 5042 12481
rect 4986 12407 5042 12416
rect 5092 12186 5120 13110
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5184 12442 5212 12582
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 5000 12158 5120 12186
rect 5000 12102 5028 12158
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 4894 11248 4950 11257
rect 4894 11183 4950 11192
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4908 8430 4936 11018
rect 5000 10282 5028 12038
rect 5276 10606 5304 13631
rect 5552 11694 5580 13926
rect 5632 13184 5684 13190
rect 5632 13126 5684 13132
rect 5644 12850 5672 13126
rect 5828 12866 5856 13926
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 5920 12986 5948 13806
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 5632 12844 5684 12850
rect 5828 12838 5948 12866
rect 5632 12786 5684 12792
rect 5630 12744 5686 12753
rect 5630 12679 5632 12688
rect 5684 12679 5686 12688
rect 5632 12650 5684 12656
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5356 11008 5408 11014
rect 5356 10950 5408 10956
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 5368 10452 5396 10950
rect 5552 10810 5580 11630
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5448 10736 5500 10742
rect 5446 10704 5448 10713
rect 5500 10704 5502 10713
rect 5446 10639 5502 10648
rect 5644 10588 5672 12650
rect 5816 11688 5868 11694
rect 5816 11630 5868 11636
rect 5184 10424 5396 10452
rect 5460 10560 5672 10588
rect 5000 10254 5120 10282
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4724 8294 4752 8366
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4724 7886 4752 8230
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 5000 6458 5028 9590
rect 5092 7546 5120 10254
rect 5184 9518 5212 10424
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5368 8566 5396 9658
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 5460 8362 5488 10560
rect 5828 10554 5856 11630
rect 5736 10526 5856 10554
rect 5538 9888 5594 9897
rect 5538 9823 5594 9832
rect 5552 9722 5580 9823
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4632 4214 4660 4422
rect 4620 4208 4672 4214
rect 4620 4150 4672 4156
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 3884 3664 3936 3670
rect 3884 3606 3936 3612
rect 3792 3120 3844 3126
rect 3792 3062 3844 3068
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3896 800 3924 3606
rect 3988 3058 4016 3878
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 4080 3505 4108 3538
rect 4632 3534 4660 3878
rect 4620 3528 4672 3534
rect 4066 3496 4122 3505
rect 4620 3470 4672 3476
rect 4066 3431 4122 3440
rect 4160 3460 4212 3466
rect 4160 3402 4212 3408
rect 4344 3460 4396 3466
rect 4344 3402 4396 3408
rect 4172 3126 4200 3402
rect 4160 3120 4212 3126
rect 4356 3097 4384 3402
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4160 3062 4212 3068
rect 4342 3088 4398 3097
rect 3976 3052 4028 3058
rect 4342 3023 4398 3032
rect 3976 2994 4028 3000
rect 4066 2952 4122 2961
rect 4066 2887 4068 2896
rect 4120 2887 4122 2896
rect 4068 2858 4120 2864
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2446 4660 3334
rect 4724 3194 4752 6190
rect 5276 5778 5304 6190
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4908 3534 4936 5510
rect 5276 5030 5304 5714
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5276 4690 5304 4966
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 5460 4010 5488 7686
rect 5552 6322 5580 7754
rect 5540 6316 5592 6322
rect 5736 6304 5764 10526
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5540 6258 5592 6264
rect 5644 6276 5764 6304
rect 5540 6180 5592 6186
rect 5540 6122 5592 6128
rect 5552 5030 5580 6122
rect 5644 6118 5672 6276
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5644 5642 5672 6054
rect 5632 5636 5684 5642
rect 5632 5578 5684 5584
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5552 3942 5580 4966
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 5184 3058 5212 3334
rect 5552 3194 5580 3334
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5356 3120 5408 3126
rect 5408 3068 5580 3074
rect 5356 3062 5580 3068
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 5172 3052 5224 3058
rect 5368 3046 5580 3062
rect 5172 2994 5224 3000
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 4712 2304 4764 2310
rect 4712 2246 4764 2252
rect 3988 2106 4016 2246
rect 3976 2100 4028 2106
rect 3976 2042 4028 2048
rect 4724 1494 4752 2246
rect 5000 1970 5028 2994
rect 5552 2825 5580 3046
rect 5538 2816 5594 2825
rect 5538 2751 5594 2760
rect 5262 2680 5318 2689
rect 5262 2615 5318 2624
rect 5276 2446 5304 2615
rect 5644 2514 5672 3878
rect 5828 3602 5856 10406
rect 5920 4010 5948 12838
rect 6012 11354 6040 15830
rect 6288 15570 6316 16934
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 6380 16250 6408 16390
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6276 15564 6328 15570
rect 6276 15506 6328 15512
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 6104 14498 6132 15098
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 6196 14618 6224 14962
rect 6184 14612 6236 14618
rect 6184 14554 6236 14560
rect 6104 14470 6224 14498
rect 6092 13932 6144 13938
rect 6092 13874 6144 13880
rect 6104 11694 6132 13874
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 6000 11076 6052 11082
rect 6000 11018 6052 11024
rect 6012 8090 6040 11018
rect 6104 10198 6132 11494
rect 6092 10192 6144 10198
rect 6092 10134 6144 10140
rect 6196 9926 6224 14470
rect 6380 13530 6408 16186
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 6276 13456 6328 13462
rect 6274 13424 6276 13433
rect 6328 13424 6330 13433
rect 6274 13359 6330 13368
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6380 12918 6408 13262
rect 6472 13190 6500 19382
rect 6642 19343 6698 19352
rect 6840 19310 6868 19751
rect 6932 19417 6960 19910
rect 7024 19514 7052 20470
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 7012 19508 7064 19514
rect 7012 19450 7064 19456
rect 6918 19408 6974 19417
rect 6918 19343 6974 19352
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6552 19168 6604 19174
rect 6552 19110 6604 19116
rect 6644 19168 6696 19174
rect 6644 19110 6696 19116
rect 6564 18902 6592 19110
rect 6552 18896 6604 18902
rect 6552 18838 6604 18844
rect 6656 18222 6684 19110
rect 7012 18692 7064 18698
rect 7012 18634 7064 18640
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 6932 18306 6960 18362
rect 6748 18278 6960 18306
rect 6644 18216 6696 18222
rect 6644 18158 6696 18164
rect 6552 18148 6604 18154
rect 6552 18090 6604 18096
rect 6564 17202 6592 18090
rect 6748 17610 6776 18278
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 6736 17604 6788 17610
rect 6736 17546 6788 17552
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6564 16658 6592 17138
rect 6840 17116 6868 17614
rect 6920 17128 6972 17134
rect 6840 17088 6920 17116
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6564 16096 6592 16594
rect 6840 16590 6868 17088
rect 6920 17070 6972 17076
rect 6920 16992 6972 16998
rect 6920 16934 6972 16940
rect 6828 16584 6880 16590
rect 6828 16526 6880 16532
rect 6644 16108 6696 16114
rect 6564 16068 6644 16096
rect 6644 16050 6696 16056
rect 6550 15192 6606 15201
rect 6550 15127 6606 15136
rect 6460 13184 6512 13190
rect 6460 13126 6512 13132
rect 6368 12912 6420 12918
rect 6368 12854 6420 12860
rect 6276 12300 6328 12306
rect 6276 12242 6328 12248
rect 6288 11218 6316 12242
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6276 11212 6328 11218
rect 6276 11154 6328 11160
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 5908 4004 5960 4010
rect 5908 3946 5960 3952
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 6012 2854 6040 4422
rect 6104 3369 6132 8774
rect 6472 7818 6500 11698
rect 6564 9976 6592 15127
rect 6656 14482 6684 16050
rect 6736 15632 6788 15638
rect 6734 15600 6736 15609
rect 6788 15600 6790 15609
rect 6734 15535 6790 15544
rect 6736 15496 6788 15502
rect 6840 15484 6868 16526
rect 6788 15456 6868 15484
rect 6736 15438 6788 15444
rect 6840 14958 6868 15456
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6644 14476 6696 14482
rect 6644 14418 6696 14424
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6642 13832 6698 13841
rect 6642 13767 6698 13776
rect 6656 11762 6684 13767
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6642 11520 6698 11529
rect 6642 11455 6698 11464
rect 6656 11354 6684 11455
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 6748 11014 6776 13874
rect 6840 13870 6868 14894
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6932 13258 6960 16934
rect 7024 14074 7052 18634
rect 7116 17746 7144 20334
rect 7196 20052 7248 20058
rect 7196 19994 7248 20000
rect 7208 18902 7236 19994
rect 7300 18970 7328 23666
rect 7392 23338 7420 24278
rect 7484 24274 7512 35566
rect 9140 31754 9168 36722
rect 9312 33312 9364 33318
rect 9312 33254 9364 33260
rect 9220 32428 9272 32434
rect 9220 32370 9272 32376
rect 9048 31726 9168 31754
rect 7656 30728 7708 30734
rect 7656 30670 7708 30676
rect 7564 24336 7616 24342
rect 7564 24278 7616 24284
rect 7472 24268 7524 24274
rect 7472 24210 7524 24216
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 7484 23497 7512 24006
rect 7576 23662 7604 24278
rect 7668 24206 7696 30670
rect 8300 29164 8352 29170
rect 8300 29106 8352 29112
rect 8208 27872 8260 27878
rect 8208 27814 8260 27820
rect 7840 27328 7892 27334
rect 7840 27270 7892 27276
rect 7852 26450 7880 27270
rect 7840 26444 7892 26450
rect 7840 26386 7892 26392
rect 7748 25900 7800 25906
rect 7748 25842 7800 25848
rect 7760 25226 7788 25842
rect 7840 25832 7892 25838
rect 7840 25774 7892 25780
rect 7748 25220 7800 25226
rect 7748 25162 7800 25168
rect 7656 24200 7708 24206
rect 7656 24142 7708 24148
rect 7654 23896 7710 23905
rect 7760 23866 7788 25162
rect 7654 23831 7710 23840
rect 7748 23860 7800 23866
rect 7668 23730 7696 23831
rect 7748 23802 7800 23808
rect 7656 23724 7708 23730
rect 7656 23666 7708 23672
rect 7564 23656 7616 23662
rect 7564 23598 7616 23604
rect 7470 23488 7526 23497
rect 7470 23423 7526 23432
rect 7392 23310 7696 23338
rect 7380 23112 7432 23118
rect 7380 23054 7432 23060
rect 7392 19802 7420 23054
rect 7472 22976 7524 22982
rect 7472 22918 7524 22924
rect 7564 22976 7616 22982
rect 7564 22918 7616 22924
rect 7484 22710 7512 22918
rect 7472 22704 7524 22710
rect 7472 22646 7524 22652
rect 7472 22160 7524 22166
rect 7472 22102 7524 22108
rect 7484 19961 7512 22102
rect 7576 20874 7604 22918
rect 7564 20868 7616 20874
rect 7564 20810 7616 20816
rect 7562 20496 7618 20505
rect 7562 20431 7618 20440
rect 7470 19952 7526 19961
rect 7576 19922 7604 20431
rect 7470 19887 7526 19896
rect 7564 19916 7616 19922
rect 7564 19858 7616 19864
rect 7392 19774 7604 19802
rect 7380 19440 7432 19446
rect 7380 19382 7432 19388
rect 7288 18964 7340 18970
rect 7288 18906 7340 18912
rect 7196 18896 7248 18902
rect 7196 18838 7248 18844
rect 7288 18692 7340 18698
rect 7288 18634 7340 18640
rect 7104 17740 7156 17746
rect 7104 17682 7156 17688
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 7116 15570 7144 15982
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 7196 15360 7248 15366
rect 7194 15328 7196 15337
rect 7248 15328 7250 15337
rect 7194 15263 7250 15272
rect 7300 15178 7328 18634
rect 7208 15150 7328 15178
rect 7102 14512 7158 14521
rect 7102 14447 7104 14456
rect 7156 14447 7158 14456
rect 7104 14418 7156 14424
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7116 13954 7144 14418
rect 7024 13926 7144 13954
rect 6920 13252 6972 13258
rect 6920 13194 6972 13200
rect 7024 12322 7052 13926
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 6932 12294 7052 12322
rect 6828 11824 6880 11830
rect 6826 11792 6828 11801
rect 6880 11792 6882 11801
rect 6826 11727 6882 11736
rect 6932 11336 6960 12294
rect 7116 12186 7144 13194
rect 7024 12158 7144 12186
rect 7024 11898 7052 12158
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 6840 11308 6960 11336
rect 6840 11098 6868 11308
rect 7116 11234 7144 11630
rect 6932 11218 7144 11234
rect 6920 11212 7144 11218
rect 6972 11206 7144 11212
rect 6920 11154 6972 11160
rect 6840 11070 7052 11098
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6920 10736 6972 10742
rect 6840 10696 6920 10724
rect 6734 10568 6790 10577
rect 6734 10503 6790 10512
rect 6644 9988 6696 9994
rect 6564 9948 6644 9976
rect 6564 9722 6592 9948
rect 6644 9930 6696 9936
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 6656 8974 6684 9658
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6656 7886 6684 8910
rect 6748 8906 6776 10503
rect 6736 8900 6788 8906
rect 6736 8842 6788 8848
rect 6748 8498 6776 8842
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6460 7812 6512 7818
rect 6460 7754 6512 7760
rect 6656 7546 6684 7822
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6564 6866 6592 7278
rect 6840 7002 6868 10696
rect 6920 10678 6972 10684
rect 6920 10260 6972 10266
rect 7024 10248 7052 11070
rect 6972 10220 7052 10248
rect 6920 10202 6972 10208
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6932 8974 6960 9862
rect 7116 9654 7144 11206
rect 7208 10146 7236 15150
rect 7288 14340 7340 14346
rect 7288 14282 7340 14288
rect 7300 13546 7328 14282
rect 7392 14074 7420 19382
rect 7472 19304 7524 19310
rect 7472 19246 7524 19252
rect 7484 18902 7512 19246
rect 7472 18896 7524 18902
rect 7472 18838 7524 18844
rect 7484 18698 7512 18838
rect 7472 18692 7524 18698
rect 7472 18634 7524 18640
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7484 16998 7512 18022
rect 7576 17610 7604 19774
rect 7668 19666 7696 23310
rect 7748 23112 7800 23118
rect 7746 23080 7748 23089
rect 7800 23080 7802 23089
rect 7746 23015 7802 23024
rect 7760 22574 7788 23015
rect 7748 22568 7800 22574
rect 7748 22510 7800 22516
rect 7748 22092 7800 22098
rect 7748 22034 7800 22040
rect 7760 20534 7788 22034
rect 7748 20528 7800 20534
rect 7748 20470 7800 20476
rect 7748 20324 7800 20330
rect 7748 20266 7800 20272
rect 7760 20058 7788 20266
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 7746 19816 7802 19825
rect 7746 19751 7748 19760
rect 7800 19751 7802 19760
rect 7852 19768 7880 25774
rect 7932 25424 7984 25430
rect 7932 25366 7984 25372
rect 7944 24750 7972 25366
rect 8024 25220 8076 25226
rect 8024 25162 8076 25168
rect 7932 24744 7984 24750
rect 7932 24686 7984 24692
rect 8036 22094 8064 25162
rect 8116 25152 8168 25158
rect 8116 25094 8168 25100
rect 8128 24818 8156 25094
rect 8220 24818 8248 27814
rect 8312 26586 8340 29106
rect 8392 28076 8444 28082
rect 8392 28018 8444 28024
rect 8404 27470 8432 28018
rect 8392 27464 8444 27470
rect 8392 27406 8444 27412
rect 8944 27464 8996 27470
rect 8944 27406 8996 27412
rect 8300 26580 8352 26586
rect 8300 26522 8352 26528
rect 8116 24812 8168 24818
rect 8116 24754 8168 24760
rect 8208 24812 8260 24818
rect 8208 24754 8260 24760
rect 8312 24682 8340 26522
rect 8208 24676 8260 24682
rect 8208 24618 8260 24624
rect 8300 24676 8352 24682
rect 8300 24618 8352 24624
rect 8852 24676 8904 24682
rect 8852 24618 8904 24624
rect 8220 24562 8248 24618
rect 8220 24534 8340 24562
rect 8208 24200 8260 24206
rect 8208 24142 8260 24148
rect 7944 22066 8064 22094
rect 7944 21894 7972 22066
rect 8114 21992 8170 22001
rect 8114 21927 8170 21936
rect 7932 21888 7984 21894
rect 7932 21830 7984 21836
rect 8128 21486 8156 21927
rect 8116 21480 8168 21486
rect 8116 21422 8168 21428
rect 8024 20596 8076 20602
rect 8024 20538 8076 20544
rect 7932 20392 7984 20398
rect 7930 20360 7932 20369
rect 7984 20360 7986 20369
rect 7930 20295 7986 20304
rect 8036 19786 8064 20538
rect 8024 19780 8076 19786
rect 7852 19740 7972 19768
rect 7748 19722 7800 19728
rect 7668 19638 7880 19666
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 7760 18154 7788 18906
rect 7748 18148 7800 18154
rect 7748 18090 7800 18096
rect 7654 17912 7710 17921
rect 7654 17847 7710 17856
rect 7564 17604 7616 17610
rect 7564 17546 7616 17552
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 7668 16522 7696 17847
rect 7852 17270 7880 19638
rect 7840 17264 7892 17270
rect 7840 17206 7892 17212
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 7656 16516 7708 16522
rect 7656 16458 7708 16464
rect 7470 16416 7526 16425
rect 7470 16351 7526 16360
rect 7484 15434 7512 16351
rect 7472 15428 7524 15434
rect 7472 15370 7524 15376
rect 7654 15056 7710 15065
rect 7654 14991 7710 15000
rect 7668 14958 7696 14991
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 7472 14340 7524 14346
rect 7472 14282 7524 14288
rect 7380 14068 7432 14074
rect 7380 14010 7432 14016
rect 7300 13518 7420 13546
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7300 10742 7328 11154
rect 7288 10736 7340 10742
rect 7288 10678 7340 10684
rect 7392 10282 7420 13518
rect 7484 10418 7512 14282
rect 7656 14272 7708 14278
rect 7656 14214 7708 14220
rect 7668 13938 7696 14214
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7760 13802 7788 16730
rect 7748 13796 7800 13802
rect 7748 13738 7800 13744
rect 7562 12472 7618 12481
rect 7760 12442 7788 13738
rect 7944 13530 7972 19740
rect 8024 19722 8076 19728
rect 8128 19666 8156 21422
rect 8220 21418 8248 24142
rect 8208 21412 8260 21418
rect 8208 21354 8260 21360
rect 8208 20528 8260 20534
rect 8208 20470 8260 20476
rect 8220 20058 8248 20470
rect 8208 20052 8260 20058
rect 8208 19994 8260 20000
rect 8036 19638 8156 19666
rect 8036 18698 8064 19638
rect 8114 19408 8170 19417
rect 8312 19394 8340 24534
rect 8864 24410 8892 24618
rect 8852 24404 8904 24410
rect 8852 24346 8904 24352
rect 8760 24268 8812 24274
rect 8760 24210 8812 24216
rect 8668 24200 8720 24206
rect 8668 24142 8720 24148
rect 8392 24132 8444 24138
rect 8392 24074 8444 24080
rect 8404 23633 8432 24074
rect 8390 23624 8446 23633
rect 8390 23559 8446 23568
rect 8392 23112 8444 23118
rect 8392 23054 8444 23060
rect 8404 22166 8432 23054
rect 8484 22704 8536 22710
rect 8484 22646 8536 22652
rect 8392 22160 8444 22166
rect 8392 22102 8444 22108
rect 8392 22024 8444 22030
rect 8392 21966 8444 21972
rect 8404 20618 8432 21966
rect 8496 20754 8524 22646
rect 8496 20726 8616 20754
rect 8404 20590 8524 20618
rect 8392 20528 8444 20534
rect 8392 20470 8444 20476
rect 8114 19343 8170 19352
rect 8220 19366 8340 19394
rect 8024 18692 8076 18698
rect 8024 18634 8076 18640
rect 8022 13968 8078 13977
rect 8022 13903 8078 13912
rect 8036 13802 8064 13903
rect 8024 13796 8076 13802
rect 8024 13738 8076 13744
rect 7932 13524 7984 13530
rect 7932 13466 7984 13472
rect 7562 12407 7618 12416
rect 7748 12436 7800 12442
rect 7576 12374 7604 12407
rect 7748 12378 7800 12384
rect 7564 12368 7616 12374
rect 7564 12310 7616 12316
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7748 12164 7800 12170
rect 7748 12106 7800 12112
rect 7484 10390 7696 10418
rect 7392 10254 7604 10282
rect 7208 10118 7420 10146
rect 7196 9988 7248 9994
rect 7196 9930 7248 9936
rect 7104 9648 7156 9654
rect 7104 9590 7156 9596
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7024 9042 7052 9522
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6564 4298 6592 5714
rect 6748 5166 6776 6802
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6840 5710 6868 6598
rect 6932 6390 6960 8910
rect 7024 8906 7052 8978
rect 7012 8900 7064 8906
rect 7012 8842 7064 8848
rect 7024 6458 7052 8842
rect 7102 8664 7158 8673
rect 7102 8599 7104 8608
rect 7156 8599 7158 8608
rect 7104 8570 7156 8576
rect 7208 8090 7236 9930
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6932 5273 6960 5850
rect 7024 5302 7052 6394
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7300 5642 7328 5850
rect 7288 5636 7340 5642
rect 7288 5578 7340 5584
rect 7012 5296 7064 5302
rect 6918 5264 6974 5273
rect 7012 5238 7064 5244
rect 6918 5199 6974 5208
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 7300 4706 7328 5578
rect 7392 4826 7420 10118
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7484 9110 7512 9862
rect 7472 9104 7524 9110
rect 7472 9046 7524 9052
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7116 4690 7328 4706
rect 7104 4684 7328 4690
rect 7156 4678 7328 4684
rect 7104 4626 7156 4632
rect 6564 4270 6684 4298
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6460 4072 6512 4078
rect 6460 4014 6512 4020
rect 6090 3360 6146 3369
rect 6090 3295 6146 3304
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 4988 1964 5040 1970
rect 4988 1906 5040 1912
rect 4712 1488 4764 1494
rect 4712 1430 4764 1436
rect 5184 800 5212 2246
rect 6472 800 6500 4014
rect 6564 3738 6592 4082
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 6656 3641 6684 4270
rect 7104 4208 7156 4214
rect 7156 4168 7236 4196
rect 7104 4150 7156 4156
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 6642 3632 6698 3641
rect 6642 3567 6698 3576
rect 7116 3466 7144 3878
rect 7104 3460 7156 3466
rect 7104 3402 7156 3408
rect 7208 3398 7236 4168
rect 7576 3505 7604 10254
rect 7668 9926 7696 10390
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7760 9178 7788 12106
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7852 8362 7880 12174
rect 7944 12102 7972 13466
rect 8128 12434 8156 19343
rect 8220 15026 8248 19366
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 8312 14346 8340 18566
rect 8404 16250 8432 20470
rect 8496 17338 8524 20590
rect 8588 19009 8616 20726
rect 8574 19000 8630 19009
rect 8574 18935 8630 18944
rect 8576 18828 8628 18834
rect 8576 18770 8628 18776
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8390 15736 8446 15745
rect 8390 15671 8446 15680
rect 8300 14340 8352 14346
rect 8300 14282 8352 14288
rect 8404 13433 8432 15671
rect 8496 14890 8524 16934
rect 8588 16454 8616 18770
rect 8680 18442 8708 24142
rect 8772 21350 8800 24210
rect 8852 22568 8904 22574
rect 8852 22510 8904 22516
rect 8864 21570 8892 22510
rect 8956 22094 8984 27406
rect 9048 24410 9076 31726
rect 9232 30938 9260 32370
rect 9220 30932 9272 30938
rect 9220 30874 9272 30880
rect 9128 25288 9180 25294
rect 9128 25230 9180 25236
rect 9140 24857 9168 25230
rect 9126 24848 9182 24857
rect 9182 24806 9260 24834
rect 9126 24783 9182 24792
rect 9128 24608 9180 24614
rect 9128 24550 9180 24556
rect 9036 24404 9088 24410
rect 9036 24346 9088 24352
rect 9140 23730 9168 24550
rect 9232 24138 9260 24806
rect 9220 24132 9272 24138
rect 9220 24074 9272 24080
rect 9324 23730 9352 33254
rect 9508 32570 9536 37130
rect 9692 37126 9720 39200
rect 9772 37256 9824 37262
rect 9772 37198 9824 37204
rect 9680 37120 9732 37126
rect 9680 37062 9732 37068
rect 9784 32570 9812 37198
rect 10980 37108 11008 39200
rect 12268 37244 12296 39200
rect 12440 37256 12492 37262
rect 12268 37216 12440 37244
rect 12440 37198 12492 37204
rect 11060 37120 11112 37126
rect 10980 37080 11060 37108
rect 11060 37062 11112 37068
rect 12440 37120 12492 37126
rect 12440 37062 12492 37068
rect 12900 37120 12952 37126
rect 13556 37108 13584 39200
rect 14200 37262 14228 39200
rect 14188 37256 14240 37262
rect 14188 37198 14240 37204
rect 14280 37256 14332 37262
rect 14280 37198 14332 37204
rect 14832 37256 14884 37262
rect 14832 37198 14884 37204
rect 13820 37120 13872 37126
rect 13556 37080 13820 37108
rect 12900 37062 12952 37068
rect 13820 37062 13872 37068
rect 10140 32768 10192 32774
rect 10140 32710 10192 32716
rect 10784 32768 10836 32774
rect 10784 32710 10836 32716
rect 9496 32564 9548 32570
rect 9496 32506 9548 32512
rect 9772 32564 9824 32570
rect 9772 32506 9824 32512
rect 9772 30864 9824 30870
rect 9772 30806 9824 30812
rect 9680 28008 9732 28014
rect 9680 27950 9732 27956
rect 9588 26512 9640 26518
rect 9588 26454 9640 26460
rect 9496 24608 9548 24614
rect 9496 24550 9548 24556
rect 9508 23730 9536 24550
rect 9128 23724 9180 23730
rect 9128 23666 9180 23672
rect 9312 23724 9364 23730
rect 9312 23666 9364 23672
rect 9496 23724 9548 23730
rect 9496 23666 9548 23672
rect 9600 23050 9628 26454
rect 9692 25838 9720 27950
rect 9680 25832 9732 25838
rect 9680 25774 9732 25780
rect 9692 24993 9720 25774
rect 9678 24984 9734 24993
rect 9678 24919 9734 24928
rect 9784 23610 9812 30806
rect 9864 30660 9916 30666
rect 9864 30602 9916 30608
rect 9692 23582 9812 23610
rect 9692 23186 9720 23582
rect 9772 23520 9824 23526
rect 9772 23462 9824 23468
rect 9680 23180 9732 23186
rect 9680 23122 9732 23128
rect 9588 23044 9640 23050
rect 9588 22986 9640 22992
rect 9404 22976 9456 22982
rect 9404 22918 9456 22924
rect 9416 22094 9444 22918
rect 9692 22710 9720 23122
rect 9680 22704 9732 22710
rect 9680 22646 9732 22652
rect 9588 22500 9640 22506
rect 9588 22442 9640 22448
rect 9600 22098 9628 22442
rect 9678 22128 9734 22137
rect 8956 22066 9076 22094
rect 9416 22066 9536 22094
rect 8956 21622 8984 21653
rect 8944 21616 8996 21622
rect 8864 21564 8944 21570
rect 8864 21558 8996 21564
rect 8864 21542 8984 21558
rect 8852 21480 8904 21486
rect 8852 21422 8904 21428
rect 8760 21344 8812 21350
rect 8760 21286 8812 21292
rect 8760 21140 8812 21146
rect 8760 21082 8812 21088
rect 8772 20466 8800 21082
rect 8760 20460 8812 20466
rect 8760 20402 8812 20408
rect 8864 20398 8892 21422
rect 8956 21418 8984 21542
rect 8944 21412 8996 21418
rect 8944 21354 8996 21360
rect 8942 20904 8998 20913
rect 8942 20839 8944 20848
rect 8996 20839 8998 20848
rect 8944 20810 8996 20816
rect 8852 20392 8904 20398
rect 8852 20334 8904 20340
rect 8942 20088 8998 20097
rect 8942 20023 8998 20032
rect 8760 19984 8812 19990
rect 8760 19926 8812 19932
rect 8772 19689 8800 19926
rect 8758 19680 8814 19689
rect 8758 19615 8814 19624
rect 8760 19304 8812 19310
rect 8812 19264 8892 19292
rect 8760 19246 8812 19252
rect 8864 18766 8892 19264
rect 8852 18760 8904 18766
rect 8852 18702 8904 18708
rect 8680 18426 8800 18442
rect 8680 18420 8812 18426
rect 8680 18414 8760 18420
rect 8760 18362 8812 18368
rect 8666 18320 8722 18329
rect 8666 18255 8722 18264
rect 8680 18222 8708 18255
rect 8668 18216 8720 18222
rect 8668 18158 8720 18164
rect 8758 17912 8814 17921
rect 8758 17847 8814 17856
rect 8772 17814 8800 17847
rect 8760 17808 8812 17814
rect 8760 17750 8812 17756
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 8680 16794 8708 17274
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8576 16448 8628 16454
rect 8772 16436 8800 17750
rect 8864 17678 8892 18702
rect 8852 17672 8904 17678
rect 8852 17614 8904 17620
rect 8864 17134 8892 17614
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8864 16658 8892 17070
rect 8852 16652 8904 16658
rect 8852 16594 8904 16600
rect 8576 16390 8628 16396
rect 8680 16408 8800 16436
rect 8680 16266 8708 16408
rect 8588 16238 8708 16266
rect 8484 14884 8536 14890
rect 8484 14826 8536 14832
rect 8588 13734 8616 16238
rect 8760 16108 8812 16114
rect 8760 16050 8812 16056
rect 8668 16040 8720 16046
rect 8772 16017 8800 16050
rect 8852 16040 8904 16046
rect 8668 15982 8720 15988
rect 8758 16008 8814 16017
rect 8576 13728 8628 13734
rect 8576 13670 8628 13676
rect 8390 13424 8446 13433
rect 8390 13359 8446 13368
rect 8128 12406 8432 12434
rect 8206 12336 8262 12345
rect 8206 12271 8262 12280
rect 8220 12238 8248 12271
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 8022 11656 8078 11665
rect 8022 11591 8078 11600
rect 8036 9450 8064 11591
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8312 10849 8340 11290
rect 8298 10840 8354 10849
rect 8298 10775 8354 10784
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 8312 10470 8340 10610
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 8024 9444 8076 9450
rect 8024 9386 8076 9392
rect 8128 9382 8156 9862
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 7840 8356 7892 8362
rect 7840 8298 7892 8304
rect 8128 7206 8156 9318
rect 8220 8974 8248 9454
rect 8404 9110 8432 12406
rect 8680 12238 8708 15982
rect 8852 15982 8904 15988
rect 8758 15943 8814 15952
rect 8864 15722 8892 15982
rect 8772 15694 8892 15722
rect 8772 13705 8800 15694
rect 8852 15632 8904 15638
rect 8852 15574 8904 15580
rect 8864 14006 8892 15574
rect 8852 14000 8904 14006
rect 8852 13942 8904 13948
rect 8852 13864 8904 13870
rect 8850 13832 8852 13841
rect 8904 13832 8906 13841
rect 8850 13767 8906 13776
rect 8758 13696 8814 13705
rect 8758 13631 8814 13640
rect 8956 12442 8984 20023
rect 9048 19446 9076 22066
rect 9508 21962 9536 22066
rect 9588 22092 9640 22098
rect 9678 22063 9734 22072
rect 9588 22034 9640 22040
rect 9404 21956 9456 21962
rect 9324 21916 9404 21944
rect 9324 21146 9352 21916
rect 9404 21898 9456 21904
rect 9496 21956 9548 21962
rect 9496 21898 9548 21904
rect 9402 21720 9458 21729
rect 9402 21655 9458 21664
rect 9312 21140 9364 21146
rect 9312 21082 9364 21088
rect 9416 21010 9444 21655
rect 9600 21418 9628 22034
rect 9692 21622 9720 22063
rect 9680 21616 9732 21622
rect 9680 21558 9732 21564
rect 9588 21412 9640 21418
rect 9588 21354 9640 21360
rect 9678 21040 9734 21049
rect 9404 21004 9456 21010
rect 9678 20975 9680 20984
rect 9404 20946 9456 20952
rect 9732 20975 9734 20984
rect 9680 20946 9732 20952
rect 9128 20936 9180 20942
rect 9128 20878 9180 20884
rect 9140 19961 9168 20878
rect 9220 20800 9272 20806
rect 9220 20742 9272 20748
rect 9404 20800 9456 20806
rect 9404 20742 9456 20748
rect 9126 19952 9182 19961
rect 9126 19887 9182 19896
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 9036 19440 9088 19446
rect 9036 19382 9088 19388
rect 9048 15162 9076 19382
rect 9140 17377 9168 19790
rect 9232 19718 9260 20742
rect 9312 20392 9364 20398
rect 9312 20334 9364 20340
rect 9324 20233 9352 20334
rect 9310 20224 9366 20233
rect 9310 20159 9366 20168
rect 9220 19712 9272 19718
rect 9220 19654 9272 19660
rect 9310 18728 9366 18737
rect 9416 18698 9444 20742
rect 9678 20632 9734 20641
rect 9678 20567 9734 20576
rect 9692 20398 9720 20567
rect 9680 20392 9732 20398
rect 9680 20334 9732 20340
rect 9496 20256 9548 20262
rect 9496 20198 9548 20204
rect 9508 19446 9536 20198
rect 9680 19780 9732 19786
rect 9680 19722 9732 19728
rect 9496 19440 9548 19446
rect 9496 19382 9548 19388
rect 9310 18663 9366 18672
rect 9404 18692 9456 18698
rect 9126 17368 9182 17377
rect 9126 17303 9182 17312
rect 9140 16425 9168 17303
rect 9220 16720 9272 16726
rect 9218 16688 9220 16697
rect 9272 16688 9274 16697
rect 9218 16623 9274 16632
rect 9324 16590 9352 18663
rect 9404 18634 9456 18640
rect 9416 16726 9444 18634
rect 9692 18154 9720 19722
rect 9784 18680 9812 23462
rect 9876 19922 9904 30602
rect 10048 27328 10100 27334
rect 10048 27270 10100 27276
rect 10060 24818 10088 27270
rect 10152 24954 10180 32710
rect 10796 32434 10824 32710
rect 10784 32428 10836 32434
rect 10784 32370 10836 32376
rect 12452 30734 12480 37062
rect 12912 30734 12940 37062
rect 14096 36780 14148 36786
rect 14096 36722 14148 36728
rect 13636 32904 13688 32910
rect 13636 32846 13688 32852
rect 12440 30728 12492 30734
rect 12440 30670 12492 30676
rect 12900 30728 12952 30734
rect 12900 30670 12952 30676
rect 10324 30592 10376 30598
rect 10324 30534 10376 30540
rect 13360 30592 13412 30598
rect 13360 30534 13412 30540
rect 10140 24948 10192 24954
rect 10140 24890 10192 24896
rect 10048 24812 10100 24818
rect 10048 24754 10100 24760
rect 10232 24064 10284 24070
rect 10232 24006 10284 24012
rect 10244 23497 10272 24006
rect 10230 23488 10286 23497
rect 10230 23423 10286 23432
rect 10336 23338 10364 30534
rect 13268 30388 13320 30394
rect 13268 30330 13320 30336
rect 11888 29504 11940 29510
rect 11888 29446 11940 29452
rect 11900 29170 11928 29446
rect 11888 29164 11940 29170
rect 11888 29106 11940 29112
rect 10600 29028 10652 29034
rect 10600 28970 10652 28976
rect 10612 27538 10640 28970
rect 12624 28076 12676 28082
rect 12624 28018 12676 28024
rect 11152 27872 11204 27878
rect 11152 27814 11204 27820
rect 10600 27532 10652 27538
rect 10600 27474 10652 27480
rect 11164 27130 11192 27814
rect 12072 27600 12124 27606
rect 12072 27542 12124 27548
rect 11980 27328 12032 27334
rect 11980 27270 12032 27276
rect 11152 27124 11204 27130
rect 11152 27066 11204 27072
rect 11060 26376 11112 26382
rect 11060 26318 11112 26324
rect 10692 25900 10744 25906
rect 10692 25842 10744 25848
rect 10704 25498 10732 25842
rect 10692 25492 10744 25498
rect 10692 25434 10744 25440
rect 10876 25288 10928 25294
rect 10876 25230 10928 25236
rect 10784 24948 10836 24954
rect 10784 24890 10836 24896
rect 10692 24676 10744 24682
rect 10692 24618 10744 24624
rect 10416 24200 10468 24206
rect 10416 24142 10468 24148
rect 10244 23310 10364 23338
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9968 21622 9996 21830
rect 9956 21616 10008 21622
rect 9956 21558 10008 21564
rect 10138 20904 10194 20913
rect 10138 20839 10140 20848
rect 10192 20839 10194 20848
rect 10140 20810 10192 20816
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 9864 19712 9916 19718
rect 9864 19654 9916 19660
rect 9876 18850 9904 19654
rect 10244 19174 10272 23310
rect 10324 22568 10376 22574
rect 10324 22510 10376 22516
rect 10336 20534 10364 22510
rect 10324 20528 10376 20534
rect 10324 20470 10376 20476
rect 10428 19514 10456 24142
rect 10600 23724 10652 23730
rect 10600 23666 10652 23672
rect 10506 21584 10562 21593
rect 10506 21519 10562 21528
rect 10416 19508 10468 19514
rect 10416 19450 10468 19456
rect 10324 19304 10376 19310
rect 10520 19258 10548 21519
rect 10324 19246 10376 19252
rect 10232 19168 10284 19174
rect 10046 19136 10102 19145
rect 10232 19110 10284 19116
rect 10046 19071 10102 19080
rect 10060 18970 10088 19071
rect 10336 18986 10364 19246
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 10244 18958 10364 18986
rect 10428 19230 10548 19258
rect 9876 18822 9996 18850
rect 9864 18692 9916 18698
rect 9784 18652 9864 18680
rect 9864 18634 9916 18640
rect 9680 18148 9732 18154
rect 9680 18090 9732 18096
rect 9404 16720 9456 16726
rect 9404 16662 9456 16668
rect 9312 16584 9364 16590
rect 9310 16552 9312 16561
rect 9364 16552 9366 16561
rect 9310 16487 9366 16496
rect 9680 16516 9732 16522
rect 9680 16458 9732 16464
rect 9126 16416 9182 16425
rect 9126 16351 9182 16360
rect 9310 16008 9366 16017
rect 9310 15943 9366 15952
rect 9126 15736 9182 15745
rect 9126 15671 9128 15680
rect 9180 15671 9182 15680
rect 9128 15642 9180 15648
rect 9324 15502 9352 15943
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9494 15192 9550 15201
rect 9036 15156 9088 15162
rect 9494 15127 9496 15136
rect 9036 15098 9088 15104
rect 9548 15127 9550 15136
rect 9496 15098 9548 15104
rect 9404 15088 9456 15094
rect 9403 15036 9404 15076
rect 9456 15036 9536 15042
rect 9403 15014 9536 15036
rect 9036 14952 9088 14958
rect 9404 14952 9456 14958
rect 9036 14894 9088 14900
rect 9324 14912 9404 14940
rect 9048 14482 9076 14894
rect 9324 14793 9352 14912
rect 9404 14894 9456 14900
rect 9404 14816 9456 14822
rect 9310 14784 9366 14793
rect 9404 14758 9456 14764
rect 9310 14719 9366 14728
rect 9310 14512 9366 14521
rect 9036 14476 9088 14482
rect 9310 14447 9366 14456
rect 9036 14418 9088 14424
rect 9324 12442 9352 14447
rect 9416 14385 9444 14758
rect 9402 14376 9458 14385
rect 9402 14311 9458 14320
rect 8944 12436 8996 12442
rect 8944 12378 8996 12384
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 8944 11552 8996 11558
rect 8942 11520 8944 11529
rect 8996 11520 8998 11529
rect 8942 11455 8998 11464
rect 8956 11286 8984 11455
rect 8944 11280 8996 11286
rect 8944 11222 8996 11228
rect 9048 11082 9076 12174
rect 9508 12170 9536 15014
rect 9692 12850 9720 16458
rect 9968 16046 9996 18822
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 10060 18465 10088 18566
rect 10046 18456 10102 18465
rect 10046 18391 10102 18400
rect 10048 18216 10100 18222
rect 10046 18184 10048 18193
rect 10100 18184 10102 18193
rect 10046 18119 10102 18128
rect 10046 17776 10102 17785
rect 10046 17711 10102 17720
rect 10060 17610 10088 17711
rect 10048 17604 10100 17610
rect 10048 17546 10100 17552
rect 10060 17338 10088 17546
rect 10048 17332 10100 17338
rect 10048 17274 10100 17280
rect 10152 17134 10180 18906
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 10244 17066 10272 18958
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10336 18290 10364 18566
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10428 17490 10456 19230
rect 10508 19168 10560 19174
rect 10508 19110 10560 19116
rect 10336 17462 10456 17490
rect 10232 17060 10284 17066
rect 10232 17002 10284 17008
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 9956 16040 10008 16046
rect 9956 15982 10008 15988
rect 10152 15570 10180 16050
rect 10140 15564 10192 15570
rect 10140 15506 10192 15512
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9784 12918 9812 13330
rect 9772 12912 9824 12918
rect 9772 12854 9824 12860
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9784 12322 9812 12854
rect 9692 12294 9812 12322
rect 9692 12238 9720 12294
rect 9680 12232 9732 12238
rect 9876 12220 9904 15438
rect 9956 15360 10008 15366
rect 9956 15302 10008 15308
rect 9968 13938 9996 15302
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9954 13832 10010 13841
rect 9954 13767 10010 13776
rect 9680 12174 9732 12180
rect 9784 12192 9904 12220
rect 9496 12164 9548 12170
rect 9496 12106 9548 12112
rect 9692 11830 9720 12174
rect 9220 11824 9272 11830
rect 9220 11766 9272 11772
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9232 11354 9260 11766
rect 9678 11656 9734 11665
rect 9416 11626 9678 11642
rect 9404 11620 9678 11626
rect 9456 11614 9678 11620
rect 9678 11591 9734 11600
rect 9404 11562 9456 11568
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 9310 11112 9366 11121
rect 9036 11076 9088 11082
rect 9310 11047 9366 11056
rect 9036 11018 9088 11024
rect 9128 10532 9180 10538
rect 9128 10474 9180 10480
rect 8576 10124 8628 10130
rect 8576 10066 8628 10072
rect 8588 9654 8616 10066
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8956 9178 8984 9522
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 8392 9104 8444 9110
rect 8392 9046 8444 9052
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8220 8430 8248 8910
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8208 6792 8260 6798
rect 7654 6760 7710 6769
rect 8208 6734 8260 6740
rect 7654 6695 7710 6704
rect 7668 6662 7696 6695
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7746 4720 7802 4729
rect 7746 4655 7802 4664
rect 7562 3496 7618 3505
rect 7562 3431 7618 3440
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 6932 2514 6960 2926
rect 7024 2774 7052 3334
rect 7286 3088 7342 3097
rect 7576 3058 7604 3431
rect 7760 3058 7788 4655
rect 7930 4584 7986 4593
rect 7930 4519 7932 4528
rect 7984 4519 7986 4528
rect 8116 4548 8168 4554
rect 7932 4490 7984 4496
rect 8116 4490 8168 4496
rect 8128 4457 8156 4490
rect 8114 4448 8170 4457
rect 8114 4383 8170 4392
rect 8128 4078 8156 4383
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 8128 3126 8156 3606
rect 8116 3120 8168 3126
rect 8116 3062 8168 3068
rect 7286 3023 7342 3032
rect 7564 3052 7616 3058
rect 7024 2746 7144 2774
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 7116 800 7144 2746
rect 7300 1562 7328 3023
rect 7564 2994 7616 3000
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 8220 2666 8248 6734
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8404 5710 8432 6054
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8392 5704 8444 5710
rect 8390 5672 8392 5681
rect 8444 5672 8446 5681
rect 8390 5607 8446 5616
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8312 4282 8340 5170
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8312 3602 8340 4218
rect 8390 3632 8446 3641
rect 8300 3596 8352 3602
rect 8390 3567 8392 3576
rect 8300 3538 8352 3544
rect 8444 3567 8446 3576
rect 8392 3538 8444 3544
rect 8312 3040 8340 3538
rect 8392 3052 8444 3058
rect 8312 3012 8392 3040
rect 8392 2994 8444 3000
rect 8496 2854 8524 5714
rect 8588 5166 8616 7142
rect 8668 6384 8720 6390
rect 8668 6326 8720 6332
rect 8680 6118 8708 6326
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8680 5953 8708 6054
rect 8666 5944 8722 5953
rect 8666 5879 8722 5888
rect 8864 5778 8892 7278
rect 9048 6866 9076 7822
rect 9140 7478 9168 10474
rect 9128 7472 9180 7478
rect 9128 7414 9180 7420
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8864 5302 8892 5714
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8956 4049 8984 6802
rect 9048 6322 9076 6802
rect 9324 6798 9352 11047
rect 9508 10742 9536 11494
rect 9784 11393 9812 12192
rect 9864 12096 9916 12102
rect 9864 12038 9916 12044
rect 9770 11384 9826 11393
rect 9770 11319 9826 11328
rect 9784 11286 9812 11319
rect 9772 11280 9824 11286
rect 9772 11222 9824 11228
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9678 10976 9734 10985
rect 9678 10911 9734 10920
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 9588 10736 9640 10742
rect 9588 10678 9640 10684
rect 9600 10577 9628 10678
rect 9586 10568 9642 10577
rect 9586 10503 9642 10512
rect 9692 10266 9720 10911
rect 9784 10810 9812 11086
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9692 9738 9720 9930
rect 9600 9710 9720 9738
rect 9600 9489 9628 9710
rect 9680 9512 9732 9518
rect 9586 9480 9642 9489
rect 9680 9454 9732 9460
rect 9586 9415 9642 9424
rect 9692 8906 9720 9454
rect 9784 9042 9812 10746
rect 9876 10062 9904 12038
rect 9968 11898 9996 13767
rect 10152 12434 10180 15506
rect 10244 13734 10272 17002
rect 10336 14074 10364 17462
rect 10414 15736 10470 15745
rect 10414 15671 10470 15680
rect 10428 15638 10456 15671
rect 10416 15632 10468 15638
rect 10416 15574 10468 15580
rect 10520 14958 10548 19110
rect 10612 17921 10640 23666
rect 10704 19310 10732 24618
rect 10796 21010 10824 24890
rect 10888 24818 10916 25230
rect 10876 24812 10928 24818
rect 10876 24754 10928 24760
rect 10888 24682 10916 24754
rect 10876 24676 10928 24682
rect 10876 24618 10928 24624
rect 11072 24614 11100 26318
rect 11060 24608 11112 24614
rect 11060 24550 11112 24556
rect 11060 24064 11112 24070
rect 11060 24006 11112 24012
rect 10876 23656 10928 23662
rect 10876 23598 10928 23604
rect 10888 21321 10916 23598
rect 11072 22710 11100 24006
rect 11164 23866 11192 27066
rect 11244 26988 11296 26994
rect 11244 26930 11296 26936
rect 11256 26586 11284 26930
rect 11244 26580 11296 26586
rect 11244 26522 11296 26528
rect 11152 23860 11204 23866
rect 11152 23802 11204 23808
rect 11152 22976 11204 22982
rect 11152 22918 11204 22924
rect 11060 22704 11112 22710
rect 11060 22646 11112 22652
rect 11060 22160 11112 22166
rect 11060 22102 11112 22108
rect 11072 21865 11100 22102
rect 11164 21962 11192 22918
rect 11152 21956 11204 21962
rect 11152 21898 11204 21904
rect 11058 21856 11114 21865
rect 11058 21791 11114 21800
rect 10968 21548 11020 21554
rect 10968 21490 11020 21496
rect 10980 21457 11008 21490
rect 10966 21448 11022 21457
rect 10966 21383 11022 21392
rect 10874 21312 10930 21321
rect 10874 21247 10930 21256
rect 10784 21004 10836 21010
rect 10784 20946 10836 20952
rect 10782 20496 10838 20505
rect 10782 20431 10784 20440
rect 10836 20431 10838 20440
rect 10784 20402 10836 20408
rect 10692 19304 10744 19310
rect 10692 19246 10744 19252
rect 10598 17912 10654 17921
rect 10598 17847 10654 17856
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10704 17377 10732 17478
rect 10690 17368 10746 17377
rect 10690 17303 10746 17312
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10612 16590 10640 17138
rect 10692 17060 10744 17066
rect 10692 17002 10744 17008
rect 10704 16726 10732 17002
rect 10692 16720 10744 16726
rect 10692 16662 10744 16668
rect 10600 16584 10652 16590
rect 10600 16526 10652 16532
rect 10612 16046 10640 16526
rect 10600 16040 10652 16046
rect 10600 15982 10652 15988
rect 10612 15502 10640 15982
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10508 14952 10560 14958
rect 10508 14894 10560 14900
rect 10612 14482 10640 15438
rect 10796 15178 10824 20402
rect 10888 19718 10916 21247
rect 10966 21040 11022 21049
rect 10966 20975 11022 20984
rect 10980 19786 11008 20975
rect 11150 19952 11206 19961
rect 11150 19887 11206 19896
rect 10968 19780 11020 19786
rect 10968 19722 11020 19728
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10980 19334 11008 19722
rect 10888 19306 11008 19334
rect 11060 19372 11112 19378
rect 11060 19314 11112 19320
rect 10888 18630 10916 19306
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10874 18456 10930 18465
rect 10874 18391 10930 18400
rect 10888 18358 10916 18391
rect 10876 18352 10928 18358
rect 10876 18294 10928 18300
rect 10980 18154 11008 19110
rect 10968 18148 11020 18154
rect 10968 18090 11020 18096
rect 10876 17808 10928 17814
rect 10874 17776 10876 17785
rect 10928 17776 10930 17785
rect 10874 17711 10930 17720
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10888 15366 10916 17614
rect 11072 17270 11100 19314
rect 11164 17678 11192 19887
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 11152 17536 11204 17542
rect 11150 17504 11152 17513
rect 11204 17504 11206 17513
rect 11150 17439 11206 17448
rect 11150 17368 11206 17377
rect 11150 17303 11206 17312
rect 11164 17270 11192 17303
rect 11060 17264 11112 17270
rect 11060 17206 11112 17212
rect 11152 17264 11204 17270
rect 11152 17206 11204 17212
rect 10966 16688 11022 16697
rect 10966 16623 11022 16632
rect 10980 16522 11008 16623
rect 10968 16516 11020 16522
rect 10968 16458 11020 16464
rect 10980 16114 11008 16458
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 11152 16448 11204 16454
rect 11152 16390 11204 16396
rect 11072 16114 11100 16390
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 11164 15994 11192 16390
rect 10980 15966 11192 15994
rect 10980 15910 11008 15966
rect 10968 15904 11020 15910
rect 10968 15846 11020 15852
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 11150 15328 11206 15337
rect 11150 15263 11206 15272
rect 10796 15150 10916 15178
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10336 13841 10364 14010
rect 10704 13977 10732 14758
rect 10690 13968 10746 13977
rect 10690 13903 10692 13912
rect 10744 13903 10746 13912
rect 10692 13874 10744 13880
rect 10704 13843 10732 13874
rect 10322 13832 10378 13841
rect 10322 13767 10378 13776
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 10782 13696 10838 13705
rect 10782 13631 10838 13640
rect 10690 13424 10746 13433
rect 10690 13359 10746 13368
rect 10230 12880 10286 12889
rect 10230 12815 10286 12824
rect 10244 12646 10272 12815
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 10336 12646 10364 12718
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10060 12406 10180 12434
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 10060 11082 10088 12406
rect 10140 11824 10192 11830
rect 10140 11766 10192 11772
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9864 9172 9916 9178
rect 9864 9114 9916 9120
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9876 8974 9904 9114
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9954 8936 10010 8945
rect 9680 8900 9732 8906
rect 9954 8871 9956 8880
rect 9680 8842 9732 8848
rect 10008 8871 10010 8880
rect 9956 8842 10008 8848
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9678 7032 9734 7041
rect 9784 7002 9812 7754
rect 9862 7576 9918 7585
rect 9968 7546 9996 8842
rect 9862 7511 9918 7520
rect 9956 7540 10008 7546
rect 9678 6967 9680 6976
rect 9732 6967 9734 6976
rect 9772 6996 9824 7002
rect 9680 6938 9732 6944
rect 9772 6938 9824 6944
rect 9678 6896 9734 6905
rect 9678 6831 9734 6840
rect 9692 6798 9720 6831
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 9036 5636 9088 5642
rect 9036 5578 9088 5584
rect 9048 5409 9076 5578
rect 9034 5400 9090 5409
rect 9034 5335 9090 5344
rect 9232 4282 9260 6734
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9692 5642 9720 6598
rect 9876 6254 9904 7511
rect 9956 7482 10008 7488
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9876 5234 9904 6190
rect 10060 6118 10088 11018
rect 10152 8430 10180 11766
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10140 8424 10192 8430
rect 10140 8366 10192 8372
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 9310 4856 9366 4865
rect 9310 4791 9366 4800
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 8942 4040 8998 4049
rect 8942 3975 8998 3984
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 8680 2990 8708 3538
rect 9324 3534 9352 4791
rect 9404 4684 9456 4690
rect 9404 4626 9456 4632
rect 9416 4146 9444 4626
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 9692 4214 9720 4422
rect 9588 4208 9640 4214
rect 9586 4176 9588 4185
rect 9680 4208 9732 4214
rect 9640 4176 9642 4185
rect 9404 4140 9456 4146
rect 9680 4150 9732 4156
rect 9586 4111 9642 4120
rect 9404 4082 9456 4088
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9402 3768 9458 3777
rect 9402 3703 9458 3712
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9128 3460 9180 3466
rect 9128 3402 9180 3408
rect 8668 2984 8720 2990
rect 8668 2926 8720 2932
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8220 2638 8432 2666
rect 9140 2650 9168 3402
rect 7748 2576 7800 2582
rect 7748 2518 7800 2524
rect 7760 2446 7788 2518
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 7840 2304 7892 2310
rect 7840 2246 7892 2252
rect 7852 2038 7880 2246
rect 7840 2032 7892 2038
rect 7840 1974 7892 1980
rect 7288 1556 7340 1562
rect 7288 1498 7340 1504
rect 8404 800 8432 2638
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 9324 2582 9352 3470
rect 9312 2576 9364 2582
rect 9312 2518 9364 2524
rect 9416 2378 9444 3703
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9784 3398 9812 3538
rect 9876 3534 9904 3878
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9692 3126 9720 3334
rect 9496 3120 9548 3126
rect 9496 3062 9548 3068
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 9508 2938 9536 3062
rect 9968 2990 9996 4422
rect 10152 3398 10180 8230
rect 10244 3398 10272 8366
rect 10336 7818 10364 8774
rect 10324 7812 10376 7818
rect 10324 7754 10376 7760
rect 10428 6662 10456 12718
rect 10600 10736 10652 10742
rect 10600 10678 10652 10684
rect 10612 10577 10640 10678
rect 10704 10606 10732 13359
rect 10692 10600 10744 10606
rect 10598 10568 10654 10577
rect 10692 10542 10744 10548
rect 10598 10503 10654 10512
rect 10796 10062 10824 13631
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 10784 9648 10836 9654
rect 10784 9590 10836 9596
rect 10692 8560 10744 8566
rect 10692 8502 10744 8508
rect 10506 6896 10562 6905
rect 10506 6831 10562 6840
rect 10520 6798 10548 6831
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10324 6180 10376 6186
rect 10324 6122 10376 6128
rect 10336 5914 10364 6122
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 9956 2984 10008 2990
rect 9508 2910 9720 2938
rect 9956 2926 10008 2932
rect 9404 2372 9456 2378
rect 9404 2314 9456 2320
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 8496 1902 8524 2246
rect 8484 1896 8536 1902
rect 8484 1838 8536 1844
rect 9692 800 9720 2910
rect 10152 2446 10180 3334
rect 10336 2922 10364 5170
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 10324 2916 10376 2922
rect 10324 2858 10376 2864
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 10428 1737 10456 4966
rect 10508 4276 10560 4282
rect 10508 4218 10560 4224
rect 10520 2553 10548 4218
rect 10506 2544 10562 2553
rect 10506 2479 10562 2488
rect 10612 1834 10640 5578
rect 10704 3126 10732 8502
rect 10796 7177 10824 9590
rect 10888 7562 10916 15150
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11072 12850 11100 13126
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 10968 12096 11020 12102
rect 10966 12064 10968 12073
rect 11020 12064 11022 12073
rect 10966 11999 11022 12008
rect 11072 10742 11100 12786
rect 11060 10736 11112 10742
rect 11060 10678 11112 10684
rect 11072 9654 11100 10678
rect 11164 9994 11192 15263
rect 11256 13462 11284 26522
rect 11428 26308 11480 26314
rect 11428 26250 11480 26256
rect 11440 26217 11468 26250
rect 11426 26208 11482 26217
rect 11426 26143 11482 26152
rect 11428 25424 11480 25430
rect 11428 25366 11480 25372
rect 11336 23112 11388 23118
rect 11336 23054 11388 23060
rect 11348 21962 11376 23054
rect 11336 21956 11388 21962
rect 11336 21898 11388 21904
rect 11336 21548 11388 21554
rect 11336 21490 11388 21496
rect 11348 16658 11376 21490
rect 11440 18970 11468 25366
rect 11520 24744 11572 24750
rect 11520 24686 11572 24692
rect 11532 22094 11560 24686
rect 11704 23724 11756 23730
rect 11704 23666 11756 23672
rect 11716 23633 11744 23666
rect 11702 23624 11758 23633
rect 11702 23559 11758 23568
rect 11612 23520 11664 23526
rect 11796 23520 11848 23526
rect 11664 23480 11744 23508
rect 11612 23462 11664 23468
rect 11716 22094 11744 23480
rect 11796 23462 11848 23468
rect 11808 22710 11836 23462
rect 11796 22704 11848 22710
rect 11796 22646 11848 22652
rect 11886 22128 11942 22137
rect 11532 22066 11652 22094
rect 11716 22066 11836 22094
rect 11428 18964 11480 18970
rect 11428 18906 11480 18912
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 11532 18630 11560 18770
rect 11428 18624 11480 18630
rect 11428 18566 11480 18572
rect 11520 18624 11572 18630
rect 11520 18566 11572 18572
rect 11440 18154 11468 18566
rect 11428 18148 11480 18154
rect 11428 18090 11480 18096
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 11440 14550 11468 17818
rect 11428 14544 11480 14550
rect 11428 14486 11480 14492
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11348 14249 11376 14350
rect 11334 14240 11390 14249
rect 11334 14175 11390 14184
rect 11244 13456 11296 13462
rect 11244 13398 11296 13404
rect 11256 13326 11284 13398
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11348 12850 11376 14175
rect 11532 14074 11560 18566
rect 11624 18272 11652 22066
rect 11704 21344 11756 21350
rect 11704 21286 11756 21292
rect 11716 19009 11744 21286
rect 11808 20874 11836 22066
rect 11886 22063 11942 22072
rect 11900 21962 11928 22063
rect 11888 21956 11940 21962
rect 11888 21898 11940 21904
rect 11796 20868 11848 20874
rect 11796 20810 11848 20816
rect 11888 20528 11940 20534
rect 11888 20470 11940 20476
rect 11900 20058 11928 20470
rect 11888 20052 11940 20058
rect 11888 19994 11940 20000
rect 11992 19530 12020 27270
rect 12084 26450 12112 27542
rect 12636 27334 12664 28018
rect 13176 27464 13228 27470
rect 13176 27406 13228 27412
rect 12624 27328 12676 27334
rect 12624 27270 12676 27276
rect 12716 27328 12768 27334
rect 12716 27270 12768 27276
rect 12728 27062 12756 27270
rect 12716 27056 12768 27062
rect 12716 26998 12768 27004
rect 12716 26920 12768 26926
rect 12452 26880 12716 26908
rect 12164 26784 12216 26790
rect 12164 26726 12216 26732
rect 12072 26444 12124 26450
rect 12072 26386 12124 26392
rect 12176 26314 12204 26726
rect 12256 26512 12308 26518
rect 12256 26454 12308 26460
rect 12164 26308 12216 26314
rect 12164 26250 12216 26256
rect 12072 24608 12124 24614
rect 12072 24550 12124 24556
rect 12084 22778 12112 24550
rect 12162 22944 12218 22953
rect 12162 22879 12218 22888
rect 12072 22772 12124 22778
rect 12072 22714 12124 22720
rect 12072 22568 12124 22574
rect 12072 22510 12124 22516
rect 12084 22166 12112 22510
rect 12072 22160 12124 22166
rect 12072 22102 12124 22108
rect 12072 22024 12124 22030
rect 12072 21966 12124 21972
rect 11808 19502 12020 19530
rect 12084 19530 12112 21966
rect 12176 21010 12204 22879
rect 12268 22574 12296 26454
rect 12452 26450 12480 26880
rect 12716 26862 12768 26868
rect 13188 26586 13216 27406
rect 12992 26580 13044 26586
rect 12992 26522 13044 26528
rect 13176 26580 13228 26586
rect 13176 26522 13228 26528
rect 12440 26444 12492 26450
rect 12440 26386 12492 26392
rect 12452 23798 12480 26386
rect 13004 26382 13032 26522
rect 13280 26466 13308 30330
rect 13188 26438 13308 26466
rect 12992 26376 13044 26382
rect 12992 26318 13044 26324
rect 12716 24676 12768 24682
rect 12716 24618 12768 24624
rect 12728 24410 12756 24618
rect 12716 24404 12768 24410
rect 12716 24346 12768 24352
rect 12532 24200 12584 24206
rect 12532 24142 12584 24148
rect 12544 23798 12572 24142
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 12808 24132 12860 24138
rect 12808 24074 12860 24080
rect 12440 23792 12492 23798
rect 12440 23734 12492 23740
rect 12532 23792 12584 23798
rect 12532 23734 12584 23740
rect 12636 23730 12664 24074
rect 12624 23724 12676 23730
rect 12624 23666 12676 23672
rect 12716 22976 12768 22982
rect 12714 22944 12716 22953
rect 12768 22944 12770 22953
rect 12714 22879 12770 22888
rect 12256 22568 12308 22574
rect 12256 22510 12308 22516
rect 12622 22128 12678 22137
rect 12622 22063 12678 22072
rect 12440 21956 12492 21962
rect 12440 21898 12492 21904
rect 12452 21690 12480 21898
rect 12440 21684 12492 21690
rect 12440 21626 12492 21632
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 12256 21412 12308 21418
rect 12256 21354 12308 21360
rect 12268 21321 12296 21354
rect 12254 21312 12310 21321
rect 12254 21247 12310 21256
rect 12164 21004 12216 21010
rect 12164 20946 12216 20952
rect 12256 19780 12308 19786
rect 12256 19722 12308 19728
rect 12084 19502 12204 19530
rect 11702 19000 11758 19009
rect 11702 18935 11758 18944
rect 11624 18244 11744 18272
rect 11612 18148 11664 18154
rect 11612 18090 11664 18096
rect 11624 16250 11652 18090
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11612 14272 11664 14278
rect 11716 14249 11744 18244
rect 11808 17762 11836 19502
rect 11980 19440 12032 19446
rect 11980 19382 12032 19388
rect 12072 19440 12124 19446
rect 12072 19382 12124 19388
rect 11888 18964 11940 18970
rect 11888 18906 11940 18912
rect 11900 18358 11928 18906
rect 11888 18352 11940 18358
rect 11888 18294 11940 18300
rect 11808 17734 11928 17762
rect 11796 17672 11848 17678
rect 11796 17614 11848 17620
rect 11808 17202 11836 17614
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11900 17082 11928 17734
rect 11808 17054 11928 17082
rect 11808 14906 11836 17054
rect 11886 16960 11942 16969
rect 11886 16895 11942 16904
rect 11900 15094 11928 16895
rect 11992 16454 12020 19382
rect 12084 19310 12112 19382
rect 12072 19304 12124 19310
rect 12072 19246 12124 19252
rect 12176 18680 12204 19502
rect 12268 18970 12296 19722
rect 12348 19236 12400 19242
rect 12348 19178 12400 19184
rect 12360 19145 12388 19178
rect 12346 19136 12402 19145
rect 12346 19071 12402 19080
rect 12346 19000 12402 19009
rect 12256 18964 12308 18970
rect 12346 18935 12402 18944
rect 12256 18906 12308 18912
rect 12256 18828 12308 18834
rect 12256 18770 12308 18776
rect 12084 18652 12204 18680
rect 12084 17864 12112 18652
rect 12268 18630 12296 18770
rect 12360 18766 12388 18935
rect 12348 18760 12400 18766
rect 12348 18702 12400 18708
rect 12256 18624 12308 18630
rect 12162 18592 12218 18601
rect 12256 18566 12308 18572
rect 12162 18527 12218 18536
rect 12176 18086 12204 18527
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 12084 17836 12296 17864
rect 12164 17740 12216 17746
rect 12164 17682 12216 17688
rect 12176 17338 12204 17682
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12268 17270 12296 17836
rect 12452 17649 12480 21490
rect 12532 21344 12584 21350
rect 12532 21286 12584 21292
rect 12544 20534 12572 21286
rect 12636 21010 12664 22063
rect 12714 21992 12770 22001
rect 12714 21927 12716 21936
rect 12768 21927 12770 21936
rect 12716 21898 12768 21904
rect 12820 21729 12848 24074
rect 12900 23792 12952 23798
rect 12900 23734 12952 23740
rect 12806 21720 12862 21729
rect 12806 21655 12862 21664
rect 12624 21004 12676 21010
rect 12624 20946 12676 20952
rect 12532 20528 12584 20534
rect 12532 20470 12584 20476
rect 12808 20460 12860 20466
rect 12808 20402 12860 20408
rect 12716 20324 12768 20330
rect 12716 20266 12768 20272
rect 12532 19780 12584 19786
rect 12532 19722 12584 19728
rect 12544 18834 12572 19722
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12544 17746 12572 17818
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 12438 17640 12494 17649
rect 12348 17604 12400 17610
rect 12438 17575 12494 17584
rect 12348 17546 12400 17552
rect 12256 17264 12308 17270
rect 12256 17206 12308 17212
rect 12268 16810 12296 17206
rect 12360 16969 12388 17546
rect 12346 16960 12402 16969
rect 12346 16895 12402 16904
rect 12176 16782 12296 16810
rect 12346 16824 12402 16833
rect 12072 16720 12124 16726
rect 12072 16662 12124 16668
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 12084 15688 12112 16662
rect 11992 15660 12112 15688
rect 11888 15088 11940 15094
rect 11888 15030 11940 15036
rect 11808 14878 11928 14906
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11612 14214 11664 14220
rect 11702 14240 11758 14249
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 11348 12345 11376 12786
rect 11334 12336 11390 12345
rect 11624 12306 11652 14214
rect 11702 14175 11758 14184
rect 11704 13932 11756 13938
rect 11808 13920 11836 14758
rect 11756 13892 11836 13920
rect 11704 13874 11756 13880
rect 11716 12306 11744 13874
rect 11900 12714 11928 14878
rect 11992 14498 12020 15660
rect 12070 15600 12126 15609
rect 12070 15535 12072 15544
rect 12124 15535 12126 15544
rect 12072 15506 12124 15512
rect 12072 15020 12124 15026
rect 12072 14962 12124 14968
rect 12084 14822 12112 14962
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 12176 14550 12204 16782
rect 12346 16759 12402 16768
rect 12256 16516 12308 16522
rect 12256 16458 12308 16464
rect 12268 16425 12296 16458
rect 12254 16416 12310 16425
rect 12254 16351 12310 16360
rect 12360 15570 12388 16759
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 12530 16552 12586 16561
rect 12452 15638 12480 16526
rect 12530 16487 12586 16496
rect 12544 16454 12572 16487
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12544 15706 12572 16390
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12440 15632 12492 15638
rect 12440 15574 12492 15580
rect 12348 15564 12400 15570
rect 12348 15506 12400 15512
rect 12360 14618 12388 15506
rect 12636 15434 12664 17818
rect 12624 15428 12676 15434
rect 12624 15370 12676 15376
rect 12532 15088 12584 15094
rect 12532 15030 12584 15036
rect 12544 14822 12572 15030
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12164 14544 12216 14550
rect 11992 14470 12112 14498
rect 12164 14486 12216 14492
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11992 13802 12020 14350
rect 11980 13796 12032 13802
rect 11980 13738 12032 13744
rect 11980 13524 12032 13530
rect 11980 13466 12032 13472
rect 11992 12782 12020 13466
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11888 12708 11940 12714
rect 11888 12650 11940 12656
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 11334 12271 11390 12280
rect 11612 12300 11664 12306
rect 11348 10674 11376 12271
rect 11612 12242 11664 12248
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11808 12170 11836 12582
rect 11796 12164 11848 12170
rect 11796 12106 11848 12112
rect 11520 12096 11572 12102
rect 11520 12038 11572 12044
rect 11426 11384 11482 11393
rect 11426 11319 11482 11328
rect 11440 11132 11468 11319
rect 11532 11286 11560 12038
rect 11612 11824 11664 11830
rect 11612 11766 11664 11772
rect 11624 11506 11652 11766
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11624 11478 11744 11506
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11520 11280 11572 11286
rect 11520 11222 11572 11228
rect 11440 11104 11560 11132
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 11440 10441 11468 10950
rect 11426 10432 11482 10441
rect 11426 10367 11482 10376
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 10966 9480 11022 9489
rect 10966 9415 10968 9424
rect 11020 9415 11022 9424
rect 11426 9480 11482 9489
rect 11426 9415 11482 9424
rect 10968 9386 11020 9392
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 11072 8634 11100 8774
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 10888 7534 11284 7562
rect 10968 7472 11020 7478
rect 10966 7440 10968 7449
rect 11020 7440 11022 7449
rect 10966 7375 11022 7384
rect 10782 7168 10838 7177
rect 10782 7103 10838 7112
rect 11150 7032 11206 7041
rect 11150 6967 11206 6976
rect 11164 6866 11192 6967
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 10876 6724 10928 6730
rect 10876 6666 10928 6672
rect 10888 3602 10916 6666
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11072 6458 11100 6598
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 11164 6322 11192 6802
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 11072 5370 11100 5510
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11164 5234 11192 6258
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 10692 3120 10744 3126
rect 10692 3062 10744 3068
rect 10874 2680 10930 2689
rect 10874 2615 10930 2624
rect 10888 2446 10916 2615
rect 10876 2440 10928 2446
rect 10980 2417 11008 5170
rect 11164 4690 11192 5170
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11072 2582 11100 4558
rect 11164 3602 11192 4626
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11164 3058 11192 3402
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11256 2650 11284 7534
rect 11440 6730 11468 9415
rect 11428 6724 11480 6730
rect 11428 6666 11480 6672
rect 11336 6384 11388 6390
rect 11336 6326 11388 6332
rect 11348 3913 11376 6326
rect 11428 4480 11480 4486
rect 11428 4422 11480 4428
rect 11440 4282 11468 4422
rect 11428 4276 11480 4282
rect 11428 4218 11480 4224
rect 11532 4146 11560 11104
rect 11624 11014 11652 11290
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11716 9897 11744 11478
rect 11702 9888 11758 9897
rect 11702 9823 11758 9832
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 11612 8016 11664 8022
rect 11612 7958 11664 7964
rect 11624 7750 11652 7958
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 11716 6390 11744 9590
rect 11808 8922 11836 11698
rect 11992 11529 12020 12582
rect 12084 11665 12112 14470
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12348 14408 12400 14414
rect 12268 14368 12348 14396
rect 12164 11756 12216 11762
rect 12268 11744 12296 14368
rect 12348 14350 12400 14356
rect 12544 13705 12572 14418
rect 12728 13870 12756 20266
rect 12820 19310 12848 20402
rect 12808 19304 12860 19310
rect 12808 19246 12860 19252
rect 12808 18692 12860 18698
rect 12912 18680 12940 23734
rect 13084 23248 13136 23254
rect 13084 23190 13136 23196
rect 12992 20528 13044 20534
rect 12992 20470 13044 20476
rect 13004 19990 13032 20470
rect 12992 19984 13044 19990
rect 12992 19926 13044 19932
rect 12990 19544 13046 19553
rect 12990 19479 13046 19488
rect 13004 18834 13032 19479
rect 13096 19378 13124 23190
rect 13188 21690 13216 26438
rect 13372 24750 13400 30534
rect 13648 25362 13676 32846
rect 14108 30394 14136 36722
rect 14292 36650 14320 37198
rect 14844 36922 14872 37198
rect 15488 37126 15516 39200
rect 15476 37120 15528 37126
rect 15476 37062 15528 37068
rect 16776 36922 16804 39200
rect 17420 37126 17448 39200
rect 18512 37324 18564 37330
rect 18512 37266 18564 37272
rect 17408 37120 17460 37126
rect 17408 37062 17460 37068
rect 14832 36916 14884 36922
rect 14832 36858 14884 36864
rect 16764 36916 16816 36922
rect 16764 36858 16816 36864
rect 16856 36780 16908 36786
rect 16856 36722 16908 36728
rect 14280 36644 14332 36650
rect 14280 36586 14332 36592
rect 15384 31952 15436 31958
rect 15384 31894 15436 31900
rect 14096 30388 14148 30394
rect 14096 30330 14148 30336
rect 14280 29572 14332 29578
rect 14280 29514 14332 29520
rect 14188 25900 14240 25906
rect 14188 25842 14240 25848
rect 14096 25696 14148 25702
rect 14096 25638 14148 25644
rect 13636 25356 13688 25362
rect 13636 25298 13688 25304
rect 13360 24744 13412 24750
rect 13360 24686 13412 24692
rect 13372 23186 13400 24686
rect 13648 24274 13676 25298
rect 13636 24268 13688 24274
rect 13636 24210 13688 24216
rect 14108 24138 14136 25638
rect 14096 24132 14148 24138
rect 14096 24074 14148 24080
rect 13912 24064 13964 24070
rect 13912 24006 13964 24012
rect 13924 23594 13952 24006
rect 13912 23588 13964 23594
rect 13912 23530 13964 23536
rect 13360 23180 13412 23186
rect 13360 23122 13412 23128
rect 13268 22636 13320 22642
rect 13268 22578 13320 22584
rect 13176 21684 13228 21690
rect 13176 21626 13228 21632
rect 13176 21548 13228 21554
rect 13280 21536 13308 22578
rect 13820 22432 13872 22438
rect 13820 22374 13872 22380
rect 13544 21956 13596 21962
rect 13544 21898 13596 21904
rect 13728 21956 13780 21962
rect 13728 21898 13780 21904
rect 13556 21690 13584 21898
rect 13452 21684 13504 21690
rect 13452 21626 13504 21632
rect 13544 21684 13596 21690
rect 13544 21626 13596 21632
rect 13228 21508 13308 21536
rect 13176 21490 13228 21496
rect 13084 19372 13136 19378
rect 13084 19314 13136 19320
rect 13188 18902 13216 21490
rect 13358 20904 13414 20913
rect 13358 20839 13360 20848
rect 13412 20839 13414 20848
rect 13360 20810 13412 20816
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13280 19922 13308 20402
rect 13360 20324 13412 20330
rect 13360 20266 13412 20272
rect 13268 19916 13320 19922
rect 13268 19858 13320 19864
rect 13372 19786 13400 20266
rect 13360 19780 13412 19786
rect 13360 19722 13412 19728
rect 13464 19530 13492 21626
rect 13740 21554 13768 21898
rect 13728 21548 13780 21554
rect 13728 21490 13780 21496
rect 13636 21480 13688 21486
rect 13636 21422 13688 21428
rect 13648 21078 13676 21422
rect 13728 21344 13780 21350
rect 13728 21286 13780 21292
rect 13544 21072 13596 21078
rect 13542 21040 13544 21049
rect 13636 21072 13688 21078
rect 13596 21040 13598 21049
rect 13636 21014 13688 21020
rect 13542 20975 13598 20984
rect 13740 20942 13768 21286
rect 13832 21010 13860 22374
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 13912 21344 13964 21350
rect 13912 21286 13964 21292
rect 14004 21344 14056 21350
rect 14004 21286 14056 21292
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 13728 20936 13780 20942
rect 13728 20878 13780 20884
rect 13544 20800 13596 20806
rect 13544 20742 13596 20748
rect 13556 20466 13584 20742
rect 13924 20482 13952 21286
rect 14016 20602 14044 21286
rect 14004 20596 14056 20602
rect 14004 20538 14056 20544
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13832 20454 13952 20482
rect 13832 19718 13860 20454
rect 13912 20392 13964 20398
rect 13912 20334 13964 20340
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13360 19508 13412 19514
rect 13464 19502 13584 19530
rect 13360 19450 13412 19456
rect 13176 18896 13228 18902
rect 13176 18838 13228 18844
rect 12992 18828 13044 18834
rect 12992 18770 13044 18776
rect 13084 18828 13136 18834
rect 13084 18770 13136 18776
rect 12912 18652 13032 18680
rect 12808 18634 12860 18640
rect 12820 16522 12848 18634
rect 13004 18442 13032 18652
rect 12912 18414 13032 18442
rect 12808 16516 12860 16522
rect 12808 16458 12860 16464
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12820 15570 12848 16050
rect 12912 15745 12940 18414
rect 12992 18352 13044 18358
rect 13096 18329 13124 18770
rect 12992 18294 13044 18300
rect 13082 18320 13138 18329
rect 12898 15736 12954 15745
rect 13004 15706 13032 18294
rect 13082 18255 13138 18264
rect 13096 18222 13124 18255
rect 13084 18216 13136 18222
rect 13084 18158 13136 18164
rect 13372 18154 13400 19450
rect 13452 19372 13504 19378
rect 13452 19314 13504 19320
rect 13360 18148 13412 18154
rect 13360 18090 13412 18096
rect 13082 17912 13138 17921
rect 13082 17847 13138 17856
rect 13096 17542 13124 17847
rect 13360 17604 13412 17610
rect 13360 17546 13412 17552
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 13372 17241 13400 17546
rect 13358 17232 13414 17241
rect 13358 17167 13414 17176
rect 13176 16788 13228 16794
rect 13176 16730 13228 16736
rect 12898 15671 12954 15680
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 12806 15464 12862 15473
rect 12806 15399 12862 15408
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12530 13696 12586 13705
rect 12530 13631 12586 13640
rect 12714 13560 12770 13569
rect 12714 13495 12770 13504
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12360 13161 12388 13330
rect 12346 13152 12402 13161
rect 12346 13087 12402 13096
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12452 12889 12480 12922
rect 12438 12880 12494 12889
rect 12438 12815 12494 12824
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 12636 12646 12664 12786
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12728 12594 12756 13495
rect 12820 12730 12848 15399
rect 12992 15360 13044 15366
rect 13188 15337 13216 16730
rect 13266 16280 13322 16289
rect 13266 16215 13322 16224
rect 13360 16244 13412 16250
rect 13280 15978 13308 16215
rect 13360 16186 13412 16192
rect 13268 15972 13320 15978
rect 13268 15914 13320 15920
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 12992 15302 13044 15308
rect 13174 15328 13230 15337
rect 13004 12850 13032 15302
rect 13174 15263 13230 15272
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 13096 14346 13124 14554
rect 13084 14340 13136 14346
rect 13084 14282 13136 14288
rect 13084 12912 13136 12918
rect 13082 12880 13084 12889
rect 13136 12880 13138 12889
rect 12992 12844 13044 12850
rect 13082 12815 13138 12824
rect 12992 12786 13044 12792
rect 12820 12702 13032 12730
rect 12728 12566 12848 12594
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12216 11716 12296 11744
rect 12164 11698 12216 11704
rect 12452 11665 12480 11834
rect 12070 11656 12126 11665
rect 12438 11656 12494 11665
rect 12070 11591 12126 11600
rect 12164 11620 12216 11626
rect 12438 11591 12494 11600
rect 12164 11562 12216 11568
rect 12176 11529 12204 11562
rect 11978 11520 12034 11529
rect 11978 11455 12034 11464
rect 12162 11520 12218 11529
rect 12162 11455 12218 11464
rect 12438 11520 12494 11529
rect 12438 11455 12494 11464
rect 12452 11354 12480 11455
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11900 10577 11928 10610
rect 11886 10568 11942 10577
rect 11886 10503 11942 10512
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 11900 10266 11928 10406
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11992 9654 12020 11154
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 11900 9110 11928 9454
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 11808 8894 11928 8922
rect 11704 6384 11756 6390
rect 11704 6326 11756 6332
rect 11610 5400 11666 5409
rect 11610 5335 11666 5344
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11334 3904 11390 3913
rect 11334 3839 11390 3848
rect 11348 3482 11376 3839
rect 11348 3466 11468 3482
rect 11348 3460 11480 3466
rect 11348 3454 11428 3460
rect 11428 3402 11480 3408
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 10876 2382 10928 2388
rect 10966 2408 11022 2417
rect 11532 2378 11560 4082
rect 11624 4010 11652 5335
rect 11716 5302 11744 6326
rect 11704 5296 11756 5302
rect 11704 5238 11756 5244
rect 11612 4004 11664 4010
rect 11612 3946 11664 3952
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11716 3738 11744 3878
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 11624 2854 11652 3674
rect 11900 3058 11928 8894
rect 11992 8566 12020 9590
rect 11980 8560 12032 8566
rect 11980 8502 12032 8508
rect 11992 7954 12020 8502
rect 12084 8090 12112 10678
rect 12176 10577 12204 11018
rect 12268 10810 12296 11154
rect 12348 11076 12400 11082
rect 12348 11018 12400 11024
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12162 10568 12218 10577
rect 12162 10503 12218 10512
rect 12360 10441 12388 11018
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12162 10432 12218 10441
rect 12162 10367 12218 10376
rect 12346 10432 12402 10441
rect 12346 10367 12402 10376
rect 12176 10266 12204 10367
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12452 10033 12480 10950
rect 12544 10810 12572 12106
rect 12622 11928 12678 11937
rect 12622 11863 12678 11872
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12636 10538 12664 11863
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12820 11642 12848 12566
rect 13004 12434 13032 12702
rect 13188 12617 13216 14758
rect 13280 14550 13308 15438
rect 13268 14544 13320 14550
rect 13268 14486 13320 14492
rect 13280 13462 13308 14486
rect 13268 13456 13320 13462
rect 13268 13398 13320 13404
rect 13266 12744 13322 12753
rect 13266 12679 13322 12688
rect 13280 12646 13308 12679
rect 13268 12640 13320 12646
rect 13174 12608 13230 12617
rect 13268 12582 13320 12588
rect 13174 12543 13230 12552
rect 13174 12472 13230 12481
rect 13004 12406 13124 12434
rect 13174 12407 13230 12416
rect 12992 12300 13044 12306
rect 12992 12242 13044 12248
rect 13004 11762 13032 12242
rect 13096 12102 13124 12406
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 12728 10742 12756 11630
rect 12820 11614 13032 11642
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12912 10062 12940 10950
rect 12900 10056 12952 10062
rect 12438 10024 12494 10033
rect 12900 9998 12952 10004
rect 12438 9959 12494 9968
rect 12624 9988 12676 9994
rect 12624 9930 12676 9936
rect 12346 9888 12402 9897
rect 12346 9823 12402 9832
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 12268 9382 12296 9522
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12256 9172 12308 9178
rect 12360 9160 12388 9823
rect 12636 9178 12664 9930
rect 12308 9132 12388 9160
rect 12256 9114 12308 9120
rect 12360 8974 12388 9132
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12532 9104 12584 9110
rect 12452 9052 12532 9058
rect 12452 9046 12584 9052
rect 12452 9030 12572 9046
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 11992 7478 12020 7890
rect 11980 7472 12032 7478
rect 11980 7414 12032 7420
rect 12176 5166 12204 8842
rect 12452 8838 12480 9030
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12544 8294 12572 8774
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12532 8288 12584 8294
rect 12532 8230 12584 8236
rect 12254 6624 12310 6633
rect 12254 6559 12310 6568
rect 12268 6186 12296 6559
rect 12256 6180 12308 6186
rect 12256 6122 12308 6128
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12452 5914 12480 6054
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12636 5681 12664 8570
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12728 7342 12756 8026
rect 12912 7750 12940 9998
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 13004 7342 13032 11614
rect 13188 10742 13216 12407
rect 13268 12096 13320 12102
rect 13266 12064 13268 12073
rect 13320 12064 13322 12073
rect 13266 11999 13322 12008
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13176 10736 13228 10742
rect 13176 10678 13228 10684
rect 13280 9654 13308 11834
rect 13372 9722 13400 16186
rect 13464 13870 13492 19314
rect 13556 18834 13584 19502
rect 13924 19310 13952 20334
rect 14004 19916 14056 19922
rect 14004 19858 14056 19864
rect 13912 19304 13964 19310
rect 13912 19246 13964 19252
rect 13544 18828 13596 18834
rect 13544 18770 13596 18776
rect 13912 18760 13964 18766
rect 13912 18702 13964 18708
rect 13636 18692 13688 18698
rect 13636 18634 13688 18640
rect 13648 18601 13676 18634
rect 13634 18592 13690 18601
rect 13634 18527 13690 18536
rect 13542 18456 13598 18465
rect 13542 18391 13598 18400
rect 13556 18358 13584 18391
rect 13544 18352 13596 18358
rect 13544 18294 13596 18300
rect 13636 18352 13688 18358
rect 13636 18294 13688 18300
rect 13648 18193 13676 18294
rect 13634 18184 13690 18193
rect 13634 18119 13690 18128
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13556 15026 13584 18022
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 13636 17536 13688 17542
rect 13636 17478 13688 17484
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13648 14362 13676 17478
rect 13726 17368 13782 17377
rect 13726 17303 13782 17312
rect 13740 17134 13768 17303
rect 13832 17270 13860 17682
rect 13820 17264 13872 17270
rect 13820 17206 13872 17212
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 13740 16794 13768 17070
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13820 16176 13872 16182
rect 13820 16118 13872 16124
rect 13832 15994 13860 16118
rect 13740 15966 13860 15994
rect 13740 15473 13768 15966
rect 13924 15892 13952 18702
rect 13832 15864 13952 15892
rect 13726 15464 13782 15473
rect 13726 15399 13782 15408
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13740 14822 13768 14962
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13556 14334 13676 14362
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 13464 13433 13492 13806
rect 13450 13424 13506 13433
rect 13450 13359 13506 13368
rect 13556 13258 13584 14334
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13648 14006 13676 14214
rect 13636 14000 13688 14006
rect 13636 13942 13688 13948
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13648 13258 13676 13670
rect 13544 13252 13596 13258
rect 13544 13194 13596 13200
rect 13636 13252 13688 13258
rect 13636 13194 13688 13200
rect 13452 12912 13504 12918
rect 13452 12854 13504 12860
rect 13464 12306 13492 12854
rect 13636 12776 13688 12782
rect 13634 12744 13636 12753
rect 13688 12744 13690 12753
rect 13634 12679 13690 12688
rect 13542 12472 13598 12481
rect 13542 12407 13544 12416
rect 13596 12407 13598 12416
rect 13544 12378 13596 12384
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13832 11393 13860 15864
rect 13912 14068 13964 14074
rect 13912 14010 13964 14016
rect 13818 11384 13874 11393
rect 13818 11319 13874 11328
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 13268 9648 13320 9654
rect 13268 9590 13320 9596
rect 13452 7472 13504 7478
rect 13452 7414 13504 7420
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 12728 7002 12756 7278
rect 13464 7041 13492 7414
rect 13450 7032 13506 7041
rect 12716 6996 12768 7002
rect 13450 6967 13506 6976
rect 12716 6938 12768 6944
rect 13268 6928 13320 6934
rect 13174 6896 13230 6905
rect 13268 6870 13320 6876
rect 13174 6831 13230 6840
rect 13188 6798 13216 6831
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13280 6458 13308 6870
rect 13556 6866 13584 11018
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13740 9926 13768 10542
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13832 10130 13860 10406
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13832 9586 13860 10066
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13726 9072 13782 9081
rect 13832 9042 13860 9522
rect 13726 9007 13728 9016
rect 13780 9007 13782 9016
rect 13820 9036 13872 9042
rect 13728 8978 13780 8984
rect 13820 8978 13872 8984
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13648 8537 13676 8570
rect 13634 8528 13690 8537
rect 13832 8498 13860 8978
rect 13924 8974 13952 14010
rect 14016 13954 14044 19858
rect 14108 17814 14136 21966
rect 14096 17808 14148 17814
rect 14096 17750 14148 17756
rect 14096 16720 14148 16726
rect 14200 16708 14228 25842
rect 14292 22094 14320 29514
rect 14832 26580 14884 26586
rect 14832 26522 14884 26528
rect 14372 26376 14424 26382
rect 14370 26344 14372 26353
rect 14424 26344 14426 26353
rect 14370 26279 14426 26288
rect 14740 25696 14792 25702
rect 14740 25638 14792 25644
rect 14372 25152 14424 25158
rect 14372 25094 14424 25100
rect 14464 25152 14516 25158
rect 14464 25094 14516 25100
rect 14384 24274 14412 25094
rect 14372 24268 14424 24274
rect 14372 24210 14424 24216
rect 14476 24138 14504 25094
rect 14752 24886 14780 25638
rect 14740 24880 14792 24886
rect 14740 24822 14792 24828
rect 14844 24750 14872 26522
rect 15016 25900 15068 25906
rect 15016 25842 15068 25848
rect 14832 24744 14884 24750
rect 14832 24686 14884 24692
rect 14924 24744 14976 24750
rect 14924 24686 14976 24692
rect 14832 24268 14884 24274
rect 14832 24210 14884 24216
rect 14464 24132 14516 24138
rect 14464 24074 14516 24080
rect 14844 23662 14872 24210
rect 14832 23656 14884 23662
rect 14832 23598 14884 23604
rect 14464 23520 14516 23526
rect 14464 23462 14516 23468
rect 14476 23050 14504 23462
rect 14740 23180 14792 23186
rect 14740 23122 14792 23128
rect 14464 23044 14516 23050
rect 14464 22986 14516 22992
rect 14648 22772 14700 22778
rect 14648 22714 14700 22720
rect 14660 22098 14688 22714
rect 14292 22066 14412 22094
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14292 20777 14320 20878
rect 14278 20768 14334 20777
rect 14278 20703 14334 20712
rect 14384 19786 14412 22066
rect 14648 22092 14700 22098
rect 14648 22034 14700 22040
rect 14648 20936 14700 20942
rect 14648 20878 14700 20884
rect 14660 20602 14688 20878
rect 14648 20596 14700 20602
rect 14648 20538 14700 20544
rect 14372 19780 14424 19786
rect 14372 19722 14424 19728
rect 14384 19689 14412 19722
rect 14370 19680 14426 19689
rect 14370 19615 14426 19624
rect 14280 19508 14332 19514
rect 14280 19450 14332 19456
rect 14292 17678 14320 19450
rect 14372 19304 14424 19310
rect 14372 19246 14424 19252
rect 14384 18222 14412 19246
rect 14752 19009 14780 23122
rect 14844 19242 14872 23598
rect 14936 20942 14964 24686
rect 15028 23118 15056 25842
rect 15292 25696 15344 25702
rect 15292 25638 15344 25644
rect 15304 25226 15332 25638
rect 15292 25220 15344 25226
rect 15292 25162 15344 25168
rect 15200 25152 15252 25158
rect 15200 25094 15252 25100
rect 15212 24886 15240 25094
rect 15292 24948 15344 24954
rect 15292 24890 15344 24896
rect 15200 24880 15252 24886
rect 15200 24822 15252 24828
rect 15304 24750 15332 24890
rect 15292 24744 15344 24750
rect 15292 24686 15344 24692
rect 15292 24608 15344 24614
rect 15292 24550 15344 24556
rect 15304 24274 15332 24550
rect 15292 24268 15344 24274
rect 15292 24210 15344 24216
rect 15396 23798 15424 31894
rect 16764 29708 16816 29714
rect 16764 29650 16816 29656
rect 16212 29640 16264 29646
rect 16212 29582 16264 29588
rect 16224 28558 16252 29582
rect 16672 29164 16724 29170
rect 16672 29106 16724 29112
rect 15752 28552 15804 28558
rect 15752 28494 15804 28500
rect 16212 28552 16264 28558
rect 16212 28494 16264 28500
rect 15764 27538 15792 28494
rect 15752 27532 15804 27538
rect 15752 27474 15804 27480
rect 15476 25288 15528 25294
rect 15476 25230 15528 25236
rect 15488 24614 15516 25230
rect 15476 24608 15528 24614
rect 15476 24550 15528 24556
rect 15660 24336 15712 24342
rect 15660 24278 15712 24284
rect 15384 23792 15436 23798
rect 15384 23734 15436 23740
rect 15672 23662 15700 24278
rect 15660 23656 15712 23662
rect 15660 23598 15712 23604
rect 15016 23112 15068 23118
rect 15068 23060 15148 23066
rect 15016 23054 15148 23060
rect 15028 23038 15148 23054
rect 15014 21856 15070 21865
rect 15014 21791 15070 21800
rect 15028 21622 15056 21791
rect 15016 21616 15068 21622
rect 15016 21558 15068 21564
rect 15028 21418 15056 21558
rect 15016 21412 15068 21418
rect 15016 21354 15068 21360
rect 14924 20936 14976 20942
rect 14924 20878 14976 20884
rect 15120 20448 15148 23038
rect 15200 22976 15252 22982
rect 15200 22918 15252 22924
rect 15212 20534 15240 22918
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 15200 20528 15252 20534
rect 15200 20470 15252 20476
rect 14936 20420 15148 20448
rect 14832 19236 14884 19242
rect 14832 19178 14884 19184
rect 14738 19000 14794 19009
rect 14738 18935 14794 18944
rect 14740 18896 14792 18902
rect 14740 18838 14792 18844
rect 14464 18624 14516 18630
rect 14464 18566 14516 18572
rect 14372 18216 14424 18222
rect 14372 18158 14424 18164
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14292 17218 14320 17614
rect 14292 17190 14412 17218
rect 14280 16992 14332 16998
rect 14278 16960 14280 16969
rect 14332 16960 14334 16969
rect 14278 16895 14334 16904
rect 14148 16680 14228 16708
rect 14096 16662 14148 16668
rect 14200 14890 14228 16680
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14292 16046 14320 16526
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 14384 14890 14412 17190
rect 14476 16182 14504 18566
rect 14556 17740 14608 17746
rect 14556 17682 14608 17688
rect 14568 17270 14596 17682
rect 14556 17264 14608 17270
rect 14556 17206 14608 17212
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 14568 16658 14596 17070
rect 14556 16652 14608 16658
rect 14556 16594 14608 16600
rect 14752 16538 14780 18838
rect 14832 18216 14884 18222
rect 14832 18158 14884 18164
rect 14660 16522 14780 16538
rect 14648 16516 14780 16522
rect 14700 16510 14780 16516
rect 14648 16458 14700 16464
rect 14464 16176 14516 16182
rect 14464 16118 14516 16124
rect 14462 15872 14518 15881
rect 14462 15807 14518 15816
rect 14476 15366 14504 15807
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14464 15360 14516 15366
rect 14464 15302 14516 15308
rect 14188 14884 14240 14890
rect 14188 14826 14240 14832
rect 14372 14884 14424 14890
rect 14372 14826 14424 14832
rect 14464 14816 14516 14822
rect 14464 14758 14516 14764
rect 14016 13926 14228 13954
rect 14002 13288 14058 13297
rect 14002 13223 14058 13232
rect 14016 11014 14044 13223
rect 14200 11354 14228 13926
rect 14372 13864 14424 13870
rect 14278 13832 14334 13841
rect 14372 13806 14424 13812
rect 14278 13767 14334 13776
rect 14292 12434 14320 13767
rect 14384 13258 14412 13806
rect 14476 13258 14504 14758
rect 14568 14657 14596 15438
rect 14554 14648 14610 14657
rect 14554 14583 14610 14592
rect 14556 14340 14608 14346
rect 14556 14282 14608 14288
rect 14568 13394 14596 14282
rect 14660 13734 14688 16458
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14752 14006 14780 15302
rect 14740 14000 14792 14006
rect 14740 13942 14792 13948
rect 14648 13728 14700 13734
rect 14648 13670 14700 13676
rect 14556 13388 14608 13394
rect 14556 13330 14608 13336
rect 14372 13252 14424 13258
rect 14372 13194 14424 13200
rect 14464 13252 14516 13258
rect 14464 13194 14516 13200
rect 14292 12406 14504 12434
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 14094 11248 14150 11257
rect 14094 11183 14150 11192
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 14016 9761 14044 9998
rect 14002 9752 14058 9761
rect 14002 9687 14058 9696
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13634 8463 13690 8472
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 14108 7954 14136 11183
rect 14200 11082 14228 11290
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14188 11076 14240 11082
rect 14188 11018 14240 11024
rect 14188 10192 14240 10198
rect 14188 10134 14240 10140
rect 14200 9722 14228 10134
rect 14292 10130 14320 11086
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14384 10266 14412 10610
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14476 9926 14504 12406
rect 14568 12306 14596 13330
rect 14844 13258 14872 18158
rect 14936 14618 14964 20420
rect 15016 19780 15068 19786
rect 15016 19722 15068 19728
rect 15108 19780 15160 19786
rect 15108 19722 15160 19728
rect 15028 19553 15056 19722
rect 15014 19544 15070 19553
rect 15014 19479 15070 19488
rect 15120 18057 15148 19722
rect 15304 19718 15332 21830
rect 15660 21616 15712 21622
rect 15660 21558 15712 21564
rect 15476 21072 15528 21078
rect 15476 21014 15528 21020
rect 15488 20942 15516 21014
rect 15476 20936 15528 20942
rect 15672 20913 15700 21558
rect 15476 20878 15528 20884
rect 15658 20904 15714 20913
rect 15384 20800 15436 20806
rect 15382 20768 15384 20777
rect 15436 20768 15438 20777
rect 15382 20703 15438 20712
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15212 18578 15240 19246
rect 15396 18698 15424 20703
rect 15488 19258 15516 20878
rect 15658 20839 15714 20848
rect 15568 19712 15620 19718
rect 15568 19654 15620 19660
rect 15580 19446 15608 19654
rect 15568 19440 15620 19446
rect 15568 19382 15620 19388
rect 15488 19230 15608 19258
rect 15384 18692 15436 18698
rect 15384 18634 15436 18640
rect 15476 18692 15528 18698
rect 15476 18634 15528 18640
rect 15212 18550 15424 18578
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 15106 18048 15162 18057
rect 15106 17983 15162 17992
rect 15016 17604 15068 17610
rect 15016 17546 15068 17552
rect 15028 16794 15056 17546
rect 15016 16788 15068 16794
rect 15016 16730 15068 16736
rect 15212 16153 15240 18226
rect 15290 18184 15346 18193
rect 15290 18119 15346 18128
rect 15198 16144 15254 16153
rect 15198 16079 15254 16088
rect 15304 15994 15332 18119
rect 15108 15972 15160 15978
rect 15108 15914 15160 15920
rect 15212 15966 15332 15994
rect 15016 15904 15068 15910
rect 15016 15846 15068 15852
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 15028 14346 15056 15846
rect 15120 15473 15148 15914
rect 15106 15464 15162 15473
rect 15106 15399 15162 15408
rect 15108 14884 15160 14890
rect 15108 14826 15160 14832
rect 15016 14340 15068 14346
rect 15016 14282 15068 14288
rect 15120 14006 15148 14826
rect 15108 14000 15160 14006
rect 15108 13942 15160 13948
rect 15212 13954 15240 15966
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15304 15745 15332 15846
rect 15290 15736 15346 15745
rect 15290 15671 15346 15680
rect 15396 15620 15424 18550
rect 15488 18426 15516 18634
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15580 16289 15608 19230
rect 15672 17184 15700 20839
rect 15764 18193 15792 27474
rect 15844 26580 15896 26586
rect 15844 26522 15896 26528
rect 15856 22094 15884 26522
rect 16120 26376 16172 26382
rect 16684 26353 16712 29106
rect 16120 26318 16172 26324
rect 16670 26344 16726 26353
rect 16132 25362 16160 26318
rect 16670 26279 16726 26288
rect 16580 26240 16632 26246
rect 16580 26182 16632 26188
rect 16304 25832 16356 25838
rect 16304 25774 16356 25780
rect 16316 25362 16344 25774
rect 16120 25356 16172 25362
rect 16120 25298 16172 25304
rect 16304 25356 16356 25362
rect 16304 25298 16356 25304
rect 16592 25226 16620 26182
rect 16580 25220 16632 25226
rect 16580 25162 16632 25168
rect 16212 24744 16264 24750
rect 16212 24686 16264 24692
rect 16028 22636 16080 22642
rect 16028 22578 16080 22584
rect 15856 22066 15976 22094
rect 15948 21622 15976 22066
rect 15936 21616 15988 21622
rect 15936 21558 15988 21564
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15856 21146 15884 21490
rect 15844 21140 15896 21146
rect 15844 21082 15896 21088
rect 15936 20596 15988 20602
rect 15936 20538 15988 20544
rect 15842 19544 15898 19553
rect 15842 19479 15898 19488
rect 15856 18834 15884 19479
rect 15844 18828 15896 18834
rect 15844 18770 15896 18776
rect 15750 18184 15806 18193
rect 15750 18119 15806 18128
rect 15672 17156 15884 17184
rect 15660 17060 15712 17066
rect 15660 17002 15712 17008
rect 15672 16794 15700 17002
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 15566 16280 15622 16289
rect 15566 16215 15622 16224
rect 15476 15632 15528 15638
rect 15396 15592 15476 15620
rect 15476 15574 15528 15580
rect 15292 15428 15344 15434
rect 15292 15370 15344 15376
rect 15304 15162 15332 15370
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 14832 13252 14884 13258
rect 14660 13212 14832 13240
rect 14660 12345 14688 13212
rect 14832 13194 14884 13200
rect 14830 13152 14886 13161
rect 14830 13087 14886 13096
rect 14844 12850 14872 13087
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 14646 12336 14702 12345
rect 14556 12300 14608 12306
rect 14646 12271 14702 12280
rect 14556 12242 14608 12248
rect 14554 12200 14610 12209
rect 14554 12135 14556 12144
rect 14608 12135 14610 12144
rect 14556 12106 14608 12112
rect 14568 11354 14596 12106
rect 14844 11830 14872 12786
rect 15120 12594 15148 13942
rect 15212 13926 15332 13954
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15028 12566 15148 12594
rect 15028 12434 15056 12566
rect 14936 12406 15056 12434
rect 14832 11824 14884 11830
rect 14832 11766 14884 11772
rect 14648 11620 14700 11626
rect 14648 11562 14700 11568
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14660 11121 14688 11562
rect 14646 11112 14702 11121
rect 14646 11047 14702 11056
rect 14372 9920 14424 9926
rect 14372 9862 14424 9868
rect 14464 9920 14516 9926
rect 14936 9897 14964 12406
rect 15014 10840 15070 10849
rect 15014 10775 15070 10784
rect 15028 10606 15056 10775
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 15028 10169 15056 10542
rect 15212 10180 15240 13806
rect 15304 12850 15332 13926
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15488 12918 15516 13262
rect 15672 12918 15700 16730
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15764 12434 15792 16594
rect 15856 15144 15884 17156
rect 15948 16658 15976 20538
rect 16040 17921 16068 22578
rect 16120 22228 16172 22234
rect 16120 22170 16172 22176
rect 16026 17912 16082 17921
rect 16026 17847 16082 17856
rect 16132 17814 16160 22170
rect 16224 19854 16252 24686
rect 16488 24336 16540 24342
rect 16488 24278 16540 24284
rect 16396 24132 16448 24138
rect 16396 24074 16448 24080
rect 16408 23526 16436 24074
rect 16396 23520 16448 23526
rect 16396 23462 16448 23468
rect 16500 23254 16528 24278
rect 16580 24064 16632 24070
rect 16580 24006 16632 24012
rect 16592 23798 16620 24006
rect 16580 23792 16632 23798
rect 16580 23734 16632 23740
rect 16776 23254 16804 29650
rect 16868 29306 16896 36722
rect 17408 33856 17460 33862
rect 17408 33798 17460 33804
rect 17224 32020 17276 32026
rect 17224 31962 17276 31968
rect 16856 29300 16908 29306
rect 16856 29242 16908 29248
rect 16856 28688 16908 28694
rect 16856 28630 16908 28636
rect 16868 26790 16896 28630
rect 16948 28552 17000 28558
rect 16948 28494 17000 28500
rect 16960 28218 16988 28494
rect 16948 28212 17000 28218
rect 16948 28154 17000 28160
rect 16948 28008 17000 28014
rect 16948 27950 17000 27956
rect 16856 26784 16908 26790
rect 16856 26726 16908 26732
rect 16960 25362 16988 27950
rect 17040 27872 17092 27878
rect 17040 27814 17092 27820
rect 17052 27062 17080 27814
rect 17040 27056 17092 27062
rect 17040 26998 17092 27004
rect 16948 25356 17000 25362
rect 16948 25298 17000 25304
rect 16960 24818 16988 25298
rect 16948 24812 17000 24818
rect 16948 24754 17000 24760
rect 16488 23248 16540 23254
rect 16488 23190 16540 23196
rect 16764 23248 16816 23254
rect 16764 23190 16816 23196
rect 16580 23044 16632 23050
rect 16580 22986 16632 22992
rect 16304 21684 16356 21690
rect 16304 21626 16356 21632
rect 16316 21350 16344 21626
rect 16304 21344 16356 21350
rect 16304 21286 16356 21292
rect 16316 20534 16344 21286
rect 16592 21078 16620 22986
rect 17236 22094 17264 31962
rect 17316 23520 17368 23526
rect 17316 23462 17368 23468
rect 17328 23254 17356 23462
rect 17420 23322 17448 33798
rect 17592 31136 17644 31142
rect 17592 31078 17644 31084
rect 17500 28960 17552 28966
rect 17500 28902 17552 28908
rect 17512 28626 17540 28902
rect 17500 28620 17552 28626
rect 17500 28562 17552 28568
rect 17500 28416 17552 28422
rect 17500 28358 17552 28364
rect 17512 27538 17540 28358
rect 17500 27532 17552 27538
rect 17500 27474 17552 27480
rect 17500 27124 17552 27130
rect 17500 27066 17552 27072
rect 17408 23316 17460 23322
rect 17408 23258 17460 23264
rect 17316 23248 17368 23254
rect 17316 23190 17368 23196
rect 17328 22574 17356 23190
rect 17316 22568 17368 22574
rect 17316 22510 17368 22516
rect 17512 22386 17540 27066
rect 17604 24750 17632 31078
rect 17960 29640 18012 29646
rect 17960 29582 18012 29588
rect 17684 29504 17736 29510
rect 17684 29446 17736 29452
rect 17696 29170 17724 29446
rect 17684 29164 17736 29170
rect 17684 29106 17736 29112
rect 17684 28076 17736 28082
rect 17684 28018 17736 28024
rect 17696 27985 17724 28018
rect 17682 27976 17738 27985
rect 17682 27911 17738 27920
rect 17696 27674 17724 27911
rect 17868 27872 17920 27878
rect 17868 27814 17920 27820
rect 17684 27668 17736 27674
rect 17684 27610 17736 27616
rect 17776 26240 17828 26246
rect 17776 26182 17828 26188
rect 17788 25974 17816 26182
rect 17880 25974 17908 27814
rect 17972 27062 18000 29582
rect 18144 27328 18196 27334
rect 18144 27270 18196 27276
rect 17960 27056 18012 27062
rect 17960 26998 18012 27004
rect 17776 25968 17828 25974
rect 17776 25910 17828 25916
rect 17868 25968 17920 25974
rect 17868 25910 17920 25916
rect 17972 25838 18000 26998
rect 18156 26926 18184 27270
rect 18144 26920 18196 26926
rect 18144 26862 18196 26868
rect 17960 25832 18012 25838
rect 17960 25774 18012 25780
rect 17960 25152 18012 25158
rect 17960 25094 18012 25100
rect 17972 24886 18000 25094
rect 17960 24880 18012 24886
rect 17960 24822 18012 24828
rect 17592 24744 17644 24750
rect 17592 24686 17644 24692
rect 17868 24744 17920 24750
rect 17868 24686 17920 24692
rect 17776 24132 17828 24138
rect 17776 24074 17828 24080
rect 17592 23112 17644 23118
rect 17592 23054 17644 23060
rect 17144 22066 17264 22094
rect 17328 22358 17540 22386
rect 16580 21072 16632 21078
rect 16580 21014 16632 21020
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16948 20936 17000 20942
rect 16948 20878 17000 20884
rect 16304 20528 16356 20534
rect 16304 20470 16356 20476
rect 16396 20528 16448 20534
rect 16396 20470 16448 20476
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 16210 19000 16266 19009
rect 16210 18935 16266 18944
rect 16224 18766 16252 18935
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 16224 18358 16252 18702
rect 16212 18352 16264 18358
rect 16212 18294 16264 18300
rect 16120 17808 16172 17814
rect 16120 17750 16172 17756
rect 16212 17604 16264 17610
rect 16212 17546 16264 17552
rect 16304 17604 16356 17610
rect 16304 17546 16356 17552
rect 16118 17504 16174 17513
rect 16118 17439 16174 17448
rect 16132 16998 16160 17439
rect 16224 17338 16252 17546
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16120 16992 16172 16998
rect 16120 16934 16172 16940
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 15948 15881 15976 16390
rect 15934 15872 15990 15881
rect 15934 15807 15990 15816
rect 15856 15116 15976 15144
rect 15844 15020 15896 15026
rect 15844 14962 15896 14968
rect 15580 12406 15792 12434
rect 15580 12102 15608 12406
rect 15660 12368 15712 12374
rect 15660 12310 15712 12316
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15580 11354 15608 12038
rect 15672 11830 15700 12310
rect 15856 11937 15884 14962
rect 15948 13870 15976 15116
rect 16026 14648 16082 14657
rect 16026 14583 16028 14592
rect 16080 14583 16082 14592
rect 16028 14554 16080 14560
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 15948 12646 15976 13806
rect 16132 13802 16160 16934
rect 16316 16794 16344 17546
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16212 16584 16264 16590
rect 16212 16526 16264 16532
rect 16224 13802 16252 16526
rect 16304 16516 16356 16522
rect 16304 16458 16356 16464
rect 16316 16425 16344 16458
rect 16302 16416 16358 16425
rect 16302 16351 16358 16360
rect 16408 16250 16436 20470
rect 16592 19904 16620 20878
rect 16672 20800 16724 20806
rect 16672 20742 16724 20748
rect 16684 20330 16712 20742
rect 16672 20324 16724 20330
rect 16672 20266 16724 20272
rect 16500 19876 16620 19904
rect 16500 19786 16528 19876
rect 16488 19780 16540 19786
rect 16488 19722 16540 19728
rect 16580 19780 16632 19786
rect 16580 19722 16632 19728
rect 16592 19334 16620 19722
rect 16684 19378 16712 20266
rect 16856 20256 16908 20262
rect 16856 20198 16908 20204
rect 16764 19712 16816 19718
rect 16764 19654 16816 19660
rect 16500 19306 16620 19334
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16500 18290 16528 19306
rect 16672 18760 16724 18766
rect 16672 18702 16724 18708
rect 16488 18284 16540 18290
rect 16488 18226 16540 18232
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 16500 17338 16528 18226
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 16488 16992 16540 16998
rect 16488 16934 16540 16940
rect 16396 16244 16448 16250
rect 16396 16186 16448 16192
rect 16304 15632 16356 15638
rect 16304 15574 16356 15580
rect 16120 13796 16172 13802
rect 16120 13738 16172 13744
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 15842 11928 15898 11937
rect 15842 11863 15898 11872
rect 16040 11830 16068 13670
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16132 12102 16160 12718
rect 16212 12708 16264 12714
rect 16212 12650 16264 12656
rect 16224 12442 16252 12650
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16316 11830 16344 15574
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16408 15473 16436 15506
rect 16394 15464 16450 15473
rect 16394 15399 16450 15408
rect 16500 14804 16528 16934
rect 16592 15978 16620 18226
rect 16684 17513 16712 18702
rect 16670 17504 16726 17513
rect 16670 17439 16726 17448
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16684 16590 16712 17274
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16580 15972 16632 15978
rect 16580 15914 16632 15920
rect 16592 15570 16620 15914
rect 16580 15564 16632 15570
rect 16580 15506 16632 15512
rect 16684 15434 16712 16526
rect 16672 15428 16724 15434
rect 16672 15370 16724 15376
rect 16408 14776 16528 14804
rect 15660 11824 15712 11830
rect 15660 11766 15712 11772
rect 16028 11824 16080 11830
rect 16028 11766 16080 11772
rect 16304 11824 16356 11830
rect 16304 11766 16356 11772
rect 15660 11688 15712 11694
rect 15658 11656 15660 11665
rect 15712 11656 15714 11665
rect 15658 11591 15714 11600
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15752 11280 15804 11286
rect 15752 11222 15804 11228
rect 15660 10736 15712 10742
rect 15660 10678 15712 10684
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15474 10432 15530 10441
rect 15474 10367 15530 10376
rect 15014 10160 15070 10169
rect 15212 10152 15424 10180
rect 15014 10095 15070 10104
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 14464 9862 14516 9868
rect 14922 9888 14978 9897
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 14384 9674 14412 9862
rect 14922 9823 14978 9832
rect 15198 9752 15254 9761
rect 15198 9687 15254 9696
rect 14384 9646 14596 9674
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13740 7342 13768 7822
rect 13820 7472 13872 7478
rect 13820 7414 13872 7420
rect 13636 7336 13688 7342
rect 13636 7278 13688 7284
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 13452 6248 13504 6254
rect 13452 6190 13504 6196
rect 13464 5778 13492 6190
rect 13452 5772 13504 5778
rect 13452 5714 13504 5720
rect 12622 5672 12678 5681
rect 12256 5636 12308 5642
rect 12678 5630 13032 5658
rect 13464 5642 13492 5714
rect 12622 5607 12678 5616
rect 12256 5578 12308 5584
rect 12164 5160 12216 5166
rect 12164 5102 12216 5108
rect 12176 4554 12204 5102
rect 12164 4548 12216 4554
rect 12164 4490 12216 4496
rect 12070 4040 12126 4049
rect 12070 3975 12072 3984
rect 12124 3975 12126 3984
rect 12164 4004 12216 4010
rect 12072 3946 12124 3952
rect 12164 3946 12216 3952
rect 12176 3641 12204 3946
rect 12268 3777 12296 5578
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 13004 4026 13032 5630
rect 13452 5636 13504 5642
rect 13452 5578 13504 5584
rect 13268 5568 13320 5574
rect 13268 5510 13320 5516
rect 13176 5092 13228 5098
rect 13176 5034 13228 5040
rect 13188 4486 13216 5034
rect 13280 5001 13308 5510
rect 13360 5296 13412 5302
rect 13464 5284 13492 5578
rect 13412 5256 13492 5284
rect 13360 5238 13412 5244
rect 13266 4992 13322 5001
rect 13266 4927 13322 4936
rect 13280 4826 13308 4927
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 13360 4752 13412 4758
rect 13360 4694 13412 4700
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13372 4026 13400 4694
rect 13648 4554 13676 7278
rect 13740 6798 13768 7278
rect 13832 7002 13860 7414
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13740 6390 13768 6734
rect 13728 6384 13780 6390
rect 13728 6326 13780 6332
rect 13820 6384 13872 6390
rect 13820 6326 13872 6332
rect 13728 5296 13780 5302
rect 13728 5238 13780 5244
rect 13740 4622 13768 5238
rect 13832 4729 13860 6326
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 13910 5400 13966 5409
rect 13910 5335 13966 5344
rect 13818 4720 13874 4729
rect 13818 4655 13874 4664
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13636 4548 13688 4554
rect 13636 4490 13688 4496
rect 13452 4208 13504 4214
rect 13740 4162 13768 4558
rect 13818 4312 13874 4321
rect 13818 4247 13874 4256
rect 13832 4214 13860 4247
rect 13504 4156 13768 4162
rect 13452 4150 13768 4156
rect 13820 4208 13872 4214
rect 13820 4150 13872 4156
rect 13464 4134 13768 4150
rect 13542 4040 13598 4049
rect 12254 3768 12310 3777
rect 12254 3703 12310 3712
rect 12544 3670 12572 4014
rect 13004 3998 13124 4026
rect 13372 3998 13492 4026
rect 12624 3936 12676 3942
rect 12992 3936 13044 3942
rect 12676 3896 12940 3924
rect 12624 3878 12676 3884
rect 12532 3664 12584 3670
rect 12162 3632 12218 3641
rect 12532 3606 12584 3612
rect 12162 3567 12218 3576
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 12164 3052 12216 3058
rect 12164 2994 12216 3000
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 10966 2343 11022 2352
rect 11520 2372 11572 2378
rect 11520 2314 11572 2320
rect 11612 2372 11664 2378
rect 11612 2314 11664 2320
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 10600 1828 10652 1834
rect 10600 1770 10652 1776
rect 10414 1728 10470 1737
rect 10414 1663 10470 1672
rect 10980 800 11008 2246
rect 11624 800 11652 2314
rect 11992 2106 12020 2586
rect 12176 2378 12204 2994
rect 12164 2372 12216 2378
rect 12164 2314 12216 2320
rect 11980 2100 12032 2106
rect 11980 2042 12032 2048
rect 12532 1896 12584 1902
rect 12532 1838 12584 1844
rect 12544 1698 12572 1838
rect 12532 1692 12584 1698
rect 12532 1634 12584 1640
rect 12912 800 12940 3896
rect 12990 3904 12992 3913
rect 13044 3904 13046 3913
rect 12990 3839 13046 3848
rect 13096 3534 13124 3998
rect 13464 3738 13492 3998
rect 13542 3975 13598 3984
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 13372 3534 13400 3674
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13464 3126 13492 3674
rect 13556 3466 13584 3975
rect 13740 3602 13768 4134
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13544 3460 13596 3466
rect 13544 3402 13596 3408
rect 13648 3369 13676 3538
rect 13634 3360 13690 3369
rect 13634 3295 13690 3304
rect 13360 3120 13412 3126
rect 13360 3062 13412 3068
rect 13452 3120 13504 3126
rect 13452 3062 13504 3068
rect 13372 2938 13400 3062
rect 13740 2938 13768 3538
rect 13372 2910 13768 2938
rect 13450 2680 13506 2689
rect 13450 2615 13506 2624
rect 13464 2446 13492 2615
rect 13740 2514 13768 2910
rect 13924 2582 13952 5335
rect 14108 5166 14136 5510
rect 14200 5166 14228 9454
rect 14476 8906 14504 9454
rect 14464 8900 14516 8906
rect 14464 8842 14516 8848
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 14292 7342 14320 8230
rect 14568 7750 14596 9646
rect 14922 9344 14978 9353
rect 14922 9279 14978 9288
rect 14832 8900 14884 8906
rect 14832 8842 14884 8848
rect 14844 8809 14872 8842
rect 14830 8800 14886 8809
rect 14830 8735 14886 8744
rect 14936 8294 14964 9279
rect 15212 8294 15240 9687
rect 15304 9178 15332 9930
rect 15396 9364 15424 10152
rect 15488 9654 15516 10367
rect 15580 10198 15608 10474
rect 15568 10192 15620 10198
rect 15568 10134 15620 10140
rect 15476 9648 15528 9654
rect 15476 9590 15528 9596
rect 15568 9376 15620 9382
rect 15396 9336 15568 9364
rect 15568 9318 15620 9324
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15580 9042 15608 9318
rect 15568 9036 15620 9042
rect 15568 8978 15620 8984
rect 15568 8560 15620 8566
rect 15474 8528 15530 8537
rect 15568 8502 15620 8508
rect 15474 8463 15476 8472
rect 15528 8463 15530 8472
rect 15476 8434 15528 8440
rect 14924 8288 14976 8294
rect 15200 8288 15252 8294
rect 14924 8230 14976 8236
rect 15106 8256 15162 8265
rect 15200 8230 15252 8236
rect 15106 8191 15162 8200
rect 14832 7812 14884 7818
rect 14832 7754 14884 7760
rect 14556 7744 14608 7750
rect 14844 7721 14872 7754
rect 14556 7686 14608 7692
rect 14830 7712 14886 7721
rect 14830 7647 14886 7656
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 14556 5636 14608 5642
rect 14556 5578 14608 5584
rect 14096 5160 14148 5166
rect 14096 5102 14148 5108
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14200 4690 14228 4966
rect 14188 4684 14240 4690
rect 14188 4626 14240 4632
rect 14004 4208 14056 4214
rect 14004 4150 14056 4156
rect 14016 2990 14044 4150
rect 14568 4010 14596 5578
rect 15120 4321 15148 8191
rect 15580 7274 15608 8502
rect 15568 7268 15620 7274
rect 15568 7210 15620 7216
rect 15290 6896 15346 6905
rect 15290 6831 15346 6840
rect 15568 6860 15620 6866
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 15212 5098 15240 6190
rect 15200 5092 15252 5098
rect 15200 5034 15252 5040
rect 15106 4312 15162 4321
rect 15106 4247 15162 4256
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 14556 4004 14608 4010
rect 14556 3946 14608 3952
rect 14844 3754 14872 4082
rect 14200 3726 14872 3754
rect 14200 3670 14228 3726
rect 14188 3664 14240 3670
rect 14188 3606 14240 3612
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14844 3097 14872 3402
rect 14830 3088 14886 3097
rect 14830 3023 14886 3032
rect 14004 2984 14056 2990
rect 14004 2926 14056 2932
rect 15120 2854 15148 4247
rect 15200 4072 15252 4078
rect 15200 4014 15252 4020
rect 15212 3754 15240 4014
rect 15304 3913 15332 6831
rect 15672 6848 15700 10678
rect 15764 8809 15792 11222
rect 15934 10840 15990 10849
rect 15934 10775 15990 10784
rect 15842 10024 15898 10033
rect 15842 9959 15844 9968
rect 15896 9959 15898 9968
rect 15844 9930 15896 9936
rect 15844 9648 15896 9654
rect 15844 9590 15896 9596
rect 15856 9110 15884 9590
rect 15844 9104 15896 9110
rect 15844 9046 15896 9052
rect 15844 8900 15896 8906
rect 15844 8842 15896 8848
rect 15750 8800 15806 8809
rect 15750 8735 15806 8744
rect 15764 7342 15792 8735
rect 15752 7336 15804 7342
rect 15752 7278 15804 7284
rect 15620 6820 15700 6848
rect 15568 6802 15620 6808
rect 15856 6769 15884 8842
rect 15948 7002 15976 10775
rect 16408 10656 16436 14776
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 16684 13938 16712 14214
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16132 10628 16436 10656
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 16040 9178 16068 9522
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 16132 8362 16160 10628
rect 16394 10296 16450 10305
rect 16394 10231 16450 10240
rect 16302 9616 16358 9625
rect 16302 9551 16304 9560
rect 16356 9551 16358 9560
rect 16304 9522 16356 9528
rect 16304 8560 16356 8566
rect 16224 8520 16304 8548
rect 16120 8356 16172 8362
rect 16120 8298 16172 8304
rect 16028 8288 16080 8294
rect 16028 8230 16080 8236
rect 16040 7970 16068 8230
rect 16132 8090 16160 8298
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 16040 7942 16160 7970
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 15658 6760 15714 6769
rect 15658 6695 15714 6704
rect 15842 6760 15898 6769
rect 15842 6695 15898 6704
rect 15672 6361 15700 6695
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15658 6352 15714 6361
rect 15658 6287 15714 6296
rect 15660 6248 15712 6254
rect 15660 6190 15712 6196
rect 15384 6180 15436 6186
rect 15384 6122 15436 6128
rect 15290 3904 15346 3913
rect 15290 3839 15346 3848
rect 15396 3754 15424 6122
rect 15672 6089 15700 6190
rect 15658 6080 15714 6089
rect 15658 6015 15714 6024
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15488 4146 15516 5102
rect 15568 4548 15620 4554
rect 15568 4490 15620 4496
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 15212 3726 15424 3754
rect 15476 3120 15528 3126
rect 15476 3062 15528 3068
rect 15108 2848 15160 2854
rect 14186 2816 14242 2825
rect 15488 2825 15516 3062
rect 15108 2790 15160 2796
rect 15474 2816 15530 2825
rect 14186 2751 14242 2760
rect 15474 2751 15530 2760
rect 13912 2576 13964 2582
rect 13912 2518 13964 2524
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 13452 2440 13504 2446
rect 13452 2382 13504 2388
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 13556 1630 13584 2246
rect 13544 1624 13596 1630
rect 13544 1566 13596 1572
rect 14200 800 14228 2751
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 14464 1964 14516 1970
rect 14464 1906 14516 1912
rect 14476 1766 14504 1906
rect 14464 1760 14516 1766
rect 14464 1702 14516 1708
rect 14844 800 14872 2246
rect 15580 2038 15608 4490
rect 15568 2032 15620 2038
rect 15568 1974 15620 1980
rect 15672 1698 15700 5646
rect 15764 5386 15792 6394
rect 15948 6118 15976 6938
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 15764 5358 15884 5386
rect 15752 5296 15804 5302
rect 15752 5238 15804 5244
rect 15764 5137 15792 5238
rect 15750 5128 15806 5137
rect 15750 5063 15806 5072
rect 15856 4729 15884 5358
rect 16040 4758 16068 5714
rect 16028 4752 16080 4758
rect 15842 4720 15898 4729
rect 16028 4694 16080 4700
rect 15842 4655 15898 4664
rect 16040 4321 16068 4694
rect 16026 4312 16082 4321
rect 16026 4247 16082 4256
rect 16132 4010 16160 7942
rect 16224 4146 16252 8520
rect 16304 8502 16356 8508
rect 16408 8430 16436 10231
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16396 7948 16448 7954
rect 16500 7936 16528 13466
rect 16776 13326 16804 19654
rect 16868 19242 16896 20198
rect 16856 19236 16908 19242
rect 16856 19178 16908 19184
rect 16960 18766 16988 20878
rect 17040 19712 17092 19718
rect 17040 19654 17092 19660
rect 17052 19446 17080 19654
rect 17040 19440 17092 19446
rect 17040 19382 17092 19388
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 17052 18465 17080 18566
rect 17038 18456 17094 18465
rect 17038 18391 17094 18400
rect 17040 18352 17092 18358
rect 17040 18294 17092 18300
rect 16856 17264 16908 17270
rect 16856 17206 16908 17212
rect 16868 14006 16896 17206
rect 16948 17060 17000 17066
rect 16948 17002 17000 17008
rect 16960 16590 16988 17002
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16948 15428 17000 15434
rect 16948 15370 17000 15376
rect 16960 14074 16988 15370
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 16856 14000 16908 14006
rect 16856 13942 16908 13948
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 16672 13184 16724 13190
rect 16672 13126 16724 13132
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16592 12345 16620 12378
rect 16578 12336 16634 12345
rect 16578 12271 16634 12280
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16592 11898 16620 12106
rect 16580 11892 16632 11898
rect 16580 11834 16632 11840
rect 16580 11688 16632 11694
rect 16580 11630 16632 11636
rect 16592 10033 16620 11630
rect 16684 10062 16712 13126
rect 16960 12850 16988 13262
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 16764 12096 16816 12102
rect 16764 12038 16816 12044
rect 16776 11830 16804 12038
rect 16764 11824 16816 11830
rect 16764 11766 16816 11772
rect 16764 10464 16816 10470
rect 16764 10406 16816 10412
rect 16672 10056 16724 10062
rect 16578 10024 16634 10033
rect 16672 9998 16724 10004
rect 16578 9959 16634 9968
rect 16448 7908 16528 7936
rect 16396 7890 16448 7896
rect 16396 7812 16448 7818
rect 16396 7754 16448 7760
rect 16408 7002 16436 7754
rect 16396 6996 16448 7002
rect 16396 6938 16448 6944
rect 16500 6934 16528 7908
rect 16670 7848 16726 7857
rect 16670 7783 16672 7792
rect 16724 7783 16726 7792
rect 16672 7754 16724 7760
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16488 6928 16540 6934
rect 16488 6870 16540 6876
rect 16592 6730 16620 7142
rect 16580 6724 16632 6730
rect 16580 6666 16632 6672
rect 16486 6216 16542 6225
rect 16486 6151 16542 6160
rect 16304 6112 16356 6118
rect 16304 6054 16356 6060
rect 16316 5914 16344 6054
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 16500 5166 16528 6151
rect 16776 5760 16804 10406
rect 16868 9042 16896 12378
rect 16960 11914 16988 12786
rect 17052 12306 17080 18294
rect 17144 17610 17172 22066
rect 17328 21486 17356 22358
rect 17500 22228 17552 22234
rect 17500 22170 17552 22176
rect 17512 21622 17540 22170
rect 17604 21706 17632 23054
rect 17684 23044 17736 23050
rect 17684 22986 17736 22992
rect 17696 22545 17724 22986
rect 17682 22536 17738 22545
rect 17682 22471 17738 22480
rect 17604 21678 17724 21706
rect 17500 21616 17552 21622
rect 17500 21558 17552 21564
rect 17592 21616 17644 21622
rect 17592 21558 17644 21564
rect 17316 21480 17368 21486
rect 17316 21422 17368 21428
rect 17328 20398 17356 21422
rect 17604 21146 17632 21558
rect 17696 21486 17724 21678
rect 17684 21480 17736 21486
rect 17684 21422 17736 21428
rect 17592 21140 17644 21146
rect 17592 21082 17644 21088
rect 17696 21026 17724 21422
rect 17604 20998 17724 21026
rect 17316 20392 17368 20398
rect 17316 20334 17368 20340
rect 17604 20330 17632 20998
rect 17408 20324 17460 20330
rect 17408 20266 17460 20272
rect 17592 20324 17644 20330
rect 17592 20266 17644 20272
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 17236 20058 17264 20198
rect 17420 20058 17448 20266
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 17408 19508 17460 19514
rect 17408 19450 17460 19456
rect 17316 19304 17368 19310
rect 17316 19246 17368 19252
rect 17224 19168 17276 19174
rect 17224 19110 17276 19116
rect 17236 18698 17264 19110
rect 17224 18692 17276 18698
rect 17224 18634 17276 18640
rect 17328 17762 17356 19246
rect 17420 18630 17448 19450
rect 17408 18624 17460 18630
rect 17408 18566 17460 18572
rect 17236 17734 17356 17762
rect 17132 17604 17184 17610
rect 17132 17546 17184 17552
rect 17130 13696 17186 13705
rect 17130 13631 17186 13640
rect 17144 12918 17172 13631
rect 17132 12912 17184 12918
rect 17132 12854 17184 12860
rect 17236 12753 17264 17734
rect 17316 17672 17368 17678
rect 17314 17640 17316 17649
rect 17368 17640 17370 17649
rect 17314 17575 17370 17584
rect 17314 17232 17370 17241
rect 17314 17167 17370 17176
rect 17328 17134 17356 17167
rect 17316 17128 17368 17134
rect 17316 17070 17368 17076
rect 17316 16108 17368 16114
rect 17316 16050 17368 16056
rect 17328 15502 17356 16050
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 17328 13326 17356 15438
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17316 12912 17368 12918
rect 17314 12880 17316 12889
rect 17368 12880 17370 12889
rect 17314 12815 17370 12824
rect 17316 12776 17368 12782
rect 17222 12744 17278 12753
rect 17316 12718 17368 12724
rect 17222 12679 17278 12688
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 17224 12164 17276 12170
rect 17224 12106 17276 12112
rect 16960 11886 17080 11914
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 16960 10985 16988 11766
rect 17052 11694 17080 11886
rect 17040 11688 17092 11694
rect 17040 11630 17092 11636
rect 17038 11520 17094 11529
rect 17038 11455 17094 11464
rect 17052 11098 17080 11455
rect 17052 11070 17172 11098
rect 17040 11008 17092 11014
rect 16946 10976 17002 10985
rect 17040 10950 17092 10956
rect 16946 10911 17002 10920
rect 17052 10826 17080 10950
rect 16960 10798 17080 10826
rect 16960 10674 16988 10798
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 17144 9330 17172 11070
rect 17236 10470 17264 12106
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 17236 9722 17264 9862
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17328 9466 17356 12718
rect 17420 9586 17448 18566
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 17512 17202 17540 17614
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17512 16697 17540 17138
rect 17498 16688 17554 16697
rect 17498 16623 17554 16632
rect 17512 16590 17540 16623
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17604 14958 17632 20266
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 17696 18086 17724 18906
rect 17684 18080 17736 18086
rect 17684 18022 17736 18028
rect 17684 17604 17736 17610
rect 17684 17546 17736 17552
rect 17696 17377 17724 17546
rect 17682 17368 17738 17377
rect 17682 17303 17738 17312
rect 17788 17270 17816 24074
rect 17880 22234 17908 24686
rect 17960 24676 18012 24682
rect 17960 24618 18012 24624
rect 17868 22228 17920 22234
rect 17868 22170 17920 22176
rect 17972 22166 18000 24618
rect 18524 24206 18552 37266
rect 18708 37262 18736 39200
rect 18696 37256 18748 37262
rect 18696 37198 18748 37204
rect 19064 37188 19116 37194
rect 19064 37130 19116 37136
rect 18788 32020 18840 32026
rect 18788 31962 18840 31968
rect 18800 31754 18828 31962
rect 18616 31726 18828 31754
rect 18420 24200 18472 24206
rect 18420 24142 18472 24148
rect 18512 24200 18564 24206
rect 18512 24142 18564 24148
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 17960 22160 18012 22166
rect 17960 22102 18012 22108
rect 18064 21486 18092 23598
rect 18328 23112 18380 23118
rect 18328 23054 18380 23060
rect 18144 23044 18196 23050
rect 18144 22986 18196 22992
rect 18156 22137 18184 22986
rect 18340 22273 18368 23054
rect 18326 22264 18382 22273
rect 18326 22199 18382 22208
rect 18142 22128 18198 22137
rect 18142 22063 18198 22072
rect 18144 21956 18196 21962
rect 18144 21898 18196 21904
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 18050 21040 18106 21049
rect 18050 20975 18106 20984
rect 17960 20868 18012 20874
rect 17960 20810 18012 20816
rect 17972 20369 18000 20810
rect 17958 20360 18014 20369
rect 17958 20295 18014 20304
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 17972 18766 18000 19110
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 17776 17264 17828 17270
rect 17776 17206 17828 17212
rect 18064 17082 18092 20975
rect 18156 20398 18184 21898
rect 18326 21720 18382 21729
rect 18326 21655 18382 21664
rect 18144 20392 18196 20398
rect 18144 20334 18196 20340
rect 18156 19281 18184 20334
rect 18234 19680 18290 19689
rect 18234 19615 18290 19624
rect 18142 19272 18198 19281
rect 18142 19207 18198 19216
rect 18144 18760 18196 18766
rect 18142 18728 18144 18737
rect 18196 18728 18198 18737
rect 18142 18663 18198 18672
rect 17972 17054 18092 17082
rect 17868 16720 17920 16726
rect 17868 16662 17920 16668
rect 17682 15328 17738 15337
rect 17682 15263 17738 15272
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 17590 14784 17646 14793
rect 17590 14719 17646 14728
rect 17604 12918 17632 14719
rect 17696 14006 17724 15263
rect 17880 14958 17908 16662
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17776 14816 17828 14822
rect 17880 14793 17908 14894
rect 17776 14758 17828 14764
rect 17866 14784 17922 14793
rect 17788 14346 17816 14758
rect 17866 14719 17922 14728
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 17776 14340 17828 14346
rect 17776 14282 17828 14288
rect 17684 14000 17736 14006
rect 17684 13942 17736 13948
rect 17696 13841 17724 13942
rect 17776 13864 17828 13870
rect 17682 13832 17738 13841
rect 17776 13806 17828 13812
rect 17682 13767 17738 13776
rect 17788 13138 17816 13806
rect 17696 13110 17816 13138
rect 17592 12912 17644 12918
rect 17592 12854 17644 12860
rect 17590 12744 17646 12753
rect 17590 12679 17646 12688
rect 17604 11830 17632 12679
rect 17592 11824 17644 11830
rect 17592 11766 17644 11772
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17604 9466 17632 10066
rect 17328 9438 17632 9466
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16854 6488 16910 6497
rect 16854 6423 16910 6432
rect 16684 5732 16804 5760
rect 16488 5160 16540 5166
rect 16488 5102 16540 5108
rect 16580 4548 16632 4554
rect 16580 4490 16632 4496
rect 16592 4214 16620 4490
rect 16580 4208 16632 4214
rect 16580 4150 16632 4156
rect 16212 4140 16264 4146
rect 16212 4082 16264 4088
rect 16028 4004 16080 4010
rect 16028 3946 16080 3952
rect 16120 4004 16172 4010
rect 16120 3946 16172 3952
rect 16040 3738 16068 3946
rect 16578 3768 16634 3777
rect 16028 3732 16080 3738
rect 16578 3703 16634 3712
rect 16028 3674 16080 3680
rect 16394 3632 16450 3641
rect 16394 3567 16450 3576
rect 16408 3466 16436 3567
rect 16592 3466 16620 3703
rect 16396 3460 16448 3466
rect 16396 3402 16448 3408
rect 16580 3460 16632 3466
rect 16580 3402 16632 3408
rect 16302 3360 16358 3369
rect 16302 3295 16358 3304
rect 16316 2922 16344 3295
rect 16684 3233 16712 5732
rect 16868 5658 16896 6423
rect 16776 5630 16896 5658
rect 16776 4146 16804 5630
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16856 4072 16908 4078
rect 16856 4014 16908 4020
rect 16868 3602 16896 4014
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16762 3360 16818 3369
rect 16762 3295 16818 3304
rect 16670 3224 16726 3233
rect 16670 3159 16726 3168
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 16304 2916 16356 2922
rect 16304 2858 16356 2864
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 15948 1970 15976 2586
rect 16120 2576 16172 2582
rect 16120 2518 16172 2524
rect 15936 1964 15988 1970
rect 15936 1906 15988 1912
rect 15660 1692 15712 1698
rect 15660 1634 15712 1640
rect 16132 800 16160 2518
rect 16592 2514 16620 3062
rect 16684 3058 16712 3159
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 16776 2650 16804 3295
rect 16764 2644 16816 2650
rect 16764 2586 16816 2592
rect 16580 2508 16632 2514
rect 16580 2450 16632 2456
rect 16764 2372 16816 2378
rect 16764 2314 16816 2320
rect 16776 2038 16804 2314
rect 16764 2032 16816 2038
rect 16764 1974 16816 1980
rect 16960 1698 16988 9318
rect 17144 9302 17356 9330
rect 17224 9104 17276 9110
rect 17038 9072 17094 9081
rect 17224 9046 17276 9052
rect 17038 9007 17094 9016
rect 17052 6202 17080 9007
rect 17236 8634 17264 9046
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17130 8528 17186 8537
rect 17130 8463 17186 8472
rect 17144 6390 17172 8463
rect 17222 8392 17278 8401
rect 17222 8327 17278 8336
rect 17236 7546 17264 8327
rect 17224 7540 17276 7546
rect 17224 7482 17276 7488
rect 17132 6384 17184 6390
rect 17132 6326 17184 6332
rect 17328 6322 17356 9302
rect 17408 9036 17460 9042
rect 17408 8978 17460 8984
rect 17420 8634 17448 8978
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17604 8566 17632 9438
rect 17696 9081 17724 13110
rect 17776 12912 17828 12918
rect 17776 12854 17828 12860
rect 17682 9072 17738 9081
rect 17682 9007 17738 9016
rect 17684 8900 17736 8906
rect 17788 8888 17816 12854
rect 17880 12170 17908 14554
rect 17972 13190 18000 17054
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 18064 15026 18092 15438
rect 18248 15434 18276 19615
rect 18236 15428 18288 15434
rect 18236 15370 18288 15376
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 18052 15020 18104 15026
rect 18052 14962 18104 14968
rect 18156 14498 18184 15302
rect 18156 14470 18276 14498
rect 18144 14340 18196 14346
rect 18144 14282 18196 14288
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 17960 13184 18012 13190
rect 17960 13126 18012 13132
rect 17958 13016 18014 13025
rect 17958 12951 18014 12960
rect 17868 12164 17920 12170
rect 17868 12106 17920 12112
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17880 11150 17908 11630
rect 17972 11218 18000 12951
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17960 10804 18012 10810
rect 18064 10792 18092 14214
rect 18012 10764 18092 10792
rect 17960 10746 18012 10752
rect 17736 8860 17816 8888
rect 17684 8842 17736 8848
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 17696 7478 17724 8842
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17880 8566 17908 8774
rect 17868 8560 17920 8566
rect 17868 8502 17920 8508
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17684 7472 17736 7478
rect 17684 7414 17736 7420
rect 17592 7336 17644 7342
rect 17592 7278 17644 7284
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17052 6174 17172 6202
rect 17040 5296 17092 5302
rect 17040 5238 17092 5244
rect 17052 4826 17080 5238
rect 17040 4820 17092 4826
rect 17040 4762 17092 4768
rect 17144 2774 17172 6174
rect 17224 5296 17276 5302
rect 17224 5238 17276 5244
rect 17236 4758 17264 5238
rect 17224 4752 17276 4758
rect 17224 4694 17276 4700
rect 17236 3777 17264 4694
rect 17222 3768 17278 3777
rect 17222 3703 17278 3712
rect 17328 3369 17356 6258
rect 17420 6186 17448 6734
rect 17408 6180 17460 6186
rect 17408 6122 17460 6128
rect 17604 5778 17632 7278
rect 17684 7268 17736 7274
rect 17684 7210 17736 7216
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 17592 5772 17644 5778
rect 17592 5714 17644 5720
rect 17420 5681 17448 5714
rect 17406 5672 17462 5681
rect 17406 5607 17462 5616
rect 17590 5128 17646 5137
rect 17590 5063 17646 5072
rect 17604 4758 17632 5063
rect 17592 4752 17644 4758
rect 17592 4694 17644 4700
rect 17408 4208 17460 4214
rect 17408 4150 17460 4156
rect 17314 3360 17370 3369
rect 17314 3295 17370 3304
rect 17144 2746 17356 2774
rect 17328 2650 17356 2746
rect 17420 2650 17448 4150
rect 17592 3732 17644 3738
rect 17592 3674 17644 3680
rect 17604 2922 17632 3674
rect 17696 3126 17724 7210
rect 17774 6896 17830 6905
rect 17774 6831 17776 6840
rect 17828 6831 17830 6840
rect 17776 6802 17828 6808
rect 17776 6384 17828 6390
rect 17776 6326 17828 6332
rect 17788 3738 17816 6326
rect 17880 5681 17908 7822
rect 17866 5672 17922 5681
rect 17866 5607 17922 5616
rect 17866 5536 17922 5545
rect 17866 5471 17922 5480
rect 17880 5166 17908 5471
rect 17972 5302 18000 10746
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 18064 9450 18092 9998
rect 18156 9654 18184 14282
rect 18248 13802 18276 14470
rect 18236 13796 18288 13802
rect 18236 13738 18288 13744
rect 18340 12434 18368 21655
rect 18432 19174 18460 24142
rect 18616 23594 18644 31726
rect 18788 27328 18840 27334
rect 18788 27270 18840 27276
rect 18696 24744 18748 24750
rect 18696 24686 18748 24692
rect 18604 23588 18656 23594
rect 18604 23530 18656 23536
rect 18512 23520 18564 23526
rect 18512 23462 18564 23468
rect 18524 22506 18552 23462
rect 18512 22500 18564 22506
rect 18512 22442 18564 22448
rect 18420 19168 18472 19174
rect 18420 19110 18472 19116
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18432 18630 18460 18702
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 18524 16046 18552 22442
rect 18708 21350 18736 24686
rect 18696 21344 18748 21350
rect 18696 21286 18748 21292
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18708 19922 18736 20402
rect 18696 19916 18748 19922
rect 18696 19858 18748 19864
rect 18602 19272 18658 19281
rect 18602 19207 18658 19216
rect 18616 16833 18644 19207
rect 18602 16824 18658 16833
rect 18602 16759 18658 16768
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18512 16040 18564 16046
rect 18512 15982 18564 15988
rect 18420 14884 18472 14890
rect 18420 14826 18472 14832
rect 18432 12918 18460 14826
rect 18420 12912 18472 12918
rect 18420 12854 18472 12860
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 18432 12646 18460 12718
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18340 12406 18460 12434
rect 18432 12170 18460 12406
rect 18420 12164 18472 12170
rect 18420 12106 18472 12112
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 18248 11393 18276 11494
rect 18234 11384 18290 11393
rect 18234 11319 18290 11328
rect 18432 11286 18460 12106
rect 18236 11280 18288 11286
rect 18236 11222 18288 11228
rect 18420 11280 18472 11286
rect 18420 11222 18472 11228
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 18052 9444 18104 9450
rect 18052 9386 18104 9392
rect 18064 8498 18092 9386
rect 18144 8900 18196 8906
rect 18248 8888 18276 11222
rect 18524 11014 18552 15982
rect 18616 14958 18644 16526
rect 18696 16448 18748 16454
rect 18696 16390 18748 16396
rect 18708 16046 18736 16390
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 18696 14952 18748 14958
rect 18696 14894 18748 14900
rect 18708 14550 18736 14894
rect 18800 14822 18828 27270
rect 18880 25696 18932 25702
rect 18880 25638 18932 25644
rect 18892 23662 18920 25638
rect 19076 24410 19104 37130
rect 19996 37126 20024 39200
rect 21284 37330 21312 39200
rect 21272 37324 21324 37330
rect 21272 37266 21324 37272
rect 20076 37256 20128 37262
rect 20076 37198 20128 37204
rect 21456 37256 21508 37262
rect 21456 37198 21508 37204
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19340 36848 19392 36854
rect 19340 36790 19392 36796
rect 19248 28076 19300 28082
rect 19248 28018 19300 28024
rect 19260 27674 19288 28018
rect 19248 27668 19300 27674
rect 19248 27610 19300 27616
rect 19352 27470 19380 36790
rect 20088 36378 20116 37198
rect 20720 36576 20772 36582
rect 20720 36518 20772 36524
rect 20076 36372 20128 36378
rect 20076 36314 20128 36320
rect 19984 36168 20036 36174
rect 19984 36110 20036 36116
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19996 35290 20024 36110
rect 19984 35284 20036 35290
rect 19984 35226 20036 35232
rect 19432 35080 19484 35086
rect 19432 35022 19484 35028
rect 19340 27464 19392 27470
rect 19340 27406 19392 27412
rect 19248 25288 19300 25294
rect 19248 25230 19300 25236
rect 19064 24404 19116 24410
rect 19064 24346 19116 24352
rect 18972 23792 19024 23798
rect 18972 23734 19024 23740
rect 18880 23656 18932 23662
rect 18880 23598 18932 23604
rect 18984 23322 19012 23734
rect 18972 23316 19024 23322
rect 18972 23258 19024 23264
rect 18880 23180 18932 23186
rect 18880 23122 18932 23128
rect 18892 22982 18920 23122
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18892 22574 18920 22918
rect 18880 22568 18932 22574
rect 18880 22510 18932 22516
rect 19156 22568 19208 22574
rect 19156 22510 19208 22516
rect 18880 21480 18932 21486
rect 18880 21422 18932 21428
rect 18892 20058 18920 21422
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 18892 15162 18920 19994
rect 18970 16960 19026 16969
rect 18970 16895 19026 16904
rect 18984 16726 19012 16895
rect 18972 16720 19024 16726
rect 18972 16662 19024 16668
rect 18972 16108 19024 16114
rect 18972 16050 19024 16056
rect 18984 15570 19012 16050
rect 19168 15706 19196 22510
rect 19260 19281 19288 25230
rect 19444 23050 19472 35022
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 20732 32434 20760 36518
rect 21364 33992 21416 33998
rect 21364 33934 21416 33940
rect 20720 32428 20772 32434
rect 20720 32370 20772 32376
rect 20628 32224 20680 32230
rect 20628 32166 20680 32172
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 20352 27396 20404 27402
rect 20352 27338 20404 27344
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 20364 24410 20392 27338
rect 20640 26450 20668 32166
rect 20720 31884 20772 31890
rect 20720 31826 20772 31832
rect 20628 26444 20680 26450
rect 20628 26386 20680 26392
rect 20352 24404 20404 24410
rect 20352 24346 20404 24352
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19432 23044 19484 23050
rect 19432 22986 19484 22992
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 20168 21412 20220 21418
rect 20168 21354 20220 21360
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19352 20466 19380 20878
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19524 20528 19576 20534
rect 19524 20470 19576 20476
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 19536 20346 19564 20470
rect 19536 20330 19748 20346
rect 19536 20324 19760 20330
rect 19536 20318 19708 20324
rect 19708 20266 19760 20272
rect 20180 19854 20208 21354
rect 20168 19848 20220 19854
rect 20168 19790 20220 19796
rect 19984 19780 20036 19786
rect 19984 19722 20036 19728
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19246 19272 19302 19281
rect 19246 19207 19302 19216
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19260 17218 19288 19110
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 18426 20024 19722
rect 20364 19514 20392 24346
rect 20732 21010 20760 31826
rect 21376 28218 21404 33934
rect 21364 28212 21416 28218
rect 21364 28154 21416 28160
rect 20812 26308 20864 26314
rect 20812 26250 20864 26256
rect 20824 25498 20852 26250
rect 20812 25492 20864 25498
rect 20812 25434 20864 25440
rect 20812 25152 20864 25158
rect 20812 25094 20864 25100
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20444 19984 20496 19990
rect 20444 19926 20496 19932
rect 20628 19984 20680 19990
rect 20628 19926 20680 19932
rect 20456 19514 20484 19926
rect 20352 19508 20404 19514
rect 20352 19450 20404 19456
rect 20444 19508 20496 19514
rect 20444 19450 20496 19456
rect 20444 19372 20496 19378
rect 20444 19314 20496 19320
rect 20352 19304 20404 19310
rect 20352 19246 20404 19252
rect 20260 18760 20312 18766
rect 20260 18702 20312 18708
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 20076 18284 20128 18290
rect 20076 18226 20128 18232
rect 19890 17640 19946 17649
rect 19890 17575 19892 17584
rect 19944 17575 19946 17584
rect 19984 17604 20036 17610
rect 19892 17546 19944 17552
rect 19984 17546 20036 17552
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19996 17338 20024 17546
rect 19984 17332 20036 17338
rect 19984 17274 20036 17280
rect 19432 17264 19484 17270
rect 19260 17190 19334 17218
rect 19432 17206 19484 17212
rect 19306 17184 19334 17190
rect 19306 17156 19380 17184
rect 19352 17105 19380 17156
rect 19338 17096 19394 17105
rect 19338 17031 19394 17040
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19352 16674 19380 16934
rect 19260 16646 19380 16674
rect 19156 15700 19208 15706
rect 19156 15642 19208 15648
rect 19260 15638 19288 16646
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19248 15632 19300 15638
rect 19248 15574 19300 15580
rect 18972 15564 19024 15570
rect 18972 15506 19024 15512
rect 19064 15564 19116 15570
rect 19064 15506 19116 15512
rect 18972 15428 19024 15434
rect 18972 15370 19024 15376
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 18788 14816 18840 14822
rect 18788 14758 18840 14764
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18616 12968 18644 14010
rect 18892 13938 18920 14962
rect 18984 14346 19012 15370
rect 18972 14340 19024 14346
rect 18972 14282 19024 14288
rect 18970 14240 19026 14249
rect 18970 14175 19026 14184
rect 18984 13938 19012 14175
rect 18880 13932 18932 13938
rect 18880 13874 18932 13880
rect 18972 13932 19024 13938
rect 18972 13874 19024 13880
rect 18696 13796 18748 13802
rect 18696 13738 18748 13744
rect 18708 13326 18736 13738
rect 18786 13696 18842 13705
rect 18786 13631 18842 13640
rect 18970 13696 19026 13705
rect 18970 13631 19026 13640
rect 18800 13394 18828 13631
rect 18788 13388 18840 13394
rect 18788 13330 18840 13336
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18788 13184 18840 13190
rect 18788 13126 18840 13132
rect 18616 12940 18736 12968
rect 18602 12880 18658 12889
rect 18602 12815 18658 12824
rect 18616 12646 18644 12815
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18604 12436 18656 12442
rect 18604 12378 18656 12384
rect 18616 12170 18644 12378
rect 18604 12164 18656 12170
rect 18604 12106 18656 12112
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 18512 11008 18564 11014
rect 18512 10950 18564 10956
rect 18616 10849 18644 11630
rect 18708 11626 18736 12940
rect 18696 11620 18748 11626
rect 18696 11562 18748 11568
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18602 10840 18658 10849
rect 18602 10775 18658 10784
rect 18420 10736 18472 10742
rect 18420 10678 18472 10684
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18196 8860 18276 8888
rect 18144 8842 18196 8848
rect 18156 8634 18184 8842
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 18236 8288 18288 8294
rect 18236 8230 18288 8236
rect 18248 7993 18276 8230
rect 18340 8022 18368 10542
rect 18432 10305 18460 10678
rect 18510 10432 18566 10441
rect 18510 10367 18566 10376
rect 18418 10296 18474 10305
rect 18418 10231 18474 10240
rect 18420 9988 18472 9994
rect 18420 9930 18472 9936
rect 18432 9897 18460 9930
rect 18418 9888 18474 9897
rect 18418 9823 18474 9832
rect 18524 8906 18552 10367
rect 18604 9444 18656 9450
rect 18604 9386 18656 9392
rect 18512 8900 18564 8906
rect 18512 8842 18564 8848
rect 18328 8016 18380 8022
rect 18234 7984 18290 7993
rect 18328 7958 18380 7964
rect 18234 7919 18290 7928
rect 18248 7818 18276 7919
rect 18236 7812 18288 7818
rect 18236 7754 18288 7760
rect 18144 7472 18196 7478
rect 18144 7414 18196 7420
rect 18050 6896 18106 6905
rect 18050 6831 18106 6840
rect 18064 6633 18092 6831
rect 18050 6624 18106 6633
rect 18050 6559 18106 6568
rect 18050 6488 18106 6497
rect 18050 6423 18052 6432
rect 18104 6423 18106 6432
rect 18052 6394 18104 6400
rect 18156 6254 18184 7414
rect 18524 7206 18552 8842
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18236 6928 18288 6934
rect 18236 6870 18288 6876
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18050 5808 18106 5817
rect 18050 5743 18106 5752
rect 17960 5296 18012 5302
rect 17960 5238 18012 5244
rect 17868 5160 17920 5166
rect 18064 5137 18092 5743
rect 18156 5409 18184 6190
rect 18142 5400 18198 5409
rect 18142 5335 18198 5344
rect 18248 5234 18276 6870
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 18236 5228 18288 5234
rect 18236 5170 18288 5176
rect 17868 5102 17920 5108
rect 18050 5128 18106 5137
rect 18050 5063 18106 5072
rect 18144 5092 18196 5098
rect 18144 5034 18196 5040
rect 18052 4480 18104 4486
rect 18052 4422 18104 4428
rect 17776 3732 17828 3738
rect 17776 3674 17828 3680
rect 18064 3516 18092 4422
rect 18156 4078 18184 5034
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18328 5024 18380 5030
rect 18328 4966 18380 4972
rect 18248 4690 18276 4966
rect 18236 4684 18288 4690
rect 18236 4626 18288 4632
rect 18340 4554 18368 4966
rect 18524 4690 18552 6802
rect 18616 6118 18644 9386
rect 18708 8498 18736 11018
rect 18800 10441 18828 13126
rect 18880 11008 18932 11014
rect 18880 10950 18932 10956
rect 18786 10432 18842 10441
rect 18786 10367 18842 10376
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18696 8288 18748 8294
rect 18696 8230 18748 8236
rect 18708 7478 18736 8230
rect 18892 7478 18920 10950
rect 18984 10198 19012 13631
rect 19076 11150 19104 15506
rect 19168 15162 19288 15178
rect 19352 15162 19380 16526
rect 19156 15156 19288 15162
rect 19208 15150 19288 15156
rect 19156 15098 19208 15104
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19168 13569 19196 13874
rect 19154 13560 19210 13569
rect 19154 13495 19210 13504
rect 19156 13252 19208 13258
rect 19156 13194 19208 13200
rect 19168 11676 19196 13194
rect 19260 13025 19288 15150
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19246 13016 19302 13025
rect 19246 12951 19302 12960
rect 19248 11688 19300 11694
rect 19168 11648 19248 11676
rect 19248 11630 19300 11636
rect 19246 11520 19302 11529
rect 19246 11455 19302 11464
rect 19064 11144 19116 11150
rect 19064 11086 19116 11092
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 18972 10192 19024 10198
rect 18972 10134 19024 10140
rect 19076 9586 19104 10406
rect 19168 10198 19196 10542
rect 19156 10192 19208 10198
rect 19156 10134 19208 10140
rect 19260 9994 19288 11455
rect 19352 11336 19380 14962
rect 19444 12442 19472 17206
rect 19708 17196 19760 17202
rect 19708 17138 19760 17144
rect 19720 17105 19748 17138
rect 19706 17096 19762 17105
rect 19524 17060 19576 17066
rect 19706 17031 19762 17040
rect 19524 17002 19576 17008
rect 19536 16454 19564 17002
rect 19708 16992 19760 16998
rect 19708 16934 19760 16940
rect 19720 16522 19748 16934
rect 20088 16776 20116 18226
rect 20168 17604 20220 17610
rect 20168 17546 20220 17552
rect 20180 17066 20208 17546
rect 20168 17060 20220 17066
rect 20168 17002 20220 17008
rect 19996 16748 20208 16776
rect 19708 16516 19760 16522
rect 19708 16458 19760 16464
rect 19524 16448 19576 16454
rect 19524 16390 19576 16396
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19996 16232 20024 16748
rect 20180 16658 20208 16748
rect 20076 16652 20128 16658
rect 20076 16594 20128 16600
rect 20168 16652 20220 16658
rect 20168 16594 20220 16600
rect 20088 16250 20116 16594
rect 20272 16561 20300 18702
rect 20258 16552 20314 16561
rect 20258 16487 20314 16496
rect 19904 16204 20024 16232
rect 20076 16244 20128 16250
rect 19904 15502 19932 16204
rect 20076 16186 20128 16192
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19616 14816 19668 14822
rect 19616 14758 19668 14764
rect 19628 14414 19656 14758
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19522 13832 19578 13841
rect 19522 13767 19578 13776
rect 19536 13258 19564 13767
rect 19890 13560 19946 13569
rect 19890 13495 19946 13504
rect 19904 13394 19932 13495
rect 19892 13388 19944 13394
rect 19892 13330 19944 13336
rect 19524 13252 19576 13258
rect 19524 13194 19576 13200
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19430 12336 19486 12345
rect 19536 12306 19564 12718
rect 19892 12708 19944 12714
rect 19892 12650 19944 12656
rect 19430 12271 19486 12280
rect 19524 12300 19576 12306
rect 19444 12238 19472 12271
rect 19524 12242 19576 12248
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19904 12170 19932 12650
rect 19996 12209 20024 16050
rect 20088 15638 20116 16186
rect 20168 15904 20220 15910
rect 20168 15846 20220 15852
rect 20076 15632 20128 15638
rect 20076 15574 20128 15580
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 20088 12714 20116 12922
rect 20076 12708 20128 12714
rect 20076 12650 20128 12656
rect 20074 12608 20130 12617
rect 20074 12543 20130 12552
rect 19982 12200 20038 12209
rect 19892 12164 19944 12170
rect 19982 12135 20038 12144
rect 19892 12106 19944 12112
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19352 11308 19472 11336
rect 19444 11257 19472 11308
rect 19430 11248 19486 11257
rect 19340 11212 19392 11218
rect 19430 11183 19486 11192
rect 19616 11212 19668 11218
rect 19340 11154 19392 11160
rect 19616 11154 19668 11160
rect 19248 9988 19300 9994
rect 19248 9930 19300 9936
rect 19064 9580 19116 9586
rect 19064 9522 19116 9528
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 19062 9072 19118 9081
rect 19062 9007 19118 9016
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 18696 7472 18748 7478
rect 18880 7472 18932 7478
rect 18748 7432 18828 7460
rect 18696 7414 18748 7420
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 18694 5808 18750 5817
rect 18694 5743 18750 5752
rect 18604 5160 18656 5166
rect 18604 5102 18656 5108
rect 18512 4684 18564 4690
rect 18512 4626 18564 4632
rect 18328 4548 18380 4554
rect 18328 4490 18380 4496
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 18248 3670 18276 4082
rect 18328 3732 18380 3738
rect 18328 3674 18380 3680
rect 18236 3664 18288 3670
rect 18236 3606 18288 3612
rect 18340 3516 18368 3674
rect 17774 3496 17830 3505
rect 18064 3488 18368 3516
rect 18524 3466 18552 4626
rect 17774 3431 17776 3440
rect 17828 3431 17830 3440
rect 18512 3460 18564 3466
rect 17776 3402 17828 3408
rect 18512 3402 18564 3408
rect 18050 3360 18106 3369
rect 18050 3295 18106 3304
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 17958 3088 18014 3097
rect 18064 3074 18092 3295
rect 18142 3088 18198 3097
rect 18064 3058 18142 3074
rect 17958 3023 18014 3032
rect 18052 3052 18142 3058
rect 17592 2916 17644 2922
rect 17592 2858 17644 2864
rect 17972 2854 18000 3023
rect 18104 3046 18142 3052
rect 18142 3023 18198 3032
rect 18052 2994 18104 3000
rect 18616 2990 18644 5102
rect 18708 4321 18736 5743
rect 18800 4570 18828 7432
rect 18880 7414 18932 7420
rect 18878 7168 18934 7177
rect 18878 7103 18934 7112
rect 18892 4690 18920 7103
rect 18880 4684 18932 4690
rect 18880 4626 18932 4632
rect 18800 4542 18920 4570
rect 18694 4312 18750 4321
rect 18694 4247 18750 4256
rect 18708 3534 18736 4247
rect 18696 3528 18748 3534
rect 18892 3505 18920 4542
rect 18696 3470 18748 3476
rect 18878 3496 18934 3505
rect 18878 3431 18934 3440
rect 18892 2990 18920 3431
rect 18984 3097 19012 8434
rect 19076 7818 19104 9007
rect 19168 8906 19196 9522
rect 19352 9382 19380 11154
rect 19628 11082 19656 11154
rect 19616 11076 19668 11082
rect 19616 11018 19668 11024
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 20088 10130 20116 12543
rect 20180 11150 20208 15846
rect 20272 15609 20300 16487
rect 20258 15600 20314 15609
rect 20258 15535 20314 15544
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20272 13705 20300 15438
rect 20258 13696 20314 13705
rect 20258 13631 20314 13640
rect 20260 13456 20312 13462
rect 20260 13398 20312 13404
rect 20272 11393 20300 13398
rect 20258 11384 20314 11393
rect 20258 11319 20314 11328
rect 20168 11144 20220 11150
rect 20168 11086 20220 11092
rect 20260 11076 20312 11082
rect 20260 11018 20312 11024
rect 20272 10713 20300 11018
rect 20258 10704 20314 10713
rect 20258 10639 20314 10648
rect 20168 10532 20220 10538
rect 20168 10474 20220 10480
rect 20180 10441 20208 10474
rect 20166 10432 20222 10441
rect 20166 10367 20222 10376
rect 20364 10146 20392 19246
rect 20456 16658 20484 19314
rect 20640 19310 20668 19926
rect 20824 19922 20852 25094
rect 21468 24206 21496 37198
rect 21824 37188 21876 37194
rect 21824 37130 21876 37136
rect 21836 34202 21864 37130
rect 21928 36802 21956 39200
rect 22836 36916 22888 36922
rect 22836 36858 22888 36864
rect 21928 36786 22140 36802
rect 21928 36780 22152 36786
rect 21928 36774 22100 36780
rect 22100 36722 22152 36728
rect 22100 36644 22152 36650
rect 22100 36586 22152 36592
rect 21824 34196 21876 34202
rect 21824 34138 21876 34144
rect 22112 27470 22140 36586
rect 22100 27464 22152 27470
rect 22100 27406 22152 27412
rect 22560 27328 22612 27334
rect 22560 27270 22612 27276
rect 22100 26988 22152 26994
rect 22100 26930 22152 26936
rect 21456 24200 21508 24206
rect 21456 24142 21508 24148
rect 21468 22710 21496 24142
rect 22112 23866 22140 26930
rect 22468 26920 22520 26926
rect 22468 26862 22520 26868
rect 22100 23860 22152 23866
rect 22100 23802 22152 23808
rect 21456 22704 21508 22710
rect 21456 22646 21508 22652
rect 21364 22500 21416 22506
rect 21364 22442 21416 22448
rect 20904 20936 20956 20942
rect 20904 20878 20956 20884
rect 20916 20602 20944 20878
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20824 17746 20852 19858
rect 21088 19780 21140 19786
rect 21088 19722 21140 19728
rect 20996 17876 21048 17882
rect 20996 17818 21048 17824
rect 20812 17740 20864 17746
rect 20812 17682 20864 17688
rect 20628 17604 20680 17610
rect 20628 17546 20680 17552
rect 20536 17264 20588 17270
rect 20536 17206 20588 17212
rect 20444 16652 20496 16658
rect 20444 16594 20496 16600
rect 20444 16516 20496 16522
rect 20444 16458 20496 16464
rect 20456 15706 20484 16458
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20442 15600 20498 15609
rect 20442 15535 20498 15544
rect 20456 15026 20484 15535
rect 20444 15020 20496 15026
rect 20444 14962 20496 14968
rect 20444 14272 20496 14278
rect 20444 14214 20496 14220
rect 20456 14006 20484 14214
rect 20444 14000 20496 14006
rect 20444 13942 20496 13948
rect 20444 13252 20496 13258
rect 20444 13194 20496 13200
rect 20456 12782 20484 13194
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20456 12617 20484 12718
rect 20442 12608 20498 12617
rect 20442 12543 20498 12552
rect 20444 12436 20496 12442
rect 20444 12378 20496 12384
rect 20456 11898 20484 12378
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20444 11144 20496 11150
rect 20444 11086 20496 11092
rect 20076 10124 20128 10130
rect 20076 10066 20128 10072
rect 20272 10118 20392 10146
rect 19444 9994 19564 10010
rect 19444 9988 19576 9994
rect 19444 9982 19524 9988
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19156 8900 19208 8906
rect 19156 8842 19208 8848
rect 19444 8616 19472 9982
rect 19524 9930 19576 9936
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19444 8588 19564 8616
rect 19340 8560 19392 8566
rect 19392 8520 19472 8548
rect 19340 8502 19392 8508
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19246 8120 19302 8129
rect 19246 8055 19302 8064
rect 19260 8022 19288 8055
rect 19248 8016 19300 8022
rect 19248 7958 19300 7964
rect 19064 7812 19116 7818
rect 19064 7754 19116 7760
rect 19076 6934 19104 7754
rect 19154 7712 19210 7721
rect 19154 7647 19210 7656
rect 19168 7206 19196 7647
rect 19246 7576 19302 7585
rect 19246 7511 19302 7520
rect 19156 7200 19208 7206
rect 19156 7142 19208 7148
rect 19064 6928 19116 6934
rect 19064 6870 19116 6876
rect 19260 5846 19288 7511
rect 19352 6866 19380 8366
rect 19444 7886 19472 8520
rect 19536 7954 19564 8588
rect 19892 8084 19944 8090
rect 19892 8026 19944 8032
rect 19524 7948 19576 7954
rect 19524 7890 19576 7896
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 19444 7274 19472 7822
rect 19904 7818 19932 8026
rect 19892 7812 19944 7818
rect 19892 7754 19944 7760
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19996 7460 20024 9522
rect 20076 9376 20128 9382
rect 20168 9376 20220 9382
rect 20076 9318 20128 9324
rect 20166 9344 20168 9353
rect 20220 9344 20222 9353
rect 19904 7432 20024 7460
rect 19432 7268 19484 7274
rect 19432 7210 19484 7216
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 19904 6746 19932 7432
rect 19352 6718 19932 6746
rect 19248 5840 19300 5846
rect 19248 5782 19300 5788
rect 19156 5636 19208 5642
rect 19156 5578 19208 5584
rect 19064 5568 19116 5574
rect 19064 5510 19116 5516
rect 19076 3738 19104 5510
rect 19168 5234 19196 5578
rect 19352 5545 19380 6718
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 19444 6372 19472 6598
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19800 6452 19852 6458
rect 20088 6440 20116 9318
rect 20166 9279 20222 9288
rect 20272 7936 20300 10118
rect 20352 9988 20404 9994
rect 20352 9930 20404 9936
rect 20180 7908 20300 7936
rect 20180 7410 20208 7908
rect 20260 7812 20312 7818
rect 20260 7754 20312 7760
rect 20168 7404 20220 7410
rect 20168 7346 20220 7352
rect 19800 6394 19852 6400
rect 19904 6412 20116 6440
rect 19444 6344 19656 6372
rect 19524 6112 19576 6118
rect 19524 6054 19576 6060
rect 19536 5914 19564 6054
rect 19628 5914 19656 6344
rect 19812 6118 19840 6394
rect 19800 6112 19852 6118
rect 19800 6054 19852 6060
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19616 5908 19668 5914
rect 19616 5850 19668 5856
rect 19536 5658 19564 5850
rect 19904 5794 19932 6412
rect 20168 6316 20220 6322
rect 20168 6258 20220 6264
rect 19628 5766 19932 5794
rect 19628 5710 19656 5766
rect 19444 5630 19564 5658
rect 19616 5704 19668 5710
rect 19616 5646 19668 5652
rect 19708 5636 19760 5642
rect 19338 5536 19394 5545
rect 19338 5471 19394 5480
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 19156 5228 19208 5234
rect 19156 5170 19208 5176
rect 19246 4448 19302 4457
rect 19246 4383 19302 4392
rect 19156 4276 19208 4282
rect 19156 4218 19208 4224
rect 19064 3732 19116 3738
rect 19064 3674 19116 3680
rect 18970 3088 19026 3097
rect 18970 3023 19026 3032
rect 18604 2984 18656 2990
rect 18604 2926 18656 2932
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 18880 2984 18932 2990
rect 18880 2926 18932 2932
rect 17960 2848 18012 2854
rect 17960 2790 18012 2796
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 17408 2644 17460 2650
rect 17408 2586 17460 2592
rect 18236 2440 18288 2446
rect 18236 2382 18288 2388
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 16948 1692 17000 1698
rect 16948 1634 17000 1640
rect 17420 800 17448 2246
rect 18248 2106 18276 2382
rect 18236 2100 18288 2106
rect 18236 2042 18288 2048
rect 18052 1760 18104 1766
rect 18052 1702 18104 1708
rect 18064 800 18092 1702
rect 18800 1494 18828 2926
rect 19168 1970 19196 4218
rect 19260 4162 19288 4383
rect 19352 4321 19380 5238
rect 19444 5166 19472 5630
rect 19760 5596 20116 5624
rect 19708 5578 19760 5584
rect 20088 5545 20116 5596
rect 20074 5536 20130 5545
rect 19574 5468 19882 5477
rect 20074 5471 20130 5480
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19982 5400 20038 5409
rect 20180 5370 20208 6258
rect 20272 5914 20300 7754
rect 20364 6458 20392 9930
rect 20456 8956 20484 11086
rect 20548 9654 20576 17206
rect 20640 15570 20668 17546
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20732 15450 20760 16594
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 20640 15422 20760 15450
rect 20640 14074 20668 15422
rect 20720 14272 20772 14278
rect 20720 14214 20772 14220
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20628 13728 20680 13734
rect 20628 13670 20680 13676
rect 20640 13530 20668 13670
rect 20628 13524 20680 13530
rect 20628 13466 20680 13472
rect 20628 12164 20680 12170
rect 20628 12106 20680 12112
rect 20640 11626 20668 12106
rect 20628 11620 20680 11626
rect 20628 11562 20680 11568
rect 20626 11248 20682 11257
rect 20732 11218 20760 14214
rect 20626 11183 20682 11192
rect 20720 11212 20772 11218
rect 20640 11150 20668 11183
rect 20720 11154 20772 11160
rect 20628 11144 20680 11150
rect 20628 11086 20680 11092
rect 20628 11008 20680 11014
rect 20628 10950 20680 10956
rect 20640 10130 20668 10950
rect 20628 10124 20680 10130
rect 20628 10066 20680 10072
rect 20824 9761 20852 16050
rect 20904 14000 20956 14006
rect 20904 13942 20956 13948
rect 20916 12986 20944 13942
rect 21008 13818 21036 17818
rect 21100 16250 21128 19722
rect 21180 17876 21232 17882
rect 21180 17818 21232 17824
rect 21192 17649 21220 17818
rect 21178 17640 21234 17649
rect 21178 17575 21234 17584
rect 21088 16244 21140 16250
rect 21088 16186 21140 16192
rect 21180 15496 21232 15502
rect 21180 15438 21232 15444
rect 21192 14260 21220 15438
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 21284 14414 21312 14962
rect 21376 14550 21404 22442
rect 21548 21616 21600 21622
rect 21548 21558 21600 21564
rect 21456 21140 21508 21146
rect 21456 21082 21508 21088
rect 21468 20806 21496 21082
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 21560 18970 21588 21558
rect 21548 18964 21600 18970
rect 21548 18906 21600 18912
rect 21548 18828 21600 18834
rect 21548 18770 21600 18776
rect 21456 18148 21508 18154
rect 21456 18090 21508 18096
rect 21364 14544 21416 14550
rect 21364 14486 21416 14492
rect 21272 14408 21324 14414
rect 21272 14350 21324 14356
rect 21192 14232 21312 14260
rect 21284 13870 21312 14232
rect 21468 14006 21496 18090
rect 21456 14000 21508 14006
rect 21456 13942 21508 13948
rect 21272 13864 21324 13870
rect 21008 13790 21128 13818
rect 21272 13806 21324 13812
rect 20996 13728 21048 13734
rect 20996 13670 21048 13676
rect 21008 13258 21036 13670
rect 20996 13252 21048 13258
rect 20996 13194 21048 13200
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 20996 11212 21048 11218
rect 20996 11154 21048 11160
rect 20904 11008 20956 11014
rect 20904 10950 20956 10956
rect 20916 10742 20944 10950
rect 20904 10736 20956 10742
rect 20904 10678 20956 10684
rect 21008 10538 21036 11154
rect 21100 10538 21128 13790
rect 21272 13184 21324 13190
rect 21272 13126 21324 13132
rect 21284 12434 21312 13126
rect 21284 12406 21404 12434
rect 21272 12096 21324 12102
rect 21272 12038 21324 12044
rect 21284 11830 21312 12038
rect 21272 11824 21324 11830
rect 21272 11766 21324 11772
rect 21180 11688 21232 11694
rect 21180 11630 21232 11636
rect 21192 11354 21220 11630
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21284 11200 21312 11494
rect 21192 11172 21312 11200
rect 21192 10742 21220 11172
rect 21376 11098 21404 12406
rect 21284 11070 21404 11098
rect 21180 10736 21232 10742
rect 21180 10678 21232 10684
rect 20996 10532 21048 10538
rect 20996 10474 21048 10480
rect 21088 10532 21140 10538
rect 21088 10474 21140 10480
rect 21088 9988 21140 9994
rect 21088 9930 21140 9936
rect 20810 9752 20866 9761
rect 20810 9687 20866 9696
rect 21100 9704 21128 9930
rect 21100 9676 21220 9704
rect 20536 9648 20588 9654
rect 20536 9590 20588 9596
rect 20640 9586 21128 9602
rect 20628 9580 21128 9586
rect 20680 9574 21128 9580
rect 20628 9522 20680 9528
rect 21100 9518 21128 9574
rect 20996 9512 21048 9518
rect 20996 9454 21048 9460
rect 21088 9512 21140 9518
rect 21088 9454 21140 9460
rect 20536 8968 20588 8974
rect 20456 8928 20536 8956
rect 20536 8910 20588 8916
rect 20444 8628 20496 8634
rect 20444 8570 20496 8576
rect 20456 6798 20484 8570
rect 20444 6792 20496 6798
rect 20444 6734 20496 6740
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 20548 5794 20576 8910
rect 21008 8906 21036 9454
rect 20996 8900 21048 8906
rect 20996 8842 21048 8848
rect 20904 8832 20956 8838
rect 20904 8774 20956 8780
rect 20812 8424 20864 8430
rect 20812 8366 20864 8372
rect 20628 8356 20680 8362
rect 20628 8298 20680 8304
rect 20720 8356 20772 8362
rect 20720 8298 20772 8304
rect 20640 7426 20668 8298
rect 20732 7546 20760 8298
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 20640 7398 20760 7426
rect 20824 7410 20852 8366
rect 20732 6474 20760 7398
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 20916 7290 20944 8774
rect 21008 8634 21036 8842
rect 20996 8628 21048 8634
rect 20996 8570 21048 8576
rect 21192 8294 21220 9676
rect 21088 8288 21140 8294
rect 21088 8230 21140 8236
rect 21180 8288 21232 8294
rect 21180 8230 21232 8236
rect 21100 8106 21128 8230
rect 21100 8078 21220 8106
rect 21192 7936 21220 8078
rect 21284 7936 21312 11070
rect 21364 11008 21416 11014
rect 21364 10950 21416 10956
rect 21376 10810 21404 10950
rect 21364 10804 21416 10810
rect 21364 10746 21416 10752
rect 21364 10532 21416 10538
rect 21364 10474 21416 10480
rect 21192 7908 21312 7936
rect 21192 7818 21220 7908
rect 21180 7812 21232 7818
rect 21180 7754 21232 7760
rect 21272 7812 21324 7818
rect 21272 7754 21324 7760
rect 21284 7546 21312 7754
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 20640 6446 20760 6474
rect 20824 7262 20944 7290
rect 20640 6322 20668 6446
rect 20718 6352 20774 6361
rect 20628 6316 20680 6322
rect 20718 6287 20774 6296
rect 20628 6258 20680 6264
rect 20628 6180 20680 6186
rect 20628 6122 20680 6128
rect 20640 5914 20668 6122
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20260 5772 20312 5778
rect 20548 5766 20668 5794
rect 20260 5714 20312 5720
rect 20272 5409 20300 5714
rect 20534 5536 20590 5545
rect 20534 5471 20590 5480
rect 20258 5400 20314 5409
rect 19982 5335 19984 5344
rect 20036 5335 20038 5344
rect 20168 5364 20220 5370
rect 19984 5306 20036 5312
rect 20258 5335 20314 5344
rect 20168 5306 20220 5312
rect 19524 5296 19576 5302
rect 20260 5296 20312 5302
rect 19524 5238 19576 5244
rect 20088 5244 20260 5250
rect 20088 5238 20312 5244
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 19536 4468 19564 5238
rect 19708 5228 19760 5234
rect 20088 5222 20300 5238
rect 19760 5188 19840 5216
rect 19708 5170 19760 5176
rect 19812 5148 19840 5188
rect 20088 5148 20116 5222
rect 19812 5120 20116 5148
rect 20352 5092 20404 5098
rect 20352 5034 20404 5040
rect 20364 4978 20392 5034
rect 20364 4950 20484 4978
rect 19996 4780 20300 4808
rect 19996 4706 20024 4780
rect 19720 4678 20024 4706
rect 19720 4554 19748 4678
rect 20272 4554 20300 4780
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 19708 4548 19760 4554
rect 19708 4490 19760 4496
rect 20168 4548 20220 4554
rect 20168 4490 20220 4496
rect 20260 4548 20312 4554
rect 20260 4490 20312 4496
rect 19444 4440 19564 4468
rect 19800 4480 19852 4486
rect 19338 4312 19394 4321
rect 19338 4247 19394 4256
rect 19444 4264 19472 4440
rect 19852 4440 20024 4468
rect 19800 4422 19852 4428
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19996 4321 20024 4440
rect 19982 4312 20038 4321
rect 19616 4276 19668 4282
rect 19444 4236 19616 4264
rect 19982 4247 20038 4256
rect 20180 4298 20208 4490
rect 20364 4486 20392 4558
rect 20352 4480 20404 4486
rect 20352 4422 20404 4428
rect 20456 4298 20484 4950
rect 20548 4865 20576 5471
rect 20640 5409 20668 5766
rect 20626 5400 20682 5409
rect 20626 5335 20682 5344
rect 20534 4856 20590 4865
rect 20732 4842 20760 6287
rect 20824 5710 20852 7262
rect 20904 7200 20956 7206
rect 20904 7142 20956 7148
rect 20916 6934 20944 7142
rect 21178 7032 21234 7041
rect 21178 6967 21234 6976
rect 20904 6928 20956 6934
rect 20904 6870 20956 6876
rect 20904 6724 20956 6730
rect 20904 6666 20956 6672
rect 20916 6458 20944 6666
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 21088 6384 21140 6390
rect 21008 6344 21088 6372
rect 20904 6316 20956 6322
rect 20904 6258 20956 6264
rect 20916 6118 20944 6258
rect 20904 6112 20956 6118
rect 20904 6054 20956 6060
rect 20812 5704 20864 5710
rect 20812 5646 20864 5652
rect 20902 5672 20958 5681
rect 20902 5607 20958 5616
rect 20534 4791 20590 4800
rect 20640 4814 20760 4842
rect 20548 4622 20576 4791
rect 20536 4616 20588 4622
rect 20536 4558 20588 4564
rect 20180 4270 20484 4298
rect 20640 4298 20668 4814
rect 20718 4720 20774 4729
rect 20718 4655 20774 4664
rect 20732 4486 20760 4655
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20720 4480 20772 4486
rect 20720 4422 20772 4428
rect 20640 4270 20760 4298
rect 19616 4218 19668 4224
rect 19260 4134 19334 4162
rect 19306 4128 19334 4134
rect 19984 4140 20036 4146
rect 19306 4100 19380 4128
rect 19352 3777 19380 4100
rect 19984 4082 20036 4088
rect 19338 3768 19394 3777
rect 19338 3703 19394 3712
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19536 3534 19564 3674
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19246 3224 19302 3233
rect 19574 3227 19882 3236
rect 19246 3159 19302 3168
rect 19260 2990 19288 3159
rect 19996 3126 20024 4082
rect 19984 3120 20036 3126
rect 19984 3062 20036 3068
rect 20076 3120 20128 3126
rect 20076 3062 20128 3068
rect 19248 2984 19300 2990
rect 20088 2961 20116 3062
rect 19248 2926 19300 2932
rect 20074 2952 20130 2961
rect 20074 2887 20130 2896
rect 20180 2650 20208 4270
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 20272 2922 20300 4082
rect 20732 3534 20760 4270
rect 20824 4214 20852 4558
rect 20812 4208 20864 4214
rect 20812 4150 20864 4156
rect 20812 4072 20864 4078
rect 20812 4014 20864 4020
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20628 3460 20680 3466
rect 20628 3402 20680 3408
rect 20640 3346 20668 3402
rect 20640 3318 20760 3346
rect 20732 3126 20760 3318
rect 20824 3194 20852 4014
rect 20916 3398 20944 5607
rect 21008 3942 21036 6344
rect 21088 6326 21140 6332
rect 21088 6248 21140 6254
rect 21088 6190 21140 6196
rect 21100 6118 21128 6190
rect 21088 6112 21140 6118
rect 21088 6054 21140 6060
rect 21192 5574 21220 6967
rect 21284 6662 21312 7482
rect 21376 7410 21404 10474
rect 21468 10198 21496 13942
rect 21560 10198 21588 18770
rect 22112 18222 22140 23802
rect 22376 22976 22428 22982
rect 22376 22918 22428 22924
rect 22388 22574 22416 22918
rect 22192 22568 22244 22574
rect 22192 22510 22244 22516
rect 22376 22568 22428 22574
rect 22376 22510 22428 22516
rect 22204 22438 22232 22510
rect 22192 22432 22244 22438
rect 22192 22374 22244 22380
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 22204 20466 22232 21830
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22388 20602 22416 20878
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 22376 20392 22428 20398
rect 22376 20334 22428 20340
rect 22284 18352 22336 18358
rect 22284 18294 22336 18300
rect 22100 18216 22152 18222
rect 22100 18158 22152 18164
rect 22008 17672 22060 17678
rect 22008 17614 22060 17620
rect 22020 16658 22048 17614
rect 22008 16652 22060 16658
rect 22008 16594 22060 16600
rect 21640 16176 21692 16182
rect 21640 16118 21692 16124
rect 21652 15706 21680 16118
rect 22296 15978 22324 18294
rect 22388 17814 22416 20334
rect 22480 19922 22508 26862
rect 22572 20262 22600 27270
rect 22652 22976 22704 22982
rect 22652 22918 22704 22924
rect 22560 20256 22612 20262
rect 22560 20198 22612 20204
rect 22468 19916 22520 19922
rect 22468 19858 22520 19864
rect 22572 19718 22600 20198
rect 22664 19922 22692 22918
rect 22652 19916 22704 19922
rect 22652 19858 22704 19864
rect 22560 19712 22612 19718
rect 22560 19654 22612 19660
rect 22376 17808 22428 17814
rect 22376 17750 22428 17756
rect 22376 17128 22428 17134
rect 22376 17070 22428 17076
rect 22388 16794 22416 17070
rect 22376 16788 22428 16794
rect 22376 16730 22428 16736
rect 22560 16448 22612 16454
rect 22560 16390 22612 16396
rect 22468 16176 22520 16182
rect 22468 16118 22520 16124
rect 22284 15972 22336 15978
rect 22284 15914 22336 15920
rect 21640 15700 21692 15706
rect 21640 15642 21692 15648
rect 22374 15464 22430 15473
rect 22374 15399 22430 15408
rect 22100 14816 22152 14822
rect 22100 14758 22152 14764
rect 22112 14414 22140 14758
rect 22100 14408 22152 14414
rect 22100 14350 22152 14356
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 21640 14340 21692 14346
rect 21640 14282 21692 14288
rect 21456 10192 21508 10198
rect 21456 10134 21508 10140
rect 21548 10192 21600 10198
rect 21548 10134 21600 10140
rect 21560 9586 21588 10134
rect 21548 9580 21600 9586
rect 21548 9522 21600 9528
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 21454 7440 21510 7449
rect 21364 7404 21416 7410
rect 21454 7375 21510 7384
rect 21364 7346 21416 7352
rect 21362 6896 21418 6905
rect 21362 6831 21418 6840
rect 21272 6656 21324 6662
rect 21272 6598 21324 6604
rect 21376 6474 21404 6831
rect 21468 6662 21496 7375
rect 21560 6866 21588 9114
rect 21652 8974 21680 14282
rect 22296 13530 22324 14350
rect 22284 13524 22336 13530
rect 22284 13466 22336 13472
rect 22098 13424 22154 13433
rect 22098 13359 22154 13368
rect 22112 13326 22140 13359
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 22100 12912 22152 12918
rect 22100 12854 22152 12860
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 21824 12096 21876 12102
rect 21824 12038 21876 12044
rect 21732 11552 21784 11558
rect 21730 11520 21732 11529
rect 21784 11520 21786 11529
rect 21730 11455 21786 11464
rect 21836 11218 21864 12038
rect 22020 11665 22048 12174
rect 22006 11656 22062 11665
rect 22006 11591 22062 11600
rect 21914 11384 21970 11393
rect 21914 11319 21970 11328
rect 21824 11212 21876 11218
rect 21824 11154 21876 11160
rect 21928 11150 21956 11319
rect 21916 11144 21968 11150
rect 21916 11086 21968 11092
rect 22006 11112 22062 11121
rect 22006 11047 22062 11056
rect 21732 10600 21784 10606
rect 21732 10542 21784 10548
rect 21744 9994 21772 10542
rect 21732 9988 21784 9994
rect 21732 9930 21784 9936
rect 21916 9988 21968 9994
rect 21916 9930 21968 9936
rect 21928 9722 21956 9930
rect 22020 9926 22048 11047
rect 22008 9920 22060 9926
rect 22008 9862 22060 9868
rect 21916 9716 21968 9722
rect 21916 9658 21968 9664
rect 22112 9586 22140 12854
rect 22296 11694 22324 13466
rect 22388 11694 22416 15399
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22376 11688 22428 11694
rect 22376 11630 22428 11636
rect 22192 10668 22244 10674
rect 22192 10610 22244 10616
rect 22008 9580 22060 9586
rect 22008 9522 22060 9528
rect 22100 9580 22152 9586
rect 22100 9522 22152 9528
rect 22020 9450 22048 9522
rect 22204 9466 22232 10610
rect 22284 10056 22336 10062
rect 22284 9998 22336 10004
rect 22296 9722 22324 9998
rect 22284 9716 22336 9722
rect 22284 9658 22336 9664
rect 22284 9580 22336 9586
rect 22284 9522 22336 9528
rect 21732 9444 21784 9450
rect 21732 9386 21784 9392
rect 22008 9444 22060 9450
rect 22008 9386 22060 9392
rect 22112 9438 22232 9466
rect 21744 9178 21772 9386
rect 21732 9172 21784 9178
rect 21732 9114 21784 9120
rect 22112 8974 22140 9438
rect 22192 9376 22244 9382
rect 22192 9318 22244 9324
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 22100 8968 22152 8974
rect 22100 8910 22152 8916
rect 21548 6860 21600 6866
rect 21548 6802 21600 6808
rect 21456 6656 21508 6662
rect 21456 6598 21508 6604
rect 21376 6446 21496 6474
rect 21272 5704 21324 5710
rect 21272 5646 21324 5652
rect 21364 5704 21416 5710
rect 21364 5646 21416 5652
rect 21180 5568 21232 5574
rect 21180 5510 21232 5516
rect 21178 5400 21234 5409
rect 21178 5335 21234 5344
rect 21086 5264 21142 5273
rect 21086 5199 21088 5208
rect 21140 5199 21142 5208
rect 21088 5170 21140 5176
rect 21192 4622 21220 5335
rect 21180 4616 21232 4622
rect 21180 4558 21232 4564
rect 20996 3936 21048 3942
rect 20996 3878 21048 3884
rect 21088 3936 21140 3942
rect 21088 3878 21140 3884
rect 21100 3602 21128 3878
rect 21192 3777 21220 4558
rect 21178 3768 21234 3777
rect 21178 3703 21234 3712
rect 21088 3596 21140 3602
rect 21088 3538 21140 3544
rect 20904 3392 20956 3398
rect 20904 3334 20956 3340
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 20628 3120 20680 3126
rect 20628 3062 20680 3068
rect 20720 3120 20772 3126
rect 20720 3062 20772 3068
rect 20260 2916 20312 2922
rect 20260 2858 20312 2864
rect 20640 2774 20668 3062
rect 21284 2854 21312 5646
rect 21272 2848 21324 2854
rect 21272 2790 21324 2796
rect 20456 2746 20668 2774
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 19340 2372 19392 2378
rect 19340 2314 19392 2320
rect 19156 1964 19208 1970
rect 19156 1906 19208 1912
rect 18788 1488 18840 1494
rect 18788 1430 18840 1436
rect 19352 800 19380 2314
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 20088 1834 20116 2382
rect 20076 1828 20128 1834
rect 20076 1770 20128 1776
rect 20456 1562 20484 2746
rect 21376 2650 21404 5646
rect 21468 3534 21496 6446
rect 21652 5302 21680 8910
rect 22112 8514 22140 8910
rect 21744 8486 22140 8514
rect 21744 8265 21772 8486
rect 22008 8424 22060 8430
rect 22008 8366 22060 8372
rect 21916 8288 21968 8294
rect 21730 8256 21786 8265
rect 21916 8230 21968 8236
rect 21730 8191 21786 8200
rect 21732 6928 21784 6934
rect 21732 6870 21784 6876
rect 21548 5296 21600 5302
rect 21548 5238 21600 5244
rect 21640 5296 21692 5302
rect 21640 5238 21692 5244
rect 21560 5098 21588 5238
rect 21548 5092 21600 5098
rect 21548 5034 21600 5040
rect 21744 5030 21772 6870
rect 21822 5808 21878 5817
rect 21822 5743 21878 5752
rect 21836 5710 21864 5743
rect 21824 5704 21876 5710
rect 21824 5646 21876 5652
rect 21928 5098 21956 8230
rect 22020 7954 22048 8366
rect 22112 7954 22140 8486
rect 22008 7948 22060 7954
rect 22008 7890 22060 7896
rect 22100 7948 22152 7954
rect 22100 7890 22152 7896
rect 22204 7410 22232 9318
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 22296 7342 22324 9522
rect 22388 8498 22416 11630
rect 22376 8492 22428 8498
rect 22376 8434 22428 8440
rect 22480 8129 22508 16118
rect 22572 12170 22600 16390
rect 22848 12918 22876 36858
rect 23216 36786 23244 39200
rect 24504 37126 24532 39200
rect 25148 37262 25176 39200
rect 26436 37262 26464 39200
rect 25136 37256 25188 37262
rect 25136 37198 25188 37204
rect 26424 37256 26476 37262
rect 26424 37198 26476 37204
rect 27724 37126 27752 39200
rect 28368 37262 28396 39200
rect 29656 37262 29684 39200
rect 30944 37262 30972 39200
rect 27896 37256 27948 37262
rect 27896 37198 27948 37204
rect 28356 37256 28408 37262
rect 28356 37198 28408 37204
rect 29644 37256 29696 37262
rect 29644 37198 29696 37204
rect 30932 37256 30984 37262
rect 30932 37198 30984 37204
rect 24492 37120 24544 37126
rect 24492 37062 24544 37068
rect 25320 37120 25372 37126
rect 25320 37062 25372 37068
rect 27712 37120 27764 37126
rect 27712 37062 27764 37068
rect 23204 36780 23256 36786
rect 23204 36722 23256 36728
rect 23572 32224 23624 32230
rect 23572 32166 23624 32172
rect 23584 31958 23612 32166
rect 23572 31952 23624 31958
rect 23572 31894 23624 31900
rect 25332 31890 25360 37062
rect 27620 36236 27672 36242
rect 27620 36178 27672 36184
rect 25320 31884 25372 31890
rect 25320 31826 25372 31832
rect 27632 31822 27660 36178
rect 27804 31884 27856 31890
rect 27804 31826 27856 31832
rect 27620 31816 27672 31822
rect 27620 31758 27672 31764
rect 26148 30728 26200 30734
rect 26148 30670 26200 30676
rect 26160 25294 26188 30670
rect 27816 25702 27844 31826
rect 27908 30938 27936 37198
rect 28264 37188 28316 37194
rect 28264 37130 28316 37136
rect 28276 32910 28304 37130
rect 32232 37126 32260 39200
rect 32772 37324 32824 37330
rect 32772 37266 32824 37272
rect 32312 37256 32364 37262
rect 32312 37198 32364 37204
rect 32404 37256 32456 37262
rect 32404 37198 32456 37204
rect 28632 37120 28684 37126
rect 28632 37062 28684 37068
rect 28724 37120 28776 37126
rect 28724 37062 28776 37068
rect 32220 37120 32272 37126
rect 32220 37062 32272 37068
rect 28264 32904 28316 32910
rect 28264 32846 28316 32852
rect 28356 32768 28408 32774
rect 28356 32710 28408 32716
rect 27896 30932 27948 30938
rect 27896 30874 27948 30880
rect 28080 30592 28132 30598
rect 28080 30534 28132 30540
rect 28092 27130 28120 30534
rect 28080 27124 28132 27130
rect 28080 27066 28132 27072
rect 28368 26926 28396 32710
rect 28644 32434 28672 37062
rect 28736 36242 28764 37062
rect 32324 36922 32352 37198
rect 32312 36916 32364 36922
rect 32312 36858 32364 36864
rect 28724 36236 28776 36242
rect 28724 36178 28776 36184
rect 30472 32904 30524 32910
rect 30472 32846 30524 32852
rect 28632 32428 28684 32434
rect 28632 32370 28684 32376
rect 30484 29850 30512 32846
rect 30472 29844 30524 29850
rect 30472 29786 30524 29792
rect 32416 29714 32444 37198
rect 32784 35894 32812 37266
rect 32876 37210 32904 39200
rect 34164 39114 34192 39200
rect 34256 39114 34284 39222
rect 34164 39086 34284 39114
rect 34440 37210 34468 39222
rect 35438 39200 35494 39800
rect 36082 39200 36138 39800
rect 37370 39200 37426 39800
rect 38658 39200 38714 39800
rect 39302 39200 39358 39800
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34796 37256 34848 37262
rect 32876 37182 33180 37210
rect 34440 37182 34560 37210
rect 34796 37198 34848 37204
rect 33152 37126 33180 37182
rect 34532 37126 34560 37182
rect 33140 37120 33192 37126
rect 33140 37062 33192 37068
rect 34520 37120 34572 37126
rect 34520 37062 34572 37068
rect 33140 36644 33192 36650
rect 33140 36586 33192 36592
rect 32784 35866 32904 35894
rect 32404 29708 32456 29714
rect 32404 29650 32456 29656
rect 28356 26920 28408 26926
rect 28356 26862 28408 26868
rect 27804 25696 27856 25702
rect 27804 25638 27856 25644
rect 26148 25288 26200 25294
rect 26148 25230 26200 25236
rect 30104 25288 30156 25294
rect 30104 25230 30156 25236
rect 23296 24336 23348 24342
rect 23296 24278 23348 24284
rect 23308 23730 23336 24278
rect 30116 24274 30144 25230
rect 32680 24812 32732 24818
rect 32680 24754 32732 24760
rect 30104 24268 30156 24274
rect 30104 24210 30156 24216
rect 31116 24064 31168 24070
rect 31116 24006 31168 24012
rect 23296 23724 23348 23730
rect 23296 23666 23348 23672
rect 25412 23724 25464 23730
rect 25412 23666 25464 23672
rect 23940 23520 23992 23526
rect 23940 23462 23992 23468
rect 23848 22636 23900 22642
rect 23848 22578 23900 22584
rect 23296 22568 23348 22574
rect 23296 22510 23348 22516
rect 23204 22432 23256 22438
rect 23204 22374 23256 22380
rect 22928 22160 22980 22166
rect 22928 22102 22980 22108
rect 22940 17678 22968 22102
rect 23020 22024 23072 22030
rect 23020 21966 23072 21972
rect 23032 21554 23060 21966
rect 23216 21690 23244 22374
rect 23308 22030 23336 22510
rect 23756 22432 23808 22438
rect 23756 22374 23808 22380
rect 23296 22024 23348 22030
rect 23296 21966 23348 21972
rect 23296 21888 23348 21894
rect 23296 21830 23348 21836
rect 23204 21684 23256 21690
rect 23204 21626 23256 21632
rect 23112 21616 23164 21622
rect 23112 21558 23164 21564
rect 23020 21548 23072 21554
rect 23020 21490 23072 21496
rect 23124 21350 23152 21558
rect 23112 21344 23164 21350
rect 23112 21286 23164 21292
rect 23216 21078 23244 21626
rect 23204 21072 23256 21078
rect 23204 21014 23256 21020
rect 23112 19508 23164 19514
rect 23112 19450 23164 19456
rect 22928 17672 22980 17678
rect 22928 17614 22980 17620
rect 22940 17270 22968 17614
rect 22928 17264 22980 17270
rect 22928 17206 22980 17212
rect 23124 16182 23152 19450
rect 23204 19236 23256 19242
rect 23204 19178 23256 19184
rect 23216 18358 23244 19178
rect 23204 18352 23256 18358
rect 23204 18294 23256 18300
rect 23112 16176 23164 16182
rect 23112 16118 23164 16124
rect 23308 15065 23336 21830
rect 23768 21486 23796 22374
rect 23756 21480 23808 21486
rect 23756 21422 23808 21428
rect 23480 19168 23532 19174
rect 23480 19110 23532 19116
rect 23492 18698 23520 19110
rect 23480 18692 23532 18698
rect 23480 18634 23532 18640
rect 23860 18306 23888 22578
rect 23952 19718 23980 23462
rect 25424 23118 25452 23666
rect 25412 23112 25464 23118
rect 25412 23054 25464 23060
rect 27988 23044 28040 23050
rect 27988 22986 28040 22992
rect 24768 22432 24820 22438
rect 24768 22374 24820 22380
rect 24492 21344 24544 21350
rect 24492 21286 24544 21292
rect 24504 20806 24532 21286
rect 24492 20800 24544 20806
rect 24492 20742 24544 20748
rect 24676 20800 24728 20806
rect 24676 20742 24728 20748
rect 24400 19780 24452 19786
rect 24400 19722 24452 19728
rect 23940 19712 23992 19718
rect 23940 19654 23992 19660
rect 24124 19372 24176 19378
rect 24124 19314 24176 19320
rect 23940 18896 23992 18902
rect 23940 18838 23992 18844
rect 23952 18630 23980 18838
rect 23940 18624 23992 18630
rect 23940 18566 23992 18572
rect 23676 18278 23888 18306
rect 23388 15360 23440 15366
rect 23388 15302 23440 15308
rect 23294 15056 23350 15065
rect 23294 14991 23350 15000
rect 22836 12912 22888 12918
rect 22836 12854 22888 12860
rect 22652 12708 22704 12714
rect 22652 12650 22704 12656
rect 22560 12164 22612 12170
rect 22560 12106 22612 12112
rect 22664 11098 22692 12650
rect 23020 11892 23072 11898
rect 23020 11834 23072 11840
rect 23032 11665 23060 11834
rect 23294 11792 23350 11801
rect 23294 11727 23350 11736
rect 23018 11656 23074 11665
rect 23018 11591 23074 11600
rect 23204 11552 23256 11558
rect 23204 11494 23256 11500
rect 23112 11348 23164 11354
rect 23112 11290 23164 11296
rect 22572 11070 22692 11098
rect 22836 11144 22888 11150
rect 22836 11086 22888 11092
rect 22466 8120 22522 8129
rect 22466 8055 22522 8064
rect 22284 7336 22336 7342
rect 22284 7278 22336 7284
rect 22468 7336 22520 7342
rect 22468 7278 22520 7284
rect 22296 6934 22324 7278
rect 22284 6928 22336 6934
rect 22284 6870 22336 6876
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 21916 5092 21968 5098
rect 21916 5034 21968 5040
rect 21732 5024 21784 5030
rect 21732 4966 21784 4972
rect 22006 4992 22062 5001
rect 22006 4927 22062 4936
rect 21914 4312 21970 4321
rect 21914 4247 21970 4256
rect 21548 4072 21600 4078
rect 21546 4040 21548 4049
rect 21600 4040 21602 4049
rect 21546 3975 21602 3984
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 21928 3398 21956 4247
rect 22020 4146 22048 4927
rect 22008 4140 22060 4146
rect 22008 4082 22060 4088
rect 22112 3534 22140 6734
rect 22376 6724 22428 6730
rect 22376 6666 22428 6672
rect 22388 5914 22416 6666
rect 22284 5908 22336 5914
rect 22284 5850 22336 5856
rect 22376 5908 22428 5914
rect 22376 5850 22428 5856
rect 22296 5778 22324 5850
rect 22284 5772 22336 5778
rect 22284 5714 22336 5720
rect 22284 5364 22336 5370
rect 22284 5306 22336 5312
rect 22376 5364 22428 5370
rect 22376 5306 22428 5312
rect 22192 5296 22244 5302
rect 22192 5238 22244 5244
rect 22204 3738 22232 5238
rect 22296 4486 22324 5306
rect 22284 4480 22336 4486
rect 22284 4422 22336 4428
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 22192 3732 22244 3738
rect 22192 3674 22244 3680
rect 22100 3528 22152 3534
rect 22152 3476 22232 3482
rect 22100 3470 22232 3476
rect 22112 3454 22232 3470
rect 22296 3466 22324 4082
rect 21548 3392 21600 3398
rect 21548 3334 21600 3340
rect 21916 3392 21968 3398
rect 21916 3334 21968 3340
rect 21364 2644 21416 2650
rect 21364 2586 21416 2592
rect 21560 2514 21588 3334
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 21916 2984 21968 2990
rect 21916 2926 21968 2932
rect 21548 2508 21600 2514
rect 21548 2450 21600 2456
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 20444 1556 20496 1562
rect 20444 1498 20496 1504
rect 20640 800 20668 2382
rect 21928 800 21956 2926
rect 22020 2446 22048 3130
rect 22100 2848 22152 2854
rect 22100 2790 22152 2796
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 22112 1737 22140 2790
rect 22204 2310 22232 3454
rect 22284 3460 22336 3466
rect 22284 3402 22336 3408
rect 22192 2304 22244 2310
rect 22192 2246 22244 2252
rect 22388 2106 22416 5306
rect 22480 3058 22508 7278
rect 22572 5302 22600 11070
rect 22652 11008 22704 11014
rect 22652 10950 22704 10956
rect 22664 10266 22692 10950
rect 22742 10568 22798 10577
rect 22742 10503 22744 10512
rect 22796 10503 22798 10512
rect 22744 10474 22796 10480
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22848 9586 22876 11086
rect 23020 9988 23072 9994
rect 23020 9930 23072 9936
rect 22836 9580 22888 9586
rect 22836 9522 22888 9528
rect 22650 9480 22706 9489
rect 22650 9415 22706 9424
rect 22664 8498 22692 9415
rect 22744 8968 22796 8974
rect 22742 8936 22744 8945
rect 22796 8936 22798 8945
rect 22742 8871 22798 8880
rect 22836 8832 22888 8838
rect 22836 8774 22888 8780
rect 22848 8566 22876 8774
rect 22836 8560 22888 8566
rect 22836 8502 22888 8508
rect 22652 8492 22704 8498
rect 22652 8434 22704 8440
rect 22744 8424 22796 8430
rect 22744 8366 22796 8372
rect 22650 8120 22706 8129
rect 22650 8055 22706 8064
rect 22664 7818 22692 8055
rect 22652 7812 22704 7818
rect 22652 7754 22704 7760
rect 22652 6792 22704 6798
rect 22652 6734 22704 6740
rect 22664 5778 22692 6734
rect 22756 6458 22784 8366
rect 22836 8288 22888 8294
rect 22836 8230 22888 8236
rect 22848 7750 22876 8230
rect 22836 7744 22888 7750
rect 22836 7686 22888 7692
rect 22928 7744 22980 7750
rect 22928 7686 22980 7692
rect 22744 6452 22796 6458
rect 22744 6394 22796 6400
rect 22940 6118 22968 7686
rect 23032 6254 23060 9930
rect 23124 6798 23152 11290
rect 23216 11150 23244 11494
rect 23308 11354 23336 11727
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 23204 11144 23256 11150
rect 23400 11098 23428 15302
rect 23478 13560 23534 13569
rect 23478 13495 23534 13504
rect 23204 11086 23256 11092
rect 23308 11070 23428 11098
rect 23308 10962 23336 11070
rect 23216 10934 23336 10962
rect 23386 10976 23442 10985
rect 23216 10062 23244 10934
rect 23386 10911 23442 10920
rect 23204 10056 23256 10062
rect 23204 9998 23256 10004
rect 23112 6792 23164 6798
rect 23112 6734 23164 6740
rect 23216 6610 23244 9998
rect 23400 9586 23428 10911
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23492 9178 23520 13495
rect 23572 12844 23624 12850
rect 23572 12786 23624 12792
rect 23584 11762 23612 12786
rect 23572 11756 23624 11762
rect 23572 11698 23624 11704
rect 23676 11642 23704 18278
rect 23756 18216 23808 18222
rect 23756 18158 23808 18164
rect 23584 11614 23704 11642
rect 23584 10742 23612 11614
rect 23664 11552 23716 11558
rect 23768 11540 23796 18158
rect 24136 17882 24164 19314
rect 24124 17876 24176 17882
rect 24124 17818 24176 17824
rect 24412 16998 24440 19722
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 24504 12306 24532 20742
rect 24688 19786 24716 20742
rect 24780 19786 24808 22374
rect 28000 21554 28028 22986
rect 27068 21548 27120 21554
rect 27068 21490 27120 21496
rect 27988 21548 28040 21554
rect 27988 21490 28040 21496
rect 26240 20936 26292 20942
rect 26240 20878 26292 20884
rect 24952 19916 25004 19922
rect 24952 19858 25004 19864
rect 24676 19780 24728 19786
rect 24676 19722 24728 19728
rect 24768 19780 24820 19786
rect 24768 19722 24820 19728
rect 24584 19712 24636 19718
rect 24584 19654 24636 19660
rect 24596 16658 24624 19654
rect 24676 19304 24728 19310
rect 24676 19246 24728 19252
rect 24688 18834 24716 19246
rect 24860 19168 24912 19174
rect 24860 19110 24912 19116
rect 24676 18828 24728 18834
rect 24676 18770 24728 18776
rect 24872 18698 24900 19110
rect 24860 18692 24912 18698
rect 24860 18634 24912 18640
rect 24964 18222 24992 19858
rect 26252 19242 26280 20878
rect 26792 20256 26844 20262
rect 26792 20198 26844 20204
rect 26804 19922 26832 20198
rect 26792 19916 26844 19922
rect 26792 19858 26844 19864
rect 26240 19236 26292 19242
rect 26240 19178 26292 19184
rect 26240 18964 26292 18970
rect 26240 18906 26292 18912
rect 26252 18766 26280 18906
rect 26240 18760 26292 18766
rect 26240 18702 26292 18708
rect 25136 18284 25188 18290
rect 25136 18226 25188 18232
rect 24952 18216 25004 18222
rect 24952 18158 25004 18164
rect 24584 16652 24636 16658
rect 24584 16594 24636 16600
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 24674 13968 24730 13977
rect 24674 13903 24730 13912
rect 24492 12300 24544 12306
rect 24492 12242 24544 12248
rect 24124 11756 24176 11762
rect 24124 11698 24176 11704
rect 23716 11512 23796 11540
rect 23664 11494 23716 11500
rect 23572 10736 23624 10742
rect 23572 10678 23624 10684
rect 23584 10169 23612 10678
rect 23676 10470 23704 11494
rect 23756 10804 23808 10810
rect 23756 10746 23808 10752
rect 23664 10464 23716 10470
rect 23664 10406 23716 10412
rect 23768 10282 23796 10746
rect 23676 10254 23796 10282
rect 23570 10160 23626 10169
rect 23570 10095 23626 10104
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23386 8528 23442 8537
rect 23296 8492 23348 8498
rect 23386 8463 23388 8472
rect 23296 8434 23348 8440
rect 23440 8463 23442 8472
rect 23388 8434 23440 8440
rect 23308 8022 23336 8434
rect 23296 8016 23348 8022
rect 23296 7958 23348 7964
rect 23388 7744 23440 7750
rect 23388 7686 23440 7692
rect 23400 7478 23428 7686
rect 23388 7472 23440 7478
rect 23388 7414 23440 7420
rect 23388 6928 23440 6934
rect 23388 6870 23440 6876
rect 23296 6792 23348 6798
rect 23294 6760 23296 6769
rect 23348 6760 23350 6769
rect 23294 6695 23350 6704
rect 23124 6582 23244 6610
rect 23020 6248 23072 6254
rect 23020 6190 23072 6196
rect 23124 6186 23152 6582
rect 23204 6248 23256 6254
rect 23204 6190 23256 6196
rect 23112 6180 23164 6186
rect 23112 6122 23164 6128
rect 22928 6112 22980 6118
rect 22834 6080 22890 6089
rect 22928 6054 22980 6060
rect 22834 6015 22890 6024
rect 22652 5772 22704 5778
rect 22652 5714 22704 5720
rect 22560 5296 22612 5302
rect 22560 5238 22612 5244
rect 22664 5114 22692 5714
rect 22572 5086 22692 5114
rect 22572 3942 22600 5086
rect 22744 4004 22796 4010
rect 22744 3946 22796 3952
rect 22560 3936 22612 3942
rect 22560 3878 22612 3884
rect 22572 3097 22600 3878
rect 22652 3528 22704 3534
rect 22756 3505 22784 3946
rect 22848 3738 22876 6015
rect 23216 5778 23244 6190
rect 23294 5944 23350 5953
rect 23294 5879 23350 5888
rect 23204 5772 23256 5778
rect 23204 5714 23256 5720
rect 23216 5250 23244 5714
rect 23124 5234 23244 5250
rect 23112 5228 23244 5234
rect 23164 5222 23244 5228
rect 23112 5170 23164 5176
rect 23020 5160 23072 5166
rect 23020 5102 23072 5108
rect 22836 3732 22888 3738
rect 22836 3674 22888 3680
rect 22652 3470 22704 3476
rect 22742 3496 22798 3505
rect 22664 3194 22692 3470
rect 22742 3431 22798 3440
rect 22652 3188 22704 3194
rect 22652 3130 22704 3136
rect 22558 3088 22614 3097
rect 22468 3052 22520 3058
rect 22558 3023 22614 3032
rect 22664 3046 22968 3074
rect 22468 2994 22520 3000
rect 22664 2922 22692 3046
rect 22940 2990 22968 3046
rect 22928 2984 22980 2990
rect 22928 2926 22980 2932
rect 22652 2916 22704 2922
rect 22652 2858 22704 2864
rect 22744 2916 22796 2922
rect 22744 2858 22796 2864
rect 22756 2582 22784 2858
rect 23032 2774 23060 5102
rect 23112 4616 23164 4622
rect 23112 4558 23164 4564
rect 23124 4282 23152 4558
rect 23112 4276 23164 4282
rect 23112 4218 23164 4224
rect 23204 4208 23256 4214
rect 23204 4150 23256 4156
rect 23216 3058 23244 4150
rect 23204 3052 23256 3058
rect 23204 2994 23256 3000
rect 23308 2802 23336 5879
rect 23400 4298 23428 6870
rect 23572 4548 23624 4554
rect 23572 4490 23624 4496
rect 23584 4434 23612 4490
rect 23676 4434 23704 10254
rect 23846 10024 23902 10033
rect 23846 9959 23902 9968
rect 23754 5128 23810 5137
rect 23754 5063 23810 5072
rect 23768 4622 23796 5063
rect 23860 4826 23888 9959
rect 23940 9580 23992 9586
rect 23940 9522 23992 9528
rect 23952 8090 23980 9522
rect 24032 9444 24084 9450
rect 24032 9386 24084 9392
rect 24044 8498 24072 9386
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 23940 8084 23992 8090
rect 23940 8026 23992 8032
rect 23848 4820 23900 4826
rect 23848 4762 23900 4768
rect 23756 4616 23808 4622
rect 23756 4558 23808 4564
rect 23584 4406 23704 4434
rect 23400 4270 23612 4298
rect 23676 4282 23704 4406
rect 23584 4146 23612 4270
rect 23664 4276 23716 4282
rect 23664 4218 23716 4224
rect 23572 4140 23624 4146
rect 23572 4082 23624 4088
rect 23388 3936 23440 3942
rect 23386 3904 23388 3913
rect 23440 3904 23442 3913
rect 23386 3839 23442 3848
rect 23388 3664 23440 3670
rect 23386 3632 23388 3641
rect 23440 3632 23442 3641
rect 23386 3567 23442 3576
rect 23584 3534 23612 4082
rect 23572 3528 23624 3534
rect 23572 3470 23624 3476
rect 24032 3460 24084 3466
rect 24032 3402 24084 3408
rect 23572 3392 23624 3398
rect 23572 3334 23624 3340
rect 23480 2848 23532 2854
rect 23308 2796 23480 2802
rect 23308 2790 23532 2796
rect 23308 2774 23520 2790
rect 22940 2746 23060 2774
rect 22744 2576 22796 2582
rect 22744 2518 22796 2524
rect 22652 2440 22704 2446
rect 22652 2382 22704 2388
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 22376 2100 22428 2106
rect 22376 2042 22428 2048
rect 22098 1728 22154 1737
rect 22098 1663 22154 1672
rect 22572 800 22600 2246
rect 22664 1698 22692 2382
rect 22652 1692 22704 1698
rect 22652 1634 22704 1640
rect 22940 1630 22968 2746
rect 23388 2576 23440 2582
rect 23386 2544 23388 2553
rect 23440 2544 23442 2553
rect 23386 2479 23442 2488
rect 23584 1873 23612 3334
rect 24044 2825 24072 3402
rect 24030 2816 24086 2825
rect 24030 2751 24086 2760
rect 24136 2514 24164 11698
rect 24688 10674 24716 13903
rect 24676 10668 24728 10674
rect 24676 10610 24728 10616
rect 24872 9450 24900 15506
rect 25148 11121 25176 18226
rect 26240 18080 26292 18086
rect 26240 18022 26292 18028
rect 26148 16652 26200 16658
rect 26148 16594 26200 16600
rect 26160 16250 26188 16594
rect 26148 16244 26200 16250
rect 26148 16186 26200 16192
rect 26252 15978 26280 18022
rect 26240 15972 26292 15978
rect 26240 15914 26292 15920
rect 27080 15502 27108 21490
rect 27804 21344 27856 21350
rect 27804 21286 27856 21292
rect 27816 20466 27844 21286
rect 27804 20460 27856 20466
rect 27804 20402 27856 20408
rect 27252 19712 27304 19718
rect 27252 19654 27304 19660
rect 27264 18358 27292 19654
rect 27712 19372 27764 19378
rect 27712 19314 27764 19320
rect 27344 18624 27396 18630
rect 27344 18566 27396 18572
rect 27252 18352 27304 18358
rect 27252 18294 27304 18300
rect 27160 18216 27212 18222
rect 27160 18158 27212 18164
rect 27172 17338 27200 18158
rect 27160 17332 27212 17338
rect 27160 17274 27212 17280
rect 27264 17134 27292 18294
rect 27356 18290 27384 18566
rect 27344 18284 27396 18290
rect 27344 18226 27396 18232
rect 27344 17536 27396 17542
rect 27344 17478 27396 17484
rect 27356 17202 27384 17478
rect 27344 17196 27396 17202
rect 27344 17138 27396 17144
rect 27252 17128 27304 17134
rect 27252 17070 27304 17076
rect 27620 16992 27672 16998
rect 27620 16934 27672 16940
rect 27632 16590 27660 16934
rect 27620 16584 27672 16590
rect 27620 16526 27672 16532
rect 27632 16114 27660 16526
rect 27620 16108 27672 16114
rect 27620 16050 27672 16056
rect 27068 15496 27120 15502
rect 27068 15438 27120 15444
rect 25964 14952 26016 14958
rect 25964 14894 26016 14900
rect 25976 14482 26004 14894
rect 26148 14816 26200 14822
rect 26148 14758 26200 14764
rect 26056 14612 26108 14618
rect 26056 14554 26108 14560
rect 25964 14476 26016 14482
rect 25964 14418 26016 14424
rect 26068 13394 26096 14554
rect 26160 14482 26188 14758
rect 26148 14476 26200 14482
rect 26148 14418 26200 14424
rect 27080 14414 27108 15438
rect 27068 14408 27120 14414
rect 27068 14350 27120 14356
rect 26424 13456 26476 13462
rect 26424 13398 26476 13404
rect 26056 13388 26108 13394
rect 26056 13330 26108 13336
rect 26436 12434 26464 13398
rect 27080 13297 27108 14350
rect 27528 13320 27580 13326
rect 27066 13288 27122 13297
rect 27528 13262 27580 13268
rect 27066 13223 27122 13232
rect 27540 12986 27568 13262
rect 27724 13190 27752 19314
rect 28000 18766 28028 21490
rect 31128 20330 31156 24006
rect 32692 23866 32720 24754
rect 32680 23860 32732 23866
rect 32680 23802 32732 23808
rect 32876 23730 32904 35866
rect 33152 31346 33180 36586
rect 33232 36100 33284 36106
rect 33232 36042 33284 36048
rect 33244 33114 33272 36042
rect 33232 33108 33284 33114
rect 33232 33050 33284 33056
rect 33140 31340 33192 31346
rect 33140 31282 33192 31288
rect 34520 26512 34572 26518
rect 34520 26454 34572 26460
rect 34532 24206 34560 26454
rect 34520 24200 34572 24206
rect 34520 24142 34572 24148
rect 32864 23724 32916 23730
rect 32864 23666 32916 23672
rect 34808 22506 34836 37198
rect 35452 36786 35480 39200
rect 36096 37262 36124 39200
rect 37186 38856 37242 38865
rect 37186 38791 37242 38800
rect 36084 37256 36136 37262
rect 36084 37198 36136 37204
rect 36360 37120 36412 37126
rect 36360 37062 36412 37068
rect 35440 36780 35492 36786
rect 35440 36722 35492 36728
rect 35532 36576 35584 36582
rect 35532 36518 35584 36524
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35544 31822 35572 36518
rect 35532 31816 35584 31822
rect 35532 31758 35584 31764
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34796 22500 34848 22506
rect 34796 22442 34848 22448
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 31392 21548 31444 21554
rect 31392 21490 31444 21496
rect 31404 21146 31432 21490
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 31392 21140 31444 21146
rect 31392 21082 31444 21088
rect 35348 20868 35400 20874
rect 35348 20810 35400 20816
rect 35360 20466 35388 20810
rect 35348 20460 35400 20466
rect 35348 20402 35400 20408
rect 31116 20324 31168 20330
rect 31116 20266 31168 20272
rect 34796 20256 34848 20262
rect 34796 20198 34848 20204
rect 34520 19848 34572 19854
rect 34520 19790 34572 19796
rect 27988 18760 28040 18766
rect 27988 18702 28040 18708
rect 34532 18698 34560 19790
rect 34520 18692 34572 18698
rect 34520 18634 34572 18640
rect 28264 17672 28316 17678
rect 28264 17614 28316 17620
rect 28276 17338 28304 17614
rect 30564 17604 30616 17610
rect 30564 17546 30616 17552
rect 28264 17332 28316 17338
rect 28264 17274 28316 17280
rect 28448 17196 28500 17202
rect 28448 17138 28500 17144
rect 28460 16182 28488 17138
rect 28632 16516 28684 16522
rect 28632 16458 28684 16464
rect 28448 16176 28500 16182
rect 28448 16118 28500 16124
rect 28540 16176 28592 16182
rect 28540 16118 28592 16124
rect 28552 15570 28580 16118
rect 28540 15564 28592 15570
rect 28540 15506 28592 15512
rect 27988 15360 28040 15366
rect 27988 15302 28040 15308
rect 28000 15026 28028 15302
rect 27988 15020 28040 15026
rect 27988 14962 28040 14968
rect 27712 13184 27764 13190
rect 27712 13126 27764 13132
rect 27528 12980 27580 12986
rect 27528 12922 27580 12928
rect 28356 12844 28408 12850
rect 28356 12786 28408 12792
rect 26252 12406 26464 12434
rect 26252 12102 26280 12406
rect 28368 12238 28396 12786
rect 28356 12232 28408 12238
rect 28356 12174 28408 12180
rect 26240 12096 26292 12102
rect 26240 12038 26292 12044
rect 25964 11620 26016 11626
rect 25964 11562 26016 11568
rect 25134 11112 25190 11121
rect 25134 11047 25190 11056
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 24964 9654 24992 9862
rect 24952 9648 25004 9654
rect 24952 9590 25004 9596
rect 25044 9648 25096 9654
rect 25044 9590 25096 9596
rect 24860 9444 24912 9450
rect 24860 9386 24912 9392
rect 25056 9110 25084 9590
rect 25044 9104 25096 9110
rect 25044 9046 25096 9052
rect 24584 8968 24636 8974
rect 24584 8910 24636 8916
rect 24596 8401 24624 8910
rect 25228 8900 25280 8906
rect 25228 8842 25280 8848
rect 25240 8498 25268 8842
rect 25228 8492 25280 8498
rect 25228 8434 25280 8440
rect 24582 8392 24638 8401
rect 24582 8327 24638 8336
rect 25320 8356 25372 8362
rect 25320 8298 25372 8304
rect 24676 8288 24728 8294
rect 24676 8230 24728 8236
rect 24688 7818 24716 8230
rect 25332 7857 25360 8298
rect 25318 7848 25374 7857
rect 24676 7812 24728 7818
rect 25318 7783 25374 7792
rect 24676 7754 24728 7760
rect 24584 7744 24636 7750
rect 24584 7686 24636 7692
rect 24596 7410 24624 7686
rect 25976 7546 26004 11562
rect 26252 11150 26280 12038
rect 26240 11144 26292 11150
rect 26240 11086 26292 11092
rect 26148 11076 26200 11082
rect 26148 11018 26200 11024
rect 26056 10464 26108 10470
rect 26056 10406 26108 10412
rect 25964 7540 26016 7546
rect 25964 7482 26016 7488
rect 24584 7404 24636 7410
rect 24584 7346 24636 7352
rect 24492 5908 24544 5914
rect 24492 5850 24544 5856
rect 24400 4616 24452 4622
rect 24400 4558 24452 4564
rect 24412 4282 24440 4558
rect 24400 4276 24452 4282
rect 24400 4218 24452 4224
rect 24412 3398 24440 4218
rect 24400 3392 24452 3398
rect 24400 3334 24452 3340
rect 24504 2854 24532 5850
rect 25228 5568 25280 5574
rect 25228 5510 25280 5516
rect 24674 4584 24730 4593
rect 24674 4519 24730 4528
rect 24582 4176 24638 4185
rect 24688 4146 24716 4519
rect 24582 4111 24638 4120
rect 24676 4140 24728 4146
rect 24596 3738 24624 4111
rect 24676 4082 24728 4088
rect 25240 3738 25268 5510
rect 26068 4298 26096 10406
rect 26160 5302 26188 11018
rect 26238 7984 26294 7993
rect 26238 7919 26240 7928
rect 26292 7919 26294 7928
rect 26240 7890 26292 7896
rect 27160 7404 27212 7410
rect 27160 7346 27212 7352
rect 26424 5568 26476 5574
rect 26424 5510 26476 5516
rect 26148 5296 26200 5302
rect 26148 5238 26200 5244
rect 26436 5234 26464 5510
rect 26424 5228 26476 5234
rect 26424 5170 26476 5176
rect 26068 4270 26188 4298
rect 26056 4140 26108 4146
rect 26056 4082 26108 4088
rect 25780 4004 25832 4010
rect 25780 3946 25832 3952
rect 25320 3936 25372 3942
rect 25320 3878 25372 3884
rect 24584 3732 24636 3738
rect 24584 3674 24636 3680
rect 25228 3732 25280 3738
rect 25228 3674 25280 3680
rect 24676 3528 24728 3534
rect 24596 3488 24676 3516
rect 24596 3058 24624 3488
rect 24676 3470 24728 3476
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 24492 2848 24544 2854
rect 24492 2790 24544 2796
rect 24124 2508 24176 2514
rect 24124 2450 24176 2456
rect 24596 2446 24624 2994
rect 25228 2644 25280 2650
rect 25228 2586 25280 2592
rect 25240 2446 25268 2586
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 24676 2304 24728 2310
rect 24676 2246 24728 2252
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 24688 1902 24716 2246
rect 24676 1896 24728 1902
rect 23570 1864 23626 1873
rect 24676 1838 24728 1844
rect 23570 1799 23626 1808
rect 23848 1692 23900 1698
rect 23848 1634 23900 1640
rect 22928 1624 22980 1630
rect 22928 1566 22980 1572
rect 23860 800 23888 1634
rect 25148 800 25176 2246
rect 25332 2038 25360 3878
rect 25792 3534 25820 3946
rect 25780 3528 25832 3534
rect 25780 3470 25832 3476
rect 25412 3052 25464 3058
rect 25412 2994 25464 3000
rect 25320 2032 25372 2038
rect 25320 1974 25372 1980
rect 25424 1698 25452 2994
rect 25872 2916 25924 2922
rect 25872 2858 25924 2864
rect 25884 2446 25912 2858
rect 25872 2440 25924 2446
rect 25872 2382 25924 2388
rect 25780 2304 25832 2310
rect 25780 2246 25832 2252
rect 25412 1692 25464 1698
rect 25412 1634 25464 1640
rect 25792 800 25820 2246
rect 26068 2009 26096 4082
rect 26160 3466 26188 4270
rect 26148 3460 26200 3466
rect 26148 3402 26200 3408
rect 26240 3392 26292 3398
rect 26240 3334 26292 3340
rect 26252 3058 26280 3334
rect 27172 3194 27200 7346
rect 27804 4616 27856 4622
rect 27804 4558 27856 4564
rect 27436 3936 27488 3942
rect 27436 3878 27488 3884
rect 27252 3664 27304 3670
rect 27252 3606 27304 3612
rect 27160 3188 27212 3194
rect 27160 3130 27212 3136
rect 27264 3126 27292 3606
rect 27252 3120 27304 3126
rect 27252 3062 27304 3068
rect 26240 3052 26292 3058
rect 26240 2994 26292 3000
rect 27448 2582 27476 3878
rect 27816 2650 27844 4558
rect 28644 2650 28672 16458
rect 28724 16108 28776 16114
rect 28724 16050 28776 16056
rect 28736 11898 28764 16050
rect 30380 16040 30432 16046
rect 30380 15982 30432 15988
rect 29736 15904 29788 15910
rect 29736 15846 29788 15852
rect 29748 15502 29776 15846
rect 29736 15496 29788 15502
rect 29736 15438 29788 15444
rect 30392 13326 30420 15982
rect 30380 13320 30432 13326
rect 30380 13262 30432 13268
rect 28724 11892 28776 11898
rect 28724 11834 28776 11840
rect 30012 9376 30064 9382
rect 30012 9318 30064 9324
rect 30024 8634 30052 9318
rect 30012 8628 30064 8634
rect 30012 8570 30064 8576
rect 30104 7336 30156 7342
rect 30104 7278 30156 7284
rect 29460 5024 29512 5030
rect 29460 4966 29512 4972
rect 27804 2644 27856 2650
rect 27804 2586 27856 2592
rect 28632 2644 28684 2650
rect 28632 2586 28684 2592
rect 27436 2576 27488 2582
rect 27436 2518 27488 2524
rect 29472 2446 29500 4966
rect 30116 2650 30144 7278
rect 30576 2922 30604 17546
rect 31392 9580 31444 9586
rect 31392 9522 31444 9528
rect 30748 7880 30800 7886
rect 30748 7822 30800 7828
rect 30654 6216 30710 6225
rect 30654 6151 30656 6160
rect 30708 6151 30710 6160
rect 30656 6122 30708 6128
rect 30760 2990 30788 7822
rect 31404 4010 31432 9522
rect 33048 5024 33100 5030
rect 33048 4966 33100 4972
rect 31392 4004 31444 4010
rect 31392 3946 31444 3952
rect 30748 2984 30800 2990
rect 30748 2926 30800 2932
rect 30564 2916 30616 2922
rect 30564 2858 30616 2864
rect 30104 2644 30156 2650
rect 30104 2586 30156 2592
rect 33060 2446 33088 4966
rect 33600 3460 33652 3466
rect 33600 3402 33652 3408
rect 33612 3058 33640 3402
rect 33600 3052 33652 3058
rect 33600 2994 33652 3000
rect 33508 2848 33560 2854
rect 33508 2790 33560 2796
rect 27344 2440 27396 2446
rect 27158 2408 27214 2417
rect 27068 2372 27120 2378
rect 27344 2382 27396 2388
rect 29460 2440 29512 2446
rect 29460 2382 29512 2388
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 31576 2440 31628 2446
rect 31576 2382 31628 2388
rect 33048 2440 33100 2446
rect 33048 2382 33100 2388
rect 27158 2343 27214 2352
rect 27068 2314 27120 2320
rect 26054 2000 26110 2009
rect 26054 1935 26110 1944
rect 27080 800 27108 2314
rect 27172 2310 27200 2343
rect 27160 2304 27212 2310
rect 27160 2246 27212 2252
rect 27356 1766 27384 2382
rect 28356 2372 28408 2378
rect 28356 2314 28408 2320
rect 27344 1760 27396 1766
rect 27344 1702 27396 1708
rect 28368 800 28396 2314
rect 29644 2304 29696 2310
rect 29644 2246 29696 2252
rect 29656 800 29684 2246
rect 30300 800 30328 2382
rect 31588 800 31616 2382
rect 32864 2304 32916 2310
rect 32864 2246 32916 2252
rect 32876 800 32904 2246
rect 33520 800 33548 2790
rect 34808 2446 34836 20198
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 36372 18426 36400 37062
rect 37200 36378 37228 38791
rect 37384 37262 37412 39200
rect 38106 37496 38162 37505
rect 38106 37431 38162 37440
rect 37372 37256 37424 37262
rect 37372 37198 37424 37204
rect 37648 37120 37700 37126
rect 37648 37062 37700 37068
rect 37660 36718 37688 37062
rect 38120 36854 38148 37431
rect 38108 36848 38160 36854
rect 38108 36790 38160 36796
rect 37648 36712 37700 36718
rect 37648 36654 37700 36660
rect 38384 36644 38436 36650
rect 38384 36586 38436 36592
rect 37188 36372 37240 36378
rect 37188 36314 37240 36320
rect 38198 36136 38254 36145
rect 38198 36071 38254 36080
rect 38212 36038 38240 36071
rect 38200 36032 38252 36038
rect 38200 35974 38252 35980
rect 38108 35692 38160 35698
rect 38108 35634 38160 35640
rect 37648 35488 37700 35494
rect 38120 35465 38148 35634
rect 37648 35430 37700 35436
rect 38106 35456 38162 35465
rect 37280 34944 37332 34950
rect 37280 34886 37332 34892
rect 37292 30870 37320 34886
rect 37280 30864 37332 30870
rect 37280 30806 37332 30812
rect 37464 30728 37516 30734
rect 37462 30696 37464 30705
rect 37516 30696 37518 30705
rect 37462 30631 37518 30640
rect 37372 29640 37424 29646
rect 37372 29582 37424 29588
rect 37384 27606 37412 29582
rect 37464 28008 37516 28014
rect 37462 27976 37464 27985
rect 37516 27976 37518 27985
rect 37462 27911 37518 27920
rect 37372 27600 37424 27606
rect 37372 27542 37424 27548
rect 37556 27464 37608 27470
rect 37556 27406 37608 27412
rect 37568 27130 37596 27406
rect 37556 27124 37608 27130
rect 37556 27066 37608 27072
rect 37280 26988 37332 26994
rect 37280 26930 37332 26936
rect 36820 20460 36872 20466
rect 36820 20402 36872 20408
rect 36832 19514 36860 20402
rect 36820 19508 36872 19514
rect 36820 19450 36872 19456
rect 36360 18420 36412 18426
rect 36360 18362 36412 18368
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 37292 16114 37320 26930
rect 37372 21616 37424 21622
rect 37372 21558 37424 21564
rect 37384 20942 37412 21558
rect 37372 20936 37424 20942
rect 37372 20878 37424 20884
rect 37280 16108 37332 16114
rect 37280 16050 37332 16056
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 37280 14476 37332 14482
rect 37280 14418 37332 14424
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 37292 13326 37320 14418
rect 37280 13320 37332 13326
rect 37280 13262 37332 13268
rect 36912 13184 36964 13190
rect 36912 13126 36964 13132
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 36924 10062 36952 13126
rect 37384 11218 37412 20878
rect 37464 18760 37516 18766
rect 37464 18702 37516 18708
rect 37476 16574 37504 18702
rect 37476 16546 37596 16574
rect 37372 11212 37424 11218
rect 37372 11154 37424 11160
rect 37188 11144 37240 11150
rect 37188 11086 37240 11092
rect 37200 10985 37228 11086
rect 37186 10976 37242 10985
rect 37186 10911 37242 10920
rect 36912 10056 36964 10062
rect 36912 9998 36964 10004
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 37464 7880 37516 7886
rect 37464 7822 37516 7828
rect 37476 7585 37504 7822
rect 37462 7576 37518 7585
rect 37462 7511 37518 7520
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 37568 6914 37596 16546
rect 37660 13530 37688 35430
rect 38106 35391 38162 35400
rect 38200 34400 38252 34406
rect 38200 34342 38252 34348
rect 38212 34105 38240 34342
rect 38198 34096 38254 34105
rect 38198 34031 38254 34040
rect 38108 32836 38160 32842
rect 38108 32778 38160 32784
rect 38120 32745 38148 32778
rect 38200 32768 38252 32774
rect 38106 32736 38162 32745
rect 38200 32710 38252 32716
rect 38106 32671 38162 32680
rect 38108 32428 38160 32434
rect 38108 32370 38160 32376
rect 37924 32224 37976 32230
rect 37924 32166 37976 32172
rect 37832 28008 37884 28014
rect 37832 27950 37884 27956
rect 37740 24200 37792 24206
rect 37740 24142 37792 24148
rect 37752 20602 37780 24142
rect 37844 23118 37872 27950
rect 37832 23112 37884 23118
rect 37832 23054 37884 23060
rect 37844 22778 37872 23054
rect 37832 22772 37884 22778
rect 37832 22714 37884 22720
rect 37832 22636 37884 22642
rect 37832 22578 37884 22584
rect 37740 20596 37792 20602
rect 37740 20538 37792 20544
rect 37844 19514 37872 22578
rect 37936 22574 37964 32166
rect 38120 32065 38148 32370
rect 38106 32056 38162 32065
rect 38106 31991 38162 32000
rect 38212 29594 38240 32710
rect 38120 29566 38240 29594
rect 38016 27464 38068 27470
rect 38016 27406 38068 27412
rect 38028 25498 38056 27406
rect 38016 25492 38068 25498
rect 38016 25434 38068 25440
rect 38016 22772 38068 22778
rect 38016 22714 38068 22720
rect 37924 22568 37976 22574
rect 37924 22510 37976 22516
rect 38028 22030 38056 22714
rect 38016 22024 38068 22030
rect 38016 21966 38068 21972
rect 37924 21888 37976 21894
rect 37924 21830 37976 21836
rect 37832 19508 37884 19514
rect 37832 19450 37884 19456
rect 37832 17536 37884 17542
rect 37832 17478 37884 17484
rect 37648 13524 37700 13530
rect 37648 13466 37700 13472
rect 37740 9988 37792 9994
rect 37740 9930 37792 9936
rect 37752 7954 37780 9930
rect 37740 7948 37792 7954
rect 37740 7890 37792 7896
rect 37476 6886 37596 6914
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 37476 3738 37504 6886
rect 37752 4622 37780 7890
rect 37844 6914 37872 17478
rect 37936 14414 37964 21830
rect 38016 20936 38068 20942
rect 38016 20878 38068 20884
rect 38028 20058 38056 20878
rect 38120 20534 38148 29566
rect 38200 29504 38252 29510
rect 38200 29446 38252 29452
rect 38212 29345 38240 29446
rect 38198 29336 38254 29345
rect 38198 29271 38254 29280
rect 38200 27328 38252 27334
rect 38198 27296 38200 27305
rect 38252 27296 38254 27305
rect 38198 27231 38254 27240
rect 38292 26376 38344 26382
rect 38292 26318 38344 26324
rect 38304 25945 38332 26318
rect 38290 25936 38346 25945
rect 38290 25871 38346 25880
rect 38200 24608 38252 24614
rect 38198 24576 38200 24585
rect 38252 24576 38254 24585
rect 38198 24511 38254 24520
rect 38200 24064 38252 24070
rect 38200 24006 38252 24012
rect 38212 23905 38240 24006
rect 38198 23896 38254 23905
rect 38198 23831 38254 23840
rect 38198 22536 38254 22545
rect 38198 22471 38200 22480
rect 38252 22471 38254 22480
rect 38200 22442 38252 22448
rect 38200 21344 38252 21350
rect 38200 21286 38252 21292
rect 38212 21185 38240 21286
rect 38198 21176 38254 21185
rect 38198 21111 38254 21120
rect 38396 21010 38424 36586
rect 38476 36236 38528 36242
rect 38476 36178 38528 36184
rect 38488 21146 38516 36178
rect 38672 35086 38700 39200
rect 39316 36786 39344 39200
rect 39304 36780 39356 36786
rect 39304 36722 39356 36728
rect 38660 35080 38712 35086
rect 38660 35022 38712 35028
rect 38568 34604 38620 34610
rect 38568 34546 38620 34552
rect 38476 21140 38528 21146
rect 38476 21082 38528 21088
rect 38384 21004 38436 21010
rect 38384 20946 38436 20952
rect 38200 20800 38252 20806
rect 38200 20742 38252 20748
rect 38108 20528 38160 20534
rect 38212 20505 38240 20742
rect 38108 20470 38160 20476
rect 38198 20496 38254 20505
rect 38198 20431 38254 20440
rect 38016 20052 38068 20058
rect 38016 19994 38068 20000
rect 38016 19372 38068 19378
rect 38016 19314 38068 19320
rect 38028 18426 38056 19314
rect 38290 19136 38346 19145
rect 38290 19071 38346 19080
rect 38200 18896 38252 18902
rect 38200 18838 38252 18844
rect 38108 18624 38160 18630
rect 38108 18566 38160 18572
rect 38016 18420 38068 18426
rect 38016 18362 38068 18368
rect 38120 18290 38148 18566
rect 38108 18284 38160 18290
rect 38108 18226 38160 18232
rect 38016 16584 38068 16590
rect 38212 16574 38240 18838
rect 38304 18766 38332 19071
rect 38580 18970 38608 34546
rect 38568 18964 38620 18970
rect 38568 18906 38620 18912
rect 38292 18760 38344 18766
rect 38292 18702 38344 18708
rect 38292 18284 38344 18290
rect 38292 18226 38344 18232
rect 38304 17785 38332 18226
rect 38290 17776 38346 17785
rect 38290 17711 38346 17720
rect 38212 16546 38424 16574
rect 38016 16526 38068 16532
rect 38028 16046 38056 16526
rect 38200 16448 38252 16454
rect 38198 16416 38200 16425
rect 38252 16416 38254 16425
rect 38198 16351 38254 16360
rect 38292 16108 38344 16114
rect 38292 16050 38344 16056
rect 38016 16040 38068 16046
rect 38016 15982 38068 15988
rect 38304 15745 38332 16050
rect 38290 15736 38346 15745
rect 38290 15671 38346 15680
rect 37924 14408 37976 14414
rect 37924 14350 37976 14356
rect 38198 14376 38254 14385
rect 38198 14311 38254 14320
rect 38212 14278 38240 14311
rect 38200 14272 38252 14278
rect 38200 14214 38252 14220
rect 38200 13184 38252 13190
rect 38200 13126 38252 13132
rect 38212 13025 38240 13126
rect 38198 13016 38254 13025
rect 38198 12951 38254 12960
rect 38108 12844 38160 12850
rect 38108 12786 38160 12792
rect 38120 12345 38148 12786
rect 38198 12744 38254 12753
rect 38198 12679 38254 12688
rect 38212 12646 38240 12679
rect 38200 12640 38252 12646
rect 38200 12582 38252 12588
rect 38106 12336 38162 12345
rect 38106 12271 38162 12280
rect 38200 9920 38252 9926
rect 38200 9862 38252 9868
rect 38212 9625 38240 9862
rect 38198 9616 38254 9625
rect 38198 9551 38254 9560
rect 38396 8566 38424 16546
rect 38384 8560 38436 8566
rect 38384 8502 38436 8508
rect 38108 8492 38160 8498
rect 38108 8434 38160 8440
rect 38120 8265 38148 8434
rect 38106 8256 38162 8265
rect 38106 8191 38162 8200
rect 37844 6886 37964 6914
rect 37936 5234 37964 6886
rect 38292 6316 38344 6322
rect 38292 6258 38344 6264
rect 38304 6225 38332 6258
rect 38290 6216 38346 6225
rect 38290 6151 38346 6160
rect 37924 5228 37976 5234
rect 37924 5170 37976 5176
rect 38108 5160 38160 5166
rect 38108 5102 38160 5108
rect 37740 4616 37792 4622
rect 37740 4558 37792 4564
rect 38016 4480 38068 4486
rect 38016 4422 38068 4428
rect 37464 3732 37516 3738
rect 37464 3674 37516 3680
rect 37648 3528 37700 3534
rect 37648 3470 37700 3476
rect 36728 3120 36780 3126
rect 36728 3062 36780 3068
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 34796 2304 34848 2310
rect 34796 2246 34848 2252
rect 36084 2304 36136 2310
rect 36084 2246 36136 2252
rect 34808 800 34836 2246
rect 36096 800 36124 2246
rect 36740 800 36768 3062
rect 36912 3052 36964 3058
rect 36912 2994 36964 3000
rect 36924 1465 36952 2994
rect 36910 1456 36966 1465
rect 36910 1391 36966 1400
rect 1674 776 1730 785
rect 1674 711 1730 720
rect 1950 200 2006 800
rect 3238 200 3294 800
rect 3882 200 3938 800
rect 5170 200 5226 800
rect 6458 200 6514 800
rect 7102 200 7158 800
rect 8390 200 8446 800
rect 9678 200 9734 800
rect 10966 200 11022 800
rect 11610 200 11666 800
rect 12898 200 12954 800
rect 14186 200 14242 800
rect 14830 200 14886 800
rect 16118 200 16174 800
rect 17406 200 17462 800
rect 18050 200 18106 800
rect 19338 200 19394 800
rect 20626 200 20682 800
rect 21914 200 21970 800
rect 22558 200 22614 800
rect 23846 200 23902 800
rect 25134 200 25190 800
rect 25778 200 25834 800
rect 27066 200 27122 800
rect 28354 200 28410 800
rect 29642 200 29698 800
rect 30286 200 30342 800
rect 31574 200 31630 800
rect 32862 200 32918 800
rect 33506 200 33562 800
rect 34794 200 34850 800
rect 36082 200 36138 800
rect 36726 200 36782 800
rect 37660 785 37688 3470
rect 38028 2446 38056 4422
rect 38120 3738 38148 5102
rect 38200 5024 38252 5030
rect 38200 4966 38252 4972
rect 38212 4865 38240 4966
rect 38198 4856 38254 4865
rect 38198 4791 38254 4800
rect 38290 4176 38346 4185
rect 38290 4111 38292 4120
rect 38344 4111 38346 4120
rect 38292 4082 38344 4088
rect 38108 3732 38160 3738
rect 38108 3674 38160 3680
rect 38108 3528 38160 3534
rect 38108 3470 38160 3476
rect 38016 2440 38068 2446
rect 38016 2382 38068 2388
rect 38120 1986 38148 3470
rect 38292 3052 38344 3058
rect 38292 2994 38344 3000
rect 38304 2825 38332 2994
rect 38290 2816 38346 2825
rect 38290 2751 38346 2760
rect 39304 2304 39356 2310
rect 39304 2246 39356 2252
rect 38028 1958 38148 1986
rect 38028 800 38056 1958
rect 39316 800 39344 2246
rect 37646 776 37702 785
rect 37646 711 37702 720
rect 38014 200 38070 800
rect 39302 200 39358 800
<< via2 >>
rect 1766 38800 1822 38856
rect 1674 38120 1730 38176
rect 1582 35400 1638 35456
rect 1766 34720 1822 34776
rect 1766 33380 1822 33416
rect 1766 33360 1768 33380
rect 1768 33360 1820 33380
rect 1820 33360 1822 33380
rect 1766 32000 1822 32056
rect 1582 31320 1638 31376
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 2502 36780 2558 36816
rect 2502 36760 2504 36780
rect 2504 36760 2556 36780
rect 2556 36760 2558 36780
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 1766 29996 1768 30016
rect 1768 29996 1820 30016
rect 1820 29996 1822 30016
rect 1766 29960 1822 29996
rect 1582 29028 1638 29064
rect 1582 29008 1584 29028
rect 1584 29008 1636 29028
rect 1636 29008 1638 29028
rect 1766 28600 1822 28656
rect 846 17312 902 17368
rect 1398 24928 1454 24984
rect 1858 27648 1914 27704
rect 2042 27648 2098 27704
rect 1950 26696 2006 26752
rect 1858 26424 1914 26480
rect 1766 25200 1822 25256
rect 1766 23840 1822 23896
rect 1674 23160 1730 23216
rect 1398 7520 1454 7576
rect 1398 5480 1454 5536
rect 1766 21800 1822 21856
rect 2594 28076 2650 28112
rect 2594 28056 2596 28076
rect 2596 28056 2648 28076
rect 2648 28056 2650 28076
rect 2502 26832 2558 26888
rect 2502 26324 2504 26344
rect 2504 26324 2556 26344
rect 2556 26324 2558 26344
rect 2502 26288 2558 26324
rect 2778 26152 2834 26208
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 3238 27820 3240 27840
rect 3240 27820 3292 27840
rect 3292 27820 3294 27840
rect 3238 27784 3294 27820
rect 2226 25236 2228 25256
rect 2228 25236 2280 25256
rect 2280 25236 2282 25256
rect 2226 25200 2282 25236
rect 1858 19216 1914 19272
rect 1858 17448 1914 17504
rect 2134 19216 2190 19272
rect 2502 24012 2504 24032
rect 2504 24012 2556 24032
rect 2556 24012 2558 24032
rect 2502 23976 2558 24012
rect 2226 16360 2282 16416
rect 1582 8628 1638 8664
rect 1582 8608 1584 8628
rect 1584 8608 1636 8628
rect 1636 8608 1638 8628
rect 1858 7268 1914 7304
rect 1858 7248 1860 7268
rect 1860 7248 1912 7268
rect 1912 7248 1914 7268
rect 2226 14864 2282 14920
rect 2318 14320 2374 14376
rect 2686 22480 2742 22536
rect 2502 18944 2558 19000
rect 2870 19216 2926 19272
rect 3422 26560 3478 26616
rect 3422 23432 3478 23488
rect 3606 23432 3662 23488
rect 3330 20340 3332 20360
rect 3332 20340 3384 20360
rect 3384 20340 3386 20360
rect 3330 20304 3386 20340
rect 3054 18400 3110 18456
rect 2778 17040 2834 17096
rect 2870 16360 2926 16416
rect 2778 15680 2834 15736
rect 2778 13640 2834 13696
rect 2778 11600 2834 11656
rect 3146 16632 3202 16688
rect 3330 15952 3386 16008
rect 3698 20440 3754 20496
rect 3514 16224 3570 16280
rect 3698 19352 3754 19408
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4066 27240 4122 27296
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4618 26288 4674 26344
rect 3882 24928 3938 24984
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 3974 24148 3976 24168
rect 3976 24148 4028 24168
rect 4028 24148 4030 24168
rect 4802 24792 4858 24848
rect 3974 24112 4030 24148
rect 4802 24148 4804 24168
rect 4804 24148 4856 24168
rect 4856 24148 4858 24168
rect 3882 23860 3938 23896
rect 3882 23840 3884 23860
rect 3884 23840 3936 23860
rect 3936 23840 3938 23860
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4802 24112 4858 24148
rect 4710 23568 4766 23624
rect 3974 20440 4030 20496
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4342 21664 4398 21720
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4158 20984 4214 21040
rect 4710 20712 4766 20768
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4618 19896 4674 19952
rect 4526 19216 4582 19272
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4250 18808 4306 18864
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4802 20576 4858 20632
rect 4802 20168 4858 20224
rect 5170 24928 5226 24984
rect 5170 24792 5226 24848
rect 4986 21936 5042 21992
rect 4894 19624 4950 19680
rect 3974 17584 4030 17640
rect 4250 17604 4306 17640
rect 4250 17584 4252 17604
rect 4252 17584 4304 17604
rect 4304 17584 4306 17604
rect 4526 17584 4582 17640
rect 4710 17720 4766 17776
rect 5262 22480 5318 22536
rect 5078 21800 5134 21856
rect 5078 20168 5134 20224
rect 5354 20032 5410 20088
rect 5170 19624 5226 19680
rect 5078 19488 5134 19544
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4066 16396 4068 16416
rect 4068 16396 4120 16416
rect 4120 16396 4122 16416
rect 4066 16360 4122 16396
rect 3514 15000 3570 15056
rect 3146 12280 3202 12336
rect 3422 11600 3478 11656
rect 3422 9424 3478 9480
rect 3974 15544 4030 15600
rect 4802 17312 4858 17368
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4066 15272 4122 15328
rect 3698 13776 3754 13832
rect 3698 12144 3754 12200
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4710 14728 4766 14784
rect 3974 13912 4030 13968
rect 3974 13252 4030 13288
rect 3974 13232 3976 13252
rect 3976 13232 4028 13252
rect 4028 13232 4030 13252
rect 3974 12688 4030 12744
rect 4618 14068 4674 14104
rect 4618 14048 4620 14068
rect 4620 14048 4672 14068
rect 4672 14048 4674 14068
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4342 13368 4398 13424
rect 4250 12724 4252 12744
rect 4252 12724 4304 12744
rect 4304 12724 4306 12744
rect 4250 12688 4306 12724
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 3790 10240 3846 10296
rect 1766 6876 1768 6896
rect 1768 6876 1820 6896
rect 1820 6876 1822 6896
rect 1766 6840 1822 6876
rect 1674 4156 1676 4176
rect 1676 4156 1728 4176
rect 1728 4156 1730 4176
rect 1674 4120 1730 4156
rect 2502 2080 2558 2136
rect 2686 1944 2742 2000
rect 3422 8084 3478 8120
rect 3422 8064 3424 8084
rect 3424 8064 3476 8084
rect 3476 8064 3478 8084
rect 3146 3340 3148 3360
rect 3148 3340 3200 3360
rect 3200 3340 3202 3360
rect 3146 3304 3202 3340
rect 2870 1808 2926 1864
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4618 11056 4674 11112
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4526 9832 4582 9888
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 3974 8880 4030 8936
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4066 5788 4068 5808
rect 4068 5788 4120 5808
rect 4120 5788 4122 5808
rect 4066 5752 4122 5788
rect 5262 18128 5318 18184
rect 5170 16088 5226 16144
rect 5078 14184 5134 14240
rect 5906 20168 5962 20224
rect 5538 16244 5594 16280
rect 5538 16224 5540 16244
rect 5540 16224 5592 16244
rect 5592 16224 5594 16244
rect 5814 16088 5870 16144
rect 5446 15544 5502 15600
rect 5538 15156 5594 15192
rect 5538 15136 5540 15156
rect 5540 15136 5592 15156
rect 5592 15136 5594 15156
rect 5538 14612 5594 14648
rect 5538 14592 5540 14612
rect 5540 14592 5592 14612
rect 5592 14592 5594 14612
rect 6182 17448 6238 17504
rect 6550 24792 6606 24848
rect 7194 25064 7250 25120
rect 7010 24928 7066 24984
rect 6734 22344 6790 22400
rect 6366 21936 6422 21992
rect 6366 21548 6422 21584
rect 6366 21528 6368 21548
rect 6368 21528 6420 21548
rect 6420 21528 6422 21548
rect 6458 20440 6514 20496
rect 6734 20168 6790 20224
rect 6826 19760 6882 19816
rect 6366 18708 6368 18728
rect 6368 18708 6420 18728
rect 6420 18708 6422 18728
rect 6366 18672 6422 18708
rect 5262 13640 5318 13696
rect 4986 12416 5042 12472
rect 4894 11192 4950 11248
rect 5630 12708 5686 12744
rect 5630 12688 5632 12708
rect 5632 12688 5684 12708
rect 5684 12688 5686 12708
rect 5446 10684 5448 10704
rect 5448 10684 5500 10704
rect 5500 10684 5502 10704
rect 5446 10648 5502 10684
rect 5538 9832 5594 9888
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4066 3440 4122 3496
rect 4342 3032 4398 3088
rect 4066 2916 4122 2952
rect 4066 2896 4068 2916
rect 4068 2896 4120 2916
rect 4120 2896 4122 2916
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 5538 2760 5594 2816
rect 5262 2624 5318 2680
rect 6274 13404 6276 13424
rect 6276 13404 6328 13424
rect 6328 13404 6330 13424
rect 6274 13368 6330 13404
rect 6642 19352 6698 19408
rect 6918 19352 6974 19408
rect 6550 15136 6606 15192
rect 6734 15580 6736 15600
rect 6736 15580 6788 15600
rect 6788 15580 6790 15600
rect 6734 15544 6790 15580
rect 6642 13776 6698 13832
rect 6642 11464 6698 11520
rect 7654 23840 7710 23896
rect 7470 23432 7526 23488
rect 7562 20440 7618 20496
rect 7470 19896 7526 19952
rect 7194 15308 7196 15328
rect 7196 15308 7248 15328
rect 7248 15308 7250 15328
rect 7194 15272 7250 15308
rect 7102 14476 7158 14512
rect 7102 14456 7104 14476
rect 7104 14456 7156 14476
rect 7156 14456 7158 14476
rect 6826 11772 6828 11792
rect 6828 11772 6880 11792
rect 6880 11772 6882 11792
rect 6826 11736 6882 11772
rect 6734 10512 6790 10568
rect 7746 23060 7748 23080
rect 7748 23060 7800 23080
rect 7800 23060 7802 23080
rect 7746 23024 7802 23060
rect 7746 19780 7802 19816
rect 7746 19760 7748 19780
rect 7748 19760 7800 19780
rect 7800 19760 7802 19780
rect 8114 21936 8170 21992
rect 7930 20340 7932 20360
rect 7932 20340 7984 20360
rect 7984 20340 7986 20360
rect 7930 20304 7986 20340
rect 7654 17856 7710 17912
rect 7470 16360 7526 16416
rect 7654 15000 7710 15056
rect 7562 12416 7618 12472
rect 8114 19352 8170 19408
rect 8390 23568 8446 23624
rect 8022 13912 8078 13968
rect 7102 8628 7158 8664
rect 7102 8608 7104 8628
rect 7104 8608 7156 8628
rect 7156 8608 7158 8628
rect 6918 5208 6974 5264
rect 6090 3304 6146 3360
rect 6642 3576 6698 3632
rect 8574 18944 8630 19000
rect 8390 15680 8446 15736
rect 9126 24792 9182 24848
rect 9678 24928 9734 24984
rect 8942 20868 8998 20904
rect 8942 20848 8944 20868
rect 8944 20848 8996 20868
rect 8996 20848 8998 20868
rect 8942 20032 8998 20088
rect 8758 19624 8814 19680
rect 8666 18264 8722 18320
rect 8758 17856 8814 17912
rect 8390 13368 8446 13424
rect 8206 12280 8262 12336
rect 8022 11600 8078 11656
rect 8298 10784 8354 10840
rect 8758 15952 8814 16008
rect 8850 13812 8852 13832
rect 8852 13812 8904 13832
rect 8904 13812 8906 13832
rect 8850 13776 8906 13812
rect 8758 13640 8814 13696
rect 9678 22072 9734 22128
rect 9402 21664 9458 21720
rect 9678 21004 9734 21040
rect 9678 20984 9680 21004
rect 9680 20984 9732 21004
rect 9732 20984 9734 21004
rect 9126 19896 9182 19952
rect 9310 20168 9366 20224
rect 9310 18672 9366 18728
rect 9678 20576 9734 20632
rect 9126 17312 9182 17368
rect 9218 16668 9220 16688
rect 9220 16668 9272 16688
rect 9272 16668 9274 16688
rect 9218 16632 9274 16668
rect 10230 23432 10286 23488
rect 10138 20868 10194 20904
rect 10138 20848 10140 20868
rect 10140 20848 10192 20868
rect 10192 20848 10194 20868
rect 10506 21528 10562 21584
rect 10046 19080 10102 19136
rect 9310 16532 9312 16552
rect 9312 16532 9364 16552
rect 9364 16532 9366 16552
rect 9310 16496 9366 16532
rect 9126 16360 9182 16416
rect 9310 15952 9366 16008
rect 9126 15700 9182 15736
rect 9126 15680 9128 15700
rect 9128 15680 9180 15700
rect 9180 15680 9182 15700
rect 9494 15156 9550 15192
rect 9494 15136 9496 15156
rect 9496 15136 9548 15156
rect 9548 15136 9550 15156
rect 9310 14728 9366 14784
rect 9310 14456 9366 14512
rect 9402 14320 9458 14376
rect 8942 11500 8944 11520
rect 8944 11500 8996 11520
rect 8996 11500 8998 11520
rect 8942 11464 8998 11500
rect 10046 18400 10102 18456
rect 10046 18164 10048 18184
rect 10048 18164 10100 18184
rect 10100 18164 10102 18184
rect 10046 18128 10102 18164
rect 10046 17720 10102 17776
rect 9954 13776 10010 13832
rect 9678 11600 9734 11656
rect 9310 11056 9366 11112
rect 7654 6704 7710 6760
rect 7746 4664 7802 4720
rect 7562 3440 7618 3496
rect 7286 3032 7342 3088
rect 7930 4548 7986 4584
rect 7930 4528 7932 4548
rect 7932 4528 7984 4548
rect 7984 4528 7986 4548
rect 8114 4392 8170 4448
rect 8390 5652 8392 5672
rect 8392 5652 8444 5672
rect 8444 5652 8446 5672
rect 8390 5616 8446 5652
rect 8390 3596 8446 3632
rect 8390 3576 8392 3596
rect 8392 3576 8444 3596
rect 8444 3576 8446 3596
rect 8666 5888 8722 5944
rect 9770 11328 9826 11384
rect 9678 10920 9734 10976
rect 9586 10512 9642 10568
rect 9586 9424 9642 9480
rect 10414 15680 10470 15736
rect 11058 21800 11114 21856
rect 10966 21392 11022 21448
rect 10874 21256 10930 21312
rect 10782 20460 10838 20496
rect 10782 20440 10784 20460
rect 10784 20440 10836 20460
rect 10836 20440 10838 20460
rect 10598 17856 10654 17912
rect 10690 17312 10746 17368
rect 10966 20984 11022 21040
rect 11150 19896 11206 19952
rect 10874 18400 10930 18456
rect 10874 17756 10876 17776
rect 10876 17756 10928 17776
rect 10928 17756 10930 17776
rect 10874 17720 10930 17756
rect 11150 17484 11152 17504
rect 11152 17484 11204 17504
rect 11204 17484 11206 17504
rect 11150 17448 11206 17484
rect 11150 17312 11206 17368
rect 10966 16632 11022 16688
rect 11150 15272 11206 15328
rect 10690 13932 10746 13968
rect 10690 13912 10692 13932
rect 10692 13912 10744 13932
rect 10744 13912 10746 13932
rect 10322 13776 10378 13832
rect 10782 13640 10838 13696
rect 10690 13368 10746 13424
rect 10230 12824 10286 12880
rect 9954 8900 10010 8936
rect 9954 8880 9956 8900
rect 9956 8880 10008 8900
rect 10008 8880 10010 8900
rect 9678 6996 9734 7032
rect 9862 7520 9918 7576
rect 9678 6976 9680 6996
rect 9680 6976 9732 6996
rect 9732 6976 9734 6996
rect 9678 6840 9734 6896
rect 9034 5344 9090 5400
rect 9310 4800 9366 4856
rect 8942 3984 8998 4040
rect 9586 4156 9588 4176
rect 9588 4156 9640 4176
rect 9640 4156 9642 4176
rect 9586 4120 9642 4156
rect 9402 3712 9458 3768
rect 10598 10512 10654 10568
rect 10506 6840 10562 6896
rect 10506 2488 10562 2544
rect 10966 12044 10968 12064
rect 10968 12044 11020 12064
rect 11020 12044 11022 12064
rect 10966 12008 11022 12044
rect 11426 26152 11482 26208
rect 11702 23568 11758 23624
rect 11334 14184 11390 14240
rect 11886 22072 11942 22128
rect 12162 22888 12218 22944
rect 12714 22924 12716 22944
rect 12716 22924 12768 22944
rect 12768 22924 12770 22944
rect 12714 22888 12770 22924
rect 12622 22072 12678 22128
rect 12254 21256 12310 21312
rect 11702 18944 11758 19000
rect 11886 16904 11942 16960
rect 12346 19080 12402 19136
rect 12346 18944 12402 19000
rect 12162 18536 12218 18592
rect 12714 21956 12770 21992
rect 12714 21936 12716 21956
rect 12716 21936 12768 21956
rect 12768 21936 12770 21956
rect 12806 21664 12862 21720
rect 12438 17584 12494 17640
rect 12346 16904 12402 16960
rect 11334 12280 11390 12336
rect 11702 14184 11758 14240
rect 12070 15564 12126 15600
rect 12070 15544 12072 15564
rect 12072 15544 12124 15564
rect 12124 15544 12126 15564
rect 12346 16768 12402 16824
rect 12254 16360 12310 16416
rect 12530 16496 12586 16552
rect 11426 11328 11482 11384
rect 11426 10376 11482 10432
rect 10966 9444 11022 9480
rect 10966 9424 10968 9444
rect 10968 9424 11020 9444
rect 11020 9424 11022 9444
rect 11426 9424 11482 9480
rect 10966 7420 10968 7440
rect 10968 7420 11020 7440
rect 11020 7420 11022 7440
rect 10966 7384 11022 7420
rect 10782 7112 10838 7168
rect 11150 6976 11206 7032
rect 10874 2624 10930 2680
rect 11702 9832 11758 9888
rect 12990 19488 13046 19544
rect 13358 20868 13414 20904
rect 13358 20848 13360 20868
rect 13360 20848 13412 20868
rect 13412 20848 13414 20868
rect 13542 21020 13544 21040
rect 13544 21020 13596 21040
rect 13596 21020 13598 21040
rect 13542 20984 13598 21020
rect 12898 15680 12954 15736
rect 13082 18264 13138 18320
rect 13082 17856 13138 17912
rect 13358 17176 13414 17232
rect 12806 15408 12862 15464
rect 12530 13640 12586 13696
rect 12714 13504 12770 13560
rect 12346 13096 12402 13152
rect 12438 12824 12494 12880
rect 13266 16224 13322 16280
rect 13174 15272 13230 15328
rect 13082 12860 13084 12880
rect 13084 12860 13136 12880
rect 13136 12860 13138 12880
rect 13082 12824 13138 12860
rect 12070 11600 12126 11656
rect 12438 11600 12494 11656
rect 11978 11464 12034 11520
rect 12162 11464 12218 11520
rect 12438 11464 12494 11520
rect 11886 10512 11942 10568
rect 11610 5344 11666 5400
rect 11334 3848 11390 3904
rect 10966 2352 11022 2408
rect 12162 10512 12218 10568
rect 12162 10376 12218 10432
rect 12346 10376 12402 10432
rect 12622 11872 12678 11928
rect 13266 12688 13322 12744
rect 13174 12552 13230 12608
rect 13174 12416 13230 12472
rect 12438 9968 12494 10024
rect 12346 9832 12402 9888
rect 12254 6568 12310 6624
rect 13266 12044 13268 12064
rect 13268 12044 13320 12064
rect 13320 12044 13322 12064
rect 13266 12008 13322 12044
rect 13634 18536 13690 18592
rect 13542 18400 13598 18456
rect 13634 18128 13690 18184
rect 13726 17312 13782 17368
rect 13726 15408 13782 15464
rect 13450 13368 13506 13424
rect 13634 12724 13636 12744
rect 13636 12724 13688 12744
rect 13688 12724 13690 12744
rect 13634 12688 13690 12724
rect 13542 12436 13598 12472
rect 13542 12416 13544 12436
rect 13544 12416 13596 12436
rect 13596 12416 13598 12436
rect 13818 11328 13874 11384
rect 13450 6976 13506 7032
rect 13174 6840 13230 6896
rect 13726 9036 13782 9072
rect 13726 9016 13728 9036
rect 13728 9016 13780 9036
rect 13780 9016 13782 9036
rect 13634 8472 13690 8528
rect 14370 26324 14372 26344
rect 14372 26324 14424 26344
rect 14424 26324 14426 26344
rect 14370 26288 14426 26324
rect 14278 20712 14334 20768
rect 14370 19624 14426 19680
rect 15014 21800 15070 21856
rect 14738 18944 14794 19000
rect 14278 16940 14280 16960
rect 14280 16940 14332 16960
rect 14332 16940 14334 16960
rect 14278 16904 14334 16940
rect 14462 15816 14518 15872
rect 14002 13232 14058 13288
rect 14278 13776 14334 13832
rect 14554 14592 14610 14648
rect 14094 11192 14150 11248
rect 14002 9696 14058 9752
rect 15014 19488 15070 19544
rect 15382 20748 15384 20768
rect 15384 20748 15436 20768
rect 15436 20748 15438 20768
rect 15382 20712 15438 20748
rect 15658 20848 15714 20904
rect 15106 17992 15162 18048
rect 15290 18128 15346 18184
rect 15198 16088 15254 16144
rect 15106 15408 15162 15464
rect 15290 15680 15346 15736
rect 16670 26288 16726 26344
rect 15842 19488 15898 19544
rect 15750 18128 15806 18184
rect 15566 16224 15622 16280
rect 14830 13096 14886 13152
rect 14646 12280 14702 12336
rect 14554 12164 14610 12200
rect 14554 12144 14556 12164
rect 14556 12144 14608 12164
rect 14608 12144 14610 12164
rect 14646 11056 14702 11112
rect 15014 10784 15070 10840
rect 16026 17856 16082 17912
rect 17682 27920 17738 27976
rect 16210 18944 16266 19000
rect 16118 17448 16174 17504
rect 15934 15816 15990 15872
rect 16026 14612 16082 14648
rect 16026 14592 16028 14612
rect 16028 14592 16080 14612
rect 16080 14592 16082 14612
rect 16302 16360 16358 16416
rect 15842 11872 15898 11928
rect 16394 15408 16450 15464
rect 16670 17448 16726 17504
rect 15658 11636 15660 11656
rect 15660 11636 15712 11656
rect 15712 11636 15714 11656
rect 15658 11600 15714 11636
rect 15474 10376 15530 10432
rect 15014 10104 15070 10160
rect 14922 9832 14978 9888
rect 15198 9696 15254 9752
rect 12622 5616 12678 5672
rect 12070 4004 12126 4040
rect 12070 3984 12072 4004
rect 12072 3984 12124 4004
rect 12124 3984 12126 4004
rect 13266 4936 13322 4992
rect 13910 5344 13966 5400
rect 13818 4664 13874 4720
rect 13818 4256 13874 4312
rect 12254 3712 12310 3768
rect 12162 3576 12218 3632
rect 10414 1672 10470 1728
rect 12990 3884 12992 3904
rect 12992 3884 13044 3904
rect 13044 3884 13046 3904
rect 12990 3848 13046 3884
rect 13542 3984 13598 4040
rect 13634 3304 13690 3360
rect 13450 2624 13506 2680
rect 14922 9288 14978 9344
rect 14830 8744 14886 8800
rect 15474 8492 15530 8528
rect 15474 8472 15476 8492
rect 15476 8472 15528 8492
rect 15528 8472 15530 8492
rect 15106 8200 15162 8256
rect 14830 7656 14886 7712
rect 15290 6840 15346 6896
rect 15106 4256 15162 4312
rect 14830 3032 14886 3088
rect 15934 10784 15990 10840
rect 15842 9988 15898 10024
rect 15842 9968 15844 9988
rect 15844 9968 15896 9988
rect 15896 9968 15898 9988
rect 15750 8744 15806 8800
rect 16394 10240 16450 10296
rect 16302 9580 16358 9616
rect 16302 9560 16304 9580
rect 16304 9560 16356 9580
rect 16356 9560 16358 9580
rect 15658 6704 15714 6760
rect 15842 6704 15898 6760
rect 15658 6296 15714 6352
rect 15290 3848 15346 3904
rect 15658 6024 15714 6080
rect 14186 2760 14242 2816
rect 15474 2760 15530 2816
rect 15750 5072 15806 5128
rect 15842 4664 15898 4720
rect 16026 4256 16082 4312
rect 17038 18400 17094 18456
rect 16578 12280 16634 12336
rect 16578 9968 16634 10024
rect 16670 7812 16726 7848
rect 16670 7792 16672 7812
rect 16672 7792 16724 7812
rect 16724 7792 16726 7812
rect 16486 6160 16542 6216
rect 17682 22480 17738 22536
rect 17130 13640 17186 13696
rect 17314 17620 17316 17640
rect 17316 17620 17368 17640
rect 17368 17620 17370 17640
rect 17314 17584 17370 17620
rect 17314 17176 17370 17232
rect 17314 12860 17316 12880
rect 17316 12860 17368 12880
rect 17368 12860 17370 12880
rect 17314 12824 17370 12860
rect 17222 12688 17278 12744
rect 17038 11464 17094 11520
rect 16946 10920 17002 10976
rect 17498 16632 17554 16688
rect 17682 17312 17738 17368
rect 18326 22208 18382 22264
rect 18142 22072 18198 22128
rect 18050 20984 18106 21040
rect 17958 20304 18014 20360
rect 18326 21664 18382 21720
rect 18234 19624 18290 19680
rect 18142 19216 18198 19272
rect 18142 18708 18144 18728
rect 18144 18708 18196 18728
rect 18196 18708 18198 18728
rect 18142 18672 18198 18708
rect 17682 15272 17738 15328
rect 17590 14728 17646 14784
rect 17866 14728 17922 14784
rect 17682 13776 17738 13832
rect 17590 12688 17646 12744
rect 16854 6432 16910 6488
rect 16578 3712 16634 3768
rect 16394 3576 16450 3632
rect 16302 3304 16358 3360
rect 16762 3304 16818 3360
rect 16670 3168 16726 3224
rect 17038 9016 17094 9072
rect 17130 8472 17186 8528
rect 17222 8336 17278 8392
rect 17682 9016 17738 9072
rect 17958 12960 18014 13016
rect 17222 3712 17278 3768
rect 17406 5616 17462 5672
rect 17590 5072 17646 5128
rect 17314 3304 17370 3360
rect 17774 6860 17830 6896
rect 17774 6840 17776 6860
rect 17776 6840 17828 6860
rect 17828 6840 17830 6860
rect 17866 5616 17922 5672
rect 17866 5480 17922 5536
rect 18602 19216 18658 19272
rect 18602 16768 18658 16824
rect 18234 11328 18290 11384
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 18970 16904 19026 16960
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19246 19216 19302 19272
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19890 17604 19946 17640
rect 19890 17584 19892 17604
rect 19892 17584 19944 17604
rect 19944 17584 19946 17604
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19338 17040 19394 17096
rect 18970 14184 19026 14240
rect 18786 13640 18842 13696
rect 18970 13640 19026 13696
rect 18602 12824 18658 12880
rect 18602 10784 18658 10840
rect 18510 10376 18566 10432
rect 18418 10240 18474 10296
rect 18418 9832 18474 9888
rect 18234 7928 18290 7984
rect 18050 6840 18106 6896
rect 18050 6568 18106 6624
rect 18050 6452 18106 6488
rect 18050 6432 18052 6452
rect 18052 6432 18104 6452
rect 18104 6432 18106 6452
rect 18050 5752 18106 5808
rect 18142 5344 18198 5400
rect 18050 5072 18106 5128
rect 18786 10376 18842 10432
rect 19154 13504 19210 13560
rect 19246 12960 19302 13016
rect 19246 11464 19302 11520
rect 19706 17040 19762 17096
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 20258 16496 20314 16552
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19522 13776 19578 13832
rect 19890 13504 19946 13560
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19430 12280 19486 12336
rect 20074 12552 20130 12608
rect 19982 12144 20038 12200
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19430 11192 19486 11248
rect 19062 9016 19118 9072
rect 18694 5752 18750 5808
rect 17774 3460 17830 3496
rect 17774 3440 17776 3460
rect 17776 3440 17828 3460
rect 17828 3440 17830 3460
rect 18050 3304 18106 3360
rect 17958 3032 18014 3088
rect 18142 3032 18198 3088
rect 18878 7112 18934 7168
rect 18694 4256 18750 4312
rect 18878 3440 18934 3496
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 20258 15544 20314 15600
rect 20258 13640 20314 13696
rect 20258 11328 20314 11384
rect 20258 10648 20314 10704
rect 20166 10376 20222 10432
rect 20442 15544 20498 15600
rect 20442 12552 20498 12608
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19246 8064 19302 8120
rect 19154 7656 19210 7712
rect 19246 7520 19302 7576
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 20166 9324 20168 9344
rect 20168 9324 20220 9344
rect 20220 9324 20222 9344
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 20166 9288 20222 9324
rect 19338 5480 19394 5536
rect 19246 4392 19302 4448
rect 18970 3032 19026 3088
rect 20074 5480 20130 5536
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19982 5364 20038 5400
rect 20626 11192 20682 11248
rect 21178 17584 21234 17640
rect 20810 9696 20866 9752
rect 20718 6296 20774 6352
rect 20534 5480 20590 5536
rect 19982 5344 19984 5364
rect 19984 5344 20036 5364
rect 20036 5344 20038 5364
rect 20258 5344 20314 5400
rect 19338 4256 19394 4312
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19982 4256 20038 4312
rect 20626 5344 20682 5400
rect 20534 4800 20590 4856
rect 21178 6976 21234 7032
rect 20902 5616 20958 5672
rect 20718 4664 20774 4720
rect 19338 3712 19394 3768
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19246 3168 19302 3224
rect 20074 2896 20130 2952
rect 22374 15408 22430 15464
rect 21454 7384 21510 7440
rect 21362 6840 21418 6896
rect 22098 13368 22154 13424
rect 21730 11500 21732 11520
rect 21732 11500 21784 11520
rect 21784 11500 21786 11520
rect 21730 11464 21786 11500
rect 22006 11600 22062 11656
rect 21914 11328 21970 11384
rect 22006 11056 22062 11112
rect 21178 5344 21234 5400
rect 21086 5228 21142 5264
rect 21086 5208 21088 5228
rect 21088 5208 21140 5228
rect 21140 5208 21142 5228
rect 21178 3712 21234 3768
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 21730 8200 21786 8256
rect 21822 5752 21878 5808
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 23294 15000 23350 15056
rect 23294 11736 23350 11792
rect 23018 11600 23074 11656
rect 22466 8064 22522 8120
rect 22006 4936 22062 4992
rect 21914 4256 21970 4312
rect 21546 4020 21548 4040
rect 21548 4020 21600 4040
rect 21600 4020 21602 4040
rect 21546 3984 21602 4020
rect 22742 10532 22798 10568
rect 22742 10512 22744 10532
rect 22744 10512 22796 10532
rect 22796 10512 22798 10532
rect 22650 9424 22706 9480
rect 22742 8916 22744 8936
rect 22744 8916 22796 8936
rect 22796 8916 22798 8936
rect 22742 8880 22798 8916
rect 22650 8064 22706 8120
rect 23478 13504 23534 13560
rect 23386 10920 23442 10976
rect 24674 13912 24730 13968
rect 23570 10104 23626 10160
rect 23386 8492 23442 8528
rect 23386 8472 23388 8492
rect 23388 8472 23440 8492
rect 23440 8472 23442 8492
rect 23294 6740 23296 6760
rect 23296 6740 23348 6760
rect 23348 6740 23350 6760
rect 23294 6704 23350 6740
rect 22834 6024 22890 6080
rect 23294 5888 23350 5944
rect 22742 3440 22798 3496
rect 22558 3032 22614 3088
rect 23846 9968 23902 10024
rect 23754 5072 23810 5128
rect 23386 3884 23388 3904
rect 23388 3884 23440 3904
rect 23440 3884 23442 3904
rect 23386 3848 23442 3884
rect 23386 3612 23388 3632
rect 23388 3612 23440 3632
rect 23440 3612 23442 3632
rect 23386 3576 23442 3612
rect 22098 1672 22154 1728
rect 23386 2524 23388 2544
rect 23388 2524 23440 2544
rect 23440 2524 23442 2544
rect 23386 2488 23442 2524
rect 24030 2760 24086 2816
rect 27066 13232 27122 13288
rect 37186 38800 37242 38856
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 25134 11056 25190 11112
rect 24582 8336 24638 8392
rect 25318 7792 25374 7848
rect 24674 4528 24730 4584
rect 24582 4120 24638 4176
rect 26238 7948 26294 7984
rect 26238 7928 26240 7948
rect 26240 7928 26292 7948
rect 26292 7928 26294 7948
rect 23570 1808 23626 1864
rect 30654 6180 30710 6216
rect 30654 6160 30656 6180
rect 30656 6160 30708 6180
rect 30708 6160 30710 6180
rect 27158 2352 27214 2408
rect 26054 1944 26110 2000
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 38106 37440 38162 37496
rect 38198 36080 38254 36136
rect 37462 30676 37464 30696
rect 37464 30676 37516 30696
rect 37516 30676 37518 30696
rect 37462 30640 37518 30676
rect 37462 27956 37464 27976
rect 37464 27956 37516 27976
rect 37516 27956 37518 27976
rect 37462 27920 37518 27956
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 37186 10920 37242 10976
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 37462 7520 37518 7576
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 38106 35400 38162 35456
rect 38198 34040 38254 34096
rect 38106 32680 38162 32736
rect 38106 32000 38162 32056
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 38198 29280 38254 29336
rect 38198 27276 38200 27296
rect 38200 27276 38252 27296
rect 38252 27276 38254 27296
rect 38198 27240 38254 27276
rect 38290 25880 38346 25936
rect 38198 24556 38200 24576
rect 38200 24556 38252 24576
rect 38252 24556 38254 24576
rect 38198 24520 38254 24556
rect 38198 23840 38254 23896
rect 38198 22500 38254 22536
rect 38198 22480 38200 22500
rect 38200 22480 38252 22500
rect 38252 22480 38254 22500
rect 38198 21120 38254 21176
rect 38198 20440 38254 20496
rect 38290 19080 38346 19136
rect 38290 17720 38346 17776
rect 38198 16396 38200 16416
rect 38200 16396 38252 16416
rect 38252 16396 38254 16416
rect 38198 16360 38254 16396
rect 38290 15680 38346 15736
rect 38198 14320 38254 14376
rect 38198 12960 38254 13016
rect 38198 12688 38254 12744
rect 38106 12280 38162 12336
rect 38198 9560 38254 9616
rect 38106 8200 38162 8256
rect 38290 6160 38346 6216
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 36910 1400 36966 1456
rect 1674 720 1730 776
rect 38198 4800 38254 4856
rect 38290 4140 38346 4176
rect 38290 4120 38292 4140
rect 38292 4120 38344 4140
rect 38344 4120 38346 4140
rect 38290 2760 38346 2816
rect 37646 720 37702 776
<< metal3 >>
rect 200 38858 800 38888
rect 1761 38858 1827 38861
rect 200 38856 1827 38858
rect 200 38800 1766 38856
rect 1822 38800 1827 38856
rect 200 38798 1827 38800
rect 200 38768 800 38798
rect 1761 38795 1827 38798
rect 37181 38858 37247 38861
rect 39200 38858 39800 38888
rect 37181 38856 39800 38858
rect 37181 38800 37186 38856
rect 37242 38800 39800 38856
rect 37181 38798 39800 38800
rect 37181 38795 37247 38798
rect 39200 38768 39800 38798
rect 200 38178 800 38208
rect 1669 38178 1735 38181
rect 200 38176 1735 38178
rect 200 38120 1674 38176
rect 1730 38120 1735 38176
rect 200 38118 1735 38120
rect 200 38088 800 38118
rect 1669 38115 1735 38118
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 38101 37498 38167 37501
rect 39200 37498 39800 37528
rect 38101 37496 39800 37498
rect 38101 37440 38106 37496
rect 38162 37440 39800 37496
rect 38101 37438 39800 37440
rect 38101 37435 38167 37438
rect 39200 37408 39800 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 200 36818 800 36848
rect 2497 36818 2563 36821
rect 200 36816 2563 36818
rect 200 36760 2502 36816
rect 2558 36760 2563 36816
rect 200 36758 2563 36760
rect 200 36728 800 36758
rect 2497 36755 2563 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 38193 36138 38259 36141
rect 39200 36138 39800 36168
rect 38193 36136 39800 36138
rect 38193 36080 38198 36136
rect 38254 36080 39800 36136
rect 38193 36078 39800 36080
rect 38193 36075 38259 36078
rect 39200 36048 39800 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 200 35458 800 35488
rect 1577 35458 1643 35461
rect 200 35456 1643 35458
rect 200 35400 1582 35456
rect 1638 35400 1643 35456
rect 200 35398 1643 35400
rect 200 35368 800 35398
rect 1577 35395 1643 35398
rect 38101 35458 38167 35461
rect 39200 35458 39800 35488
rect 38101 35456 39800 35458
rect 38101 35400 38106 35456
rect 38162 35400 39800 35456
rect 38101 35398 39800 35400
rect 38101 35395 38167 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 39200 35368 39800 35398
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 200 34778 800 34808
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 1761 34778 1827 34781
rect 200 34776 1827 34778
rect 200 34720 1766 34776
rect 1822 34720 1827 34776
rect 200 34718 1827 34720
rect 200 34688 800 34718
rect 1761 34715 1827 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 38193 34098 38259 34101
rect 39200 34098 39800 34128
rect 38193 34096 39800 34098
rect 38193 34040 38198 34096
rect 38254 34040 39800 34096
rect 38193 34038 39800 34040
rect 38193 34035 38259 34038
rect 39200 34008 39800 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 200 33418 800 33448
rect 1761 33418 1827 33421
rect 200 33416 1827 33418
rect 200 33360 1766 33416
rect 1822 33360 1827 33416
rect 200 33358 1827 33360
rect 200 33328 800 33358
rect 1761 33355 1827 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 38101 32738 38167 32741
rect 39200 32738 39800 32768
rect 38101 32736 39800 32738
rect 38101 32680 38106 32736
rect 38162 32680 39800 32736
rect 38101 32678 39800 32680
rect 38101 32675 38167 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 39200 32648 39800 32678
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 200 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1761 32058 1827 32061
rect 200 32056 1827 32058
rect 200 32000 1766 32056
rect 1822 32000 1827 32056
rect 200 31998 1827 32000
rect 200 31968 800 31998
rect 1761 31995 1827 31998
rect 38101 32058 38167 32061
rect 39200 32058 39800 32088
rect 38101 32056 39800 32058
rect 38101 32000 38106 32056
rect 38162 32000 39800 32056
rect 38101 31998 39800 32000
rect 38101 31995 38167 31998
rect 39200 31968 39800 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 200 31378 800 31408
rect 1577 31378 1643 31381
rect 200 31376 1643 31378
rect 200 31320 1582 31376
rect 1638 31320 1643 31376
rect 200 31318 1643 31320
rect 200 31288 800 31318
rect 1577 31315 1643 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 37457 30698 37523 30701
rect 39200 30698 39800 30728
rect 37457 30696 39800 30698
rect 37457 30640 37462 30696
rect 37518 30640 39800 30696
rect 37457 30638 39800 30640
rect 37457 30635 37523 30638
rect 39200 30608 39800 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 200 30018 800 30048
rect 1761 30018 1827 30021
rect 200 30016 1827 30018
rect 200 29960 1766 30016
rect 1822 29960 1827 30016
rect 200 29958 1827 29960
rect 200 29928 800 29958
rect 1761 29955 1827 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 38193 29338 38259 29341
rect 39200 29338 39800 29368
rect 38193 29336 39800 29338
rect 38193 29280 38198 29336
rect 38254 29280 39800 29336
rect 38193 29278 39800 29280
rect 38193 29275 38259 29278
rect 39200 29248 39800 29278
rect 1577 29066 1643 29069
rect 1894 29066 1900 29068
rect 1577 29064 1900 29066
rect 1577 29008 1582 29064
rect 1638 29008 1900 29064
rect 1577 29006 1900 29008
rect 1577 29003 1643 29006
rect 1894 29004 1900 29006
rect 1964 29004 1970 29068
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 200 28658 800 28688
rect 1761 28658 1827 28661
rect 200 28656 1827 28658
rect 200 28600 1766 28656
rect 1822 28600 1827 28656
rect 200 28598 1827 28600
rect 200 28568 800 28598
rect 1761 28595 1827 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 2589 28114 2655 28117
rect 12566 28114 12572 28116
rect 2589 28112 12572 28114
rect 2589 28056 2594 28112
rect 2650 28056 12572 28112
rect 2589 28054 12572 28056
rect 2589 28051 2655 28054
rect 12566 28052 12572 28054
rect 12636 28052 12642 28116
rect 13118 27916 13124 27980
rect 13188 27978 13194 27980
rect 17677 27978 17743 27981
rect 13188 27976 17743 27978
rect 13188 27920 17682 27976
rect 17738 27920 17743 27976
rect 13188 27918 17743 27920
rect 13188 27916 13194 27918
rect 17677 27915 17743 27918
rect 37457 27978 37523 27981
rect 39200 27978 39800 28008
rect 37457 27976 39800 27978
rect 37457 27920 37462 27976
rect 37518 27920 39800 27976
rect 37457 27918 39800 27920
rect 37457 27915 37523 27918
rect 39200 27888 39800 27918
rect 974 27780 980 27844
rect 1044 27842 1050 27844
rect 3233 27842 3299 27845
rect 1044 27840 3299 27842
rect 1044 27784 3238 27840
rect 3294 27784 3299 27840
rect 1044 27782 3299 27784
rect 1044 27780 1050 27782
rect 3233 27779 3299 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 1710 27644 1716 27708
rect 1780 27706 1786 27708
rect 1853 27706 1919 27709
rect 1780 27704 1919 27706
rect 1780 27648 1858 27704
rect 1914 27648 1919 27704
rect 1780 27646 1919 27648
rect 1780 27644 1786 27646
rect 1853 27643 1919 27646
rect 2037 27708 2103 27709
rect 2037 27704 2084 27708
rect 2148 27706 2154 27708
rect 2037 27648 2042 27704
rect 2037 27644 2084 27648
rect 2148 27646 2194 27706
rect 2148 27644 2154 27646
rect 2037 27643 2103 27644
rect 200 27298 800 27328
rect 4061 27298 4127 27301
rect 200 27296 4127 27298
rect 200 27240 4066 27296
rect 4122 27240 4127 27296
rect 200 27238 4127 27240
rect 200 27208 800 27238
rect 4061 27235 4127 27238
rect 38193 27298 38259 27301
rect 39200 27298 39800 27328
rect 38193 27296 39800 27298
rect 38193 27240 38198 27296
rect 38254 27240 39800 27296
rect 38193 27238 39800 27240
rect 38193 27235 38259 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 39200 27208 39800 27238
rect 19570 27167 19886 27168
rect 2497 26890 2563 26893
rect 5574 26890 5580 26892
rect 2497 26888 5580 26890
rect 2497 26832 2502 26888
rect 2558 26832 5580 26888
rect 2497 26830 5580 26832
rect 2497 26827 2563 26830
rect 5574 26828 5580 26830
rect 5644 26828 5650 26892
rect 1945 26754 2011 26757
rect 2998 26754 3004 26756
rect 1945 26752 3004 26754
rect 1945 26696 1950 26752
rect 2006 26696 3004 26752
rect 1945 26694 3004 26696
rect 1945 26691 2011 26694
rect 2998 26692 3004 26694
rect 3068 26692 3074 26756
rect 4210 26688 4526 26689
rect 200 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 3417 26618 3483 26621
rect 200 26616 3483 26618
rect 200 26560 3422 26616
rect 3478 26560 3483 26616
rect 200 26558 3483 26560
rect 200 26528 800 26558
rect 3417 26555 3483 26558
rect 1853 26482 1919 26485
rect 5758 26482 5764 26484
rect 1853 26480 5764 26482
rect 1853 26424 1858 26480
rect 1914 26424 5764 26480
rect 1853 26422 5764 26424
rect 1853 26419 1919 26422
rect 5758 26420 5764 26422
rect 5828 26420 5834 26484
rect 1158 26284 1164 26348
rect 1228 26346 1234 26348
rect 2497 26346 2563 26349
rect 1228 26344 2563 26346
rect 1228 26288 2502 26344
rect 2558 26288 2563 26344
rect 1228 26286 2563 26288
rect 1228 26284 1234 26286
rect 2497 26283 2563 26286
rect 4613 26348 4679 26349
rect 4613 26344 4660 26348
rect 4724 26346 4730 26348
rect 4613 26288 4618 26344
rect 4613 26284 4660 26288
rect 4724 26286 4770 26346
rect 4724 26284 4730 26286
rect 10542 26284 10548 26348
rect 10612 26346 10618 26348
rect 14365 26346 14431 26349
rect 16665 26346 16731 26349
rect 10612 26344 16731 26346
rect 10612 26288 14370 26344
rect 14426 26288 16670 26344
rect 16726 26288 16731 26344
rect 10612 26286 16731 26288
rect 10612 26284 10618 26286
rect 4613 26283 4679 26284
rect 14365 26283 14431 26286
rect 16665 26283 16731 26286
rect 2773 26212 2839 26213
rect 2773 26208 2820 26212
rect 2884 26210 2890 26212
rect 11421 26210 11487 26213
rect 16614 26210 16620 26212
rect 2773 26152 2778 26208
rect 2773 26148 2820 26152
rect 2884 26150 2930 26210
rect 11421 26208 16620 26210
rect 11421 26152 11426 26208
rect 11482 26152 16620 26208
rect 11421 26150 16620 26152
rect 2884 26148 2890 26150
rect 2773 26147 2839 26148
rect 11421 26147 11487 26150
rect 16614 26148 16620 26150
rect 16684 26148 16690 26212
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 38285 25938 38351 25941
rect 39200 25938 39800 25968
rect 38285 25936 39800 25938
rect 38285 25880 38290 25936
rect 38346 25880 39800 25936
rect 38285 25878 39800 25880
rect 38285 25875 38351 25878
rect 39200 25848 39800 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 200 25258 800 25288
rect 1761 25258 1827 25261
rect 200 25256 1827 25258
rect 200 25200 1766 25256
rect 1822 25200 1827 25256
rect 200 25198 1827 25200
rect 200 25168 800 25198
rect 1761 25195 1827 25198
rect 2221 25258 2287 25261
rect 9254 25258 9260 25260
rect 2221 25256 9260 25258
rect 2221 25200 2226 25256
rect 2282 25200 9260 25256
rect 2221 25198 9260 25200
rect 2221 25195 2287 25198
rect 9254 25196 9260 25198
rect 9324 25196 9330 25260
rect 7189 25124 7255 25125
rect 7189 25120 7236 25124
rect 7300 25122 7306 25124
rect 7189 25064 7194 25120
rect 7189 25060 7236 25064
rect 7300 25062 7346 25122
rect 7300 25060 7306 25062
rect 7189 25059 7255 25060
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 790 24924 796 24988
rect 860 24986 866 24988
rect 1393 24986 1459 24989
rect 860 24984 1459 24986
rect 860 24928 1398 24984
rect 1454 24928 1459 24984
rect 860 24926 1459 24928
rect 860 24924 866 24926
rect 1393 24923 1459 24926
rect 3877 24988 3943 24989
rect 3877 24984 3924 24988
rect 3988 24986 3994 24988
rect 3877 24928 3882 24984
rect 3877 24924 3924 24928
rect 3988 24926 4034 24986
rect 3988 24924 3994 24926
rect 4838 24924 4844 24988
rect 4908 24986 4914 24988
rect 5165 24986 5231 24989
rect 4908 24984 5231 24986
rect 4908 24928 5170 24984
rect 5226 24928 5231 24984
rect 4908 24926 5231 24928
rect 4908 24924 4914 24926
rect 3877 24923 3943 24924
rect 5165 24923 5231 24926
rect 7005 24988 7071 24989
rect 7005 24984 7052 24988
rect 7116 24986 7122 24988
rect 9673 24986 9739 24989
rect 15510 24986 15516 24988
rect 7005 24928 7010 24984
rect 7005 24924 7052 24928
rect 7116 24926 7162 24986
rect 9673 24984 15516 24986
rect 9673 24928 9678 24984
rect 9734 24928 15516 24984
rect 9673 24926 15516 24928
rect 7116 24924 7122 24926
rect 7005 24923 7071 24924
rect 9673 24923 9739 24926
rect 15510 24924 15516 24926
rect 15580 24924 15586 24988
rect 4797 24850 4863 24853
rect 5165 24850 5231 24853
rect 4797 24848 5231 24850
rect 4797 24792 4802 24848
rect 4858 24792 5170 24848
rect 5226 24792 5231 24848
rect 4797 24790 5231 24792
rect 4797 24787 4863 24790
rect 5165 24787 5231 24790
rect 5942 24788 5948 24852
rect 6012 24850 6018 24852
rect 6545 24850 6611 24853
rect 6012 24848 6611 24850
rect 6012 24792 6550 24848
rect 6606 24792 6611 24848
rect 6012 24790 6611 24792
rect 6012 24788 6018 24790
rect 6545 24787 6611 24790
rect 8886 24788 8892 24852
rect 8956 24850 8962 24852
rect 9121 24850 9187 24853
rect 8956 24848 9187 24850
rect 8956 24792 9126 24848
rect 9182 24792 9187 24848
rect 8956 24790 9187 24792
rect 8956 24788 8962 24790
rect 9121 24787 9187 24790
rect 38193 24578 38259 24581
rect 39200 24578 39800 24608
rect 38193 24576 39800 24578
rect 38193 24520 38198 24576
rect 38254 24520 39800 24576
rect 38193 24518 39800 24520
rect 38193 24515 38259 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 39200 24488 39800 24518
rect 34930 24447 35246 24448
rect 3550 24108 3556 24172
rect 3620 24170 3626 24172
rect 3969 24170 4035 24173
rect 4797 24170 4863 24173
rect 3620 24168 4863 24170
rect 3620 24112 3974 24168
rect 4030 24112 4802 24168
rect 4858 24112 4863 24168
rect 3620 24110 4863 24112
rect 3620 24108 3626 24110
rect 3969 24107 4035 24110
rect 4797 24107 4863 24110
rect 2497 24034 2563 24037
rect 2630 24034 2636 24036
rect 2497 24032 2636 24034
rect 2497 23976 2502 24032
rect 2558 23976 2636 24032
rect 2497 23974 2636 23976
rect 2497 23971 2563 23974
rect 2630 23972 2636 23974
rect 2700 23972 2706 24036
rect 19570 23968 19886 23969
rect 200 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 1761 23898 1827 23901
rect 200 23896 1827 23898
rect 200 23840 1766 23896
rect 1822 23840 1827 23896
rect 200 23838 1827 23840
rect 200 23808 800 23838
rect 1761 23835 1827 23838
rect 3877 23898 3943 23901
rect 7649 23898 7715 23901
rect 3877 23896 7715 23898
rect 3877 23840 3882 23896
rect 3938 23840 7654 23896
rect 7710 23840 7715 23896
rect 3877 23838 7715 23840
rect 3877 23835 3943 23838
rect 7649 23835 7715 23838
rect 38193 23898 38259 23901
rect 39200 23898 39800 23928
rect 38193 23896 39800 23898
rect 38193 23840 38198 23896
rect 38254 23840 39800 23896
rect 38193 23838 39800 23840
rect 38193 23835 38259 23838
rect 39200 23808 39800 23838
rect 4705 23626 4771 23629
rect 8385 23626 8451 23629
rect 10910 23626 10916 23628
rect 4705 23624 8172 23626
rect 4705 23568 4710 23624
rect 4766 23568 8172 23624
rect 4705 23566 8172 23568
rect 4705 23563 4771 23566
rect 3182 23428 3188 23492
rect 3252 23490 3258 23492
rect 3417 23490 3483 23493
rect 3252 23488 3483 23490
rect 3252 23432 3422 23488
rect 3478 23432 3483 23488
rect 3252 23430 3483 23432
rect 3252 23428 3258 23430
rect 3417 23427 3483 23430
rect 3601 23490 3667 23493
rect 3734 23490 3740 23492
rect 3601 23488 3740 23490
rect 3601 23432 3606 23488
rect 3662 23432 3740 23488
rect 3601 23430 3740 23432
rect 3601 23427 3667 23430
rect 3734 23428 3740 23430
rect 3804 23428 3810 23492
rect 7465 23490 7531 23493
rect 7598 23490 7604 23492
rect 7465 23488 7604 23490
rect 7465 23432 7470 23488
rect 7526 23432 7604 23488
rect 7465 23430 7604 23432
rect 7465 23427 7531 23430
rect 7598 23428 7604 23430
rect 7668 23428 7674 23492
rect 8112 23490 8172 23566
rect 8385 23624 10916 23626
rect 8385 23568 8390 23624
rect 8446 23568 10916 23624
rect 8385 23566 10916 23568
rect 8385 23563 8451 23566
rect 10910 23564 10916 23566
rect 10980 23564 10986 23628
rect 11697 23626 11763 23629
rect 11830 23626 11836 23628
rect 11697 23624 11836 23626
rect 11697 23568 11702 23624
rect 11758 23568 11836 23624
rect 11697 23566 11836 23568
rect 11697 23563 11763 23566
rect 11830 23564 11836 23566
rect 11900 23564 11906 23628
rect 10225 23492 10291 23493
rect 9990 23490 9996 23492
rect 8112 23430 9996 23490
rect 9990 23428 9996 23430
rect 10060 23428 10066 23492
rect 10174 23490 10180 23492
rect 10134 23430 10180 23490
rect 10244 23488 10291 23492
rect 10286 23432 10291 23488
rect 10174 23428 10180 23430
rect 10244 23428 10291 23432
rect 10225 23427 10291 23428
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 200 23218 800 23248
rect 1669 23218 1735 23221
rect 200 23216 1735 23218
rect 200 23160 1674 23216
rect 1730 23160 1735 23216
rect 200 23158 1735 23160
rect 200 23128 800 23158
rect 1669 23155 1735 23158
rect 7741 23082 7807 23085
rect 14406 23082 14412 23084
rect 7741 23080 14412 23082
rect 7741 23024 7746 23080
rect 7802 23024 14412 23080
rect 7741 23022 14412 23024
rect 7741 23019 7807 23022
rect 14406 23020 14412 23022
rect 14476 23020 14482 23084
rect 12157 22946 12223 22949
rect 12709 22946 12775 22949
rect 12157 22944 12775 22946
rect 12157 22888 12162 22944
rect 12218 22888 12714 22944
rect 12770 22888 12775 22944
rect 12157 22886 12775 22888
rect 12157 22883 12223 22886
rect 12709 22883 12775 22886
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 2681 22538 2747 22541
rect 5257 22538 5323 22541
rect 2681 22536 5323 22538
rect 2681 22480 2686 22536
rect 2742 22480 5262 22536
rect 5318 22480 5323 22536
rect 2681 22478 5323 22480
rect 2681 22475 2747 22478
rect 5257 22475 5323 22478
rect 17677 22538 17743 22541
rect 20110 22538 20116 22540
rect 17677 22536 20116 22538
rect 17677 22480 17682 22536
rect 17738 22480 20116 22536
rect 17677 22478 20116 22480
rect 17677 22475 17743 22478
rect 20110 22476 20116 22478
rect 20180 22476 20186 22540
rect 38193 22538 38259 22541
rect 39200 22538 39800 22568
rect 38193 22536 39800 22538
rect 38193 22480 38198 22536
rect 38254 22480 39800 22536
rect 38193 22478 39800 22480
rect 38193 22475 38259 22478
rect 39200 22448 39800 22478
rect 6494 22340 6500 22404
rect 6564 22402 6570 22404
rect 6729 22402 6795 22405
rect 6564 22400 6795 22402
rect 6564 22344 6734 22400
rect 6790 22344 6795 22400
rect 6564 22342 6795 22344
rect 6564 22340 6570 22342
rect 6729 22339 6795 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 11094 22204 11100 22268
rect 11164 22266 11170 22268
rect 18321 22266 18387 22269
rect 11164 22264 18387 22266
rect 11164 22208 18326 22264
rect 18382 22208 18387 22264
rect 11164 22206 18387 22208
rect 11164 22204 11170 22206
rect 18321 22203 18387 22206
rect 9673 22130 9739 22133
rect 11881 22130 11947 22133
rect 12617 22130 12683 22133
rect 18137 22130 18203 22133
rect 9673 22128 18203 22130
rect 9673 22072 9678 22128
rect 9734 22072 11886 22128
rect 11942 22072 12622 22128
rect 12678 22072 18142 22128
rect 18198 22072 18203 22128
rect 9673 22070 18203 22072
rect 9673 22067 9739 22070
rect 11881 22067 11947 22070
rect 12617 22067 12683 22070
rect 18137 22067 18203 22070
rect 3734 21932 3740 21996
rect 3804 21994 3810 21996
rect 4981 21994 5047 21997
rect 3804 21992 5047 21994
rect 3804 21936 4986 21992
rect 5042 21936 5047 21992
rect 3804 21934 5047 21936
rect 3804 21932 3810 21934
rect 4981 21931 5047 21934
rect 6361 21994 6427 21997
rect 6862 21994 6868 21996
rect 6361 21992 6868 21994
rect 6361 21936 6366 21992
rect 6422 21936 6868 21992
rect 6361 21934 6868 21936
rect 6361 21931 6427 21934
rect 6862 21932 6868 21934
rect 6932 21932 6938 21996
rect 8109 21994 8175 21997
rect 12709 21994 12775 21997
rect 8109 21992 12775 21994
rect 8109 21936 8114 21992
rect 8170 21936 12714 21992
rect 12770 21936 12775 21992
rect 8109 21934 12775 21936
rect 8109 21931 8175 21934
rect 12709 21931 12775 21934
rect 200 21858 800 21888
rect 1761 21858 1827 21861
rect 5073 21860 5139 21861
rect 200 21856 1827 21858
rect 200 21800 1766 21856
rect 1822 21800 1827 21856
rect 200 21798 1827 21800
rect 200 21768 800 21798
rect 1761 21795 1827 21798
rect 5022 21796 5028 21860
rect 5092 21858 5139 21860
rect 11053 21858 11119 21861
rect 15009 21858 15075 21861
rect 5092 21856 5184 21858
rect 5134 21800 5184 21856
rect 5092 21798 5184 21800
rect 11053 21856 15075 21858
rect 11053 21800 11058 21856
rect 11114 21800 15014 21856
rect 15070 21800 15075 21856
rect 11053 21798 15075 21800
rect 5092 21796 5139 21798
rect 5073 21795 5139 21796
rect 11053 21795 11119 21798
rect 15009 21795 15075 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4337 21722 4403 21725
rect 9397 21722 9463 21725
rect 4337 21720 9463 21722
rect 4337 21664 4342 21720
rect 4398 21664 9402 21720
rect 9458 21664 9463 21720
rect 4337 21662 9463 21664
rect 4337 21659 4403 21662
rect 9397 21659 9463 21662
rect 12801 21722 12867 21725
rect 18321 21722 18387 21725
rect 12801 21720 18387 21722
rect 12801 21664 12806 21720
rect 12862 21664 18326 21720
rect 18382 21664 18387 21720
rect 12801 21662 18387 21664
rect 12801 21659 12867 21662
rect 18321 21659 18387 21662
rect 6361 21586 6427 21589
rect 10501 21586 10567 21589
rect 11094 21586 11100 21588
rect 6361 21584 11100 21586
rect 6361 21528 6366 21584
rect 6422 21528 10506 21584
rect 10562 21528 11100 21584
rect 6361 21526 11100 21528
rect 6361 21523 6427 21526
rect 10501 21523 10567 21526
rect 11094 21524 11100 21526
rect 11164 21524 11170 21588
rect 3918 21388 3924 21452
rect 3988 21450 3994 21452
rect 10961 21450 11027 21453
rect 3988 21448 11027 21450
rect 3988 21392 10966 21448
rect 11022 21392 11027 21448
rect 3988 21390 11027 21392
rect 3988 21388 3994 21390
rect 10961 21387 11027 21390
rect 10869 21314 10935 21317
rect 12249 21314 12315 21317
rect 10869 21312 12315 21314
rect 10869 21256 10874 21312
rect 10930 21256 12254 21312
rect 12310 21256 12315 21312
rect 10869 21254 12315 21256
rect 10869 21251 10935 21254
rect 12249 21251 12315 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 38193 21178 38259 21181
rect 39200 21178 39800 21208
rect 38193 21176 39800 21178
rect 38193 21120 38198 21176
rect 38254 21120 39800 21176
rect 38193 21118 39800 21120
rect 38193 21115 38259 21118
rect 39200 21088 39800 21118
rect 3550 20980 3556 21044
rect 3620 21042 3626 21044
rect 4153 21042 4219 21045
rect 3620 21040 4219 21042
rect 3620 20984 4158 21040
rect 4214 20984 4219 21040
rect 3620 20982 4219 20984
rect 3620 20980 3626 20982
rect 4153 20979 4219 20982
rect 9673 21042 9739 21045
rect 10961 21042 11027 21045
rect 9673 21040 11027 21042
rect 9673 20984 9678 21040
rect 9734 20984 10966 21040
rect 11022 20984 11027 21040
rect 9673 20982 11027 20984
rect 9673 20979 9739 20982
rect 10961 20979 11027 20982
rect 13537 21042 13603 21045
rect 18045 21042 18111 21045
rect 13537 21040 18111 21042
rect 13537 20984 13542 21040
rect 13598 20984 18050 21040
rect 18106 20984 18111 21040
rect 13537 20982 18111 20984
rect 13537 20979 13603 20982
rect 18045 20979 18111 20982
rect 8937 20906 9003 20909
rect 10133 20906 10199 20909
rect 8937 20904 10199 20906
rect 8937 20848 8942 20904
rect 8998 20848 10138 20904
rect 10194 20848 10199 20904
rect 8937 20846 10199 20848
rect 8937 20843 9003 20846
rect 10133 20843 10199 20846
rect 13353 20906 13419 20909
rect 15653 20906 15719 20909
rect 13353 20904 15719 20906
rect 13353 20848 13358 20904
rect 13414 20848 15658 20904
rect 15714 20848 15719 20904
rect 13353 20846 15719 20848
rect 13353 20843 13419 20846
rect 15653 20843 15719 20846
rect 4705 20772 4771 20773
rect 4654 20770 4660 20772
rect 4614 20710 4660 20770
rect 4724 20768 4771 20772
rect 4766 20712 4771 20768
rect 4654 20708 4660 20710
rect 4724 20708 4771 20712
rect 4705 20707 4771 20708
rect 14273 20770 14339 20773
rect 15377 20770 15443 20773
rect 14273 20768 15443 20770
rect 14273 20712 14278 20768
rect 14334 20712 15382 20768
rect 15438 20712 15443 20768
rect 14273 20710 15443 20712
rect 14273 20707 14339 20710
rect 15377 20707 15443 20710
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4797 20634 4863 20637
rect 9673 20634 9739 20637
rect 4797 20632 9739 20634
rect 4797 20576 4802 20632
rect 4858 20576 9678 20632
rect 9734 20576 9739 20632
rect 4797 20574 9739 20576
rect 4797 20571 4863 20574
rect 9673 20571 9739 20574
rect 200 20498 800 20528
rect 3693 20498 3759 20501
rect 200 20496 3759 20498
rect 200 20440 3698 20496
rect 3754 20440 3759 20496
rect 200 20438 3759 20440
rect 200 20408 800 20438
rect 3693 20435 3759 20438
rect 3969 20498 4035 20501
rect 6453 20498 6519 20501
rect 7557 20498 7623 20501
rect 3969 20496 6194 20498
rect 3969 20440 3974 20496
rect 4030 20440 6194 20496
rect 3969 20438 6194 20440
rect 3969 20435 4035 20438
rect 3325 20362 3391 20365
rect 5942 20362 5948 20364
rect 3325 20360 5948 20362
rect 3325 20304 3330 20360
rect 3386 20304 5948 20360
rect 3325 20302 5948 20304
rect 3325 20299 3391 20302
rect 5942 20300 5948 20302
rect 6012 20300 6018 20364
rect 6134 20362 6194 20438
rect 6453 20496 7623 20498
rect 6453 20440 6458 20496
rect 6514 20440 7562 20496
rect 7618 20440 7623 20496
rect 6453 20438 7623 20440
rect 6453 20435 6519 20438
rect 7557 20435 7623 20438
rect 9990 20436 9996 20500
rect 10060 20498 10066 20500
rect 10777 20498 10843 20501
rect 10060 20496 10843 20498
rect 10060 20440 10782 20496
rect 10838 20440 10843 20496
rect 10060 20438 10843 20440
rect 10060 20436 10066 20438
rect 10777 20435 10843 20438
rect 38193 20498 38259 20501
rect 39200 20498 39800 20528
rect 38193 20496 39800 20498
rect 38193 20440 38198 20496
rect 38254 20440 39800 20496
rect 38193 20438 39800 20440
rect 38193 20435 38259 20438
rect 39200 20408 39800 20438
rect 7925 20362 7991 20365
rect 17953 20362 18019 20365
rect 6134 20360 18019 20362
rect 6134 20304 7930 20360
rect 7986 20304 17958 20360
rect 18014 20304 18019 20360
rect 6134 20302 18019 20304
rect 7925 20299 7991 20302
rect 17953 20299 18019 20302
rect 4797 20226 4863 20229
rect 5073 20226 5139 20229
rect 4797 20224 5139 20226
rect 4797 20168 4802 20224
rect 4858 20168 5078 20224
rect 5134 20168 5139 20224
rect 4797 20166 5139 20168
rect 4797 20163 4863 20166
rect 5073 20163 5139 20166
rect 5901 20226 5967 20229
rect 6729 20226 6795 20229
rect 9305 20226 9371 20229
rect 5901 20224 9371 20226
rect 5901 20168 5906 20224
rect 5962 20168 6734 20224
rect 6790 20168 9310 20224
rect 9366 20168 9371 20224
rect 5901 20166 9371 20168
rect 5901 20163 5967 20166
rect 6729 20163 6795 20166
rect 9305 20163 9371 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 5349 20090 5415 20093
rect 8937 20090 9003 20093
rect 5349 20088 9003 20090
rect 5349 20032 5354 20088
rect 5410 20032 8942 20088
rect 8998 20032 9003 20088
rect 5349 20030 9003 20032
rect 5349 20027 5415 20030
rect 8937 20027 9003 20030
rect 4613 19954 4679 19957
rect 7465 19954 7531 19957
rect 4613 19952 7531 19954
rect 4613 19896 4618 19952
rect 4674 19896 7470 19952
rect 7526 19896 7531 19952
rect 4613 19894 7531 19896
rect 4613 19891 4679 19894
rect 7465 19891 7531 19894
rect 9121 19954 9187 19957
rect 11145 19954 11211 19957
rect 9121 19952 11211 19954
rect 9121 19896 9126 19952
rect 9182 19896 11150 19952
rect 11206 19896 11211 19952
rect 9121 19894 11211 19896
rect 9121 19891 9187 19894
rect 11145 19891 11211 19894
rect 6821 19818 6887 19821
rect 7741 19818 7807 19821
rect 6821 19816 7807 19818
rect 6821 19760 6826 19816
rect 6882 19760 7746 19816
rect 7802 19760 7807 19816
rect 6821 19758 7807 19760
rect 6821 19755 6887 19758
rect 7741 19755 7807 19758
rect 4889 19682 4955 19685
rect 5022 19682 5028 19684
rect 4889 19680 5028 19682
rect 4889 19624 4894 19680
rect 4950 19624 5028 19680
rect 4889 19622 5028 19624
rect 4889 19619 4955 19622
rect 5022 19620 5028 19622
rect 5092 19620 5098 19684
rect 5165 19682 5231 19685
rect 8753 19682 8819 19685
rect 5165 19680 8819 19682
rect 5165 19624 5170 19680
rect 5226 19624 8758 19680
rect 8814 19624 8819 19680
rect 5165 19622 8819 19624
rect 5165 19619 5231 19622
rect 8753 19619 8819 19622
rect 14365 19682 14431 19685
rect 18229 19682 18295 19685
rect 14365 19680 18295 19682
rect 14365 19624 14370 19680
rect 14426 19624 18234 19680
rect 18290 19624 18295 19680
rect 14365 19622 18295 19624
rect 14365 19619 14431 19622
rect 18229 19619 18295 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 5073 19546 5139 19549
rect 11094 19546 11100 19548
rect 5073 19544 11100 19546
rect 5073 19488 5078 19544
rect 5134 19488 11100 19544
rect 5073 19486 11100 19488
rect 5073 19483 5139 19486
rect 11094 19484 11100 19486
rect 11164 19484 11170 19548
rect 12985 19546 13051 19549
rect 15009 19546 15075 19549
rect 15837 19546 15903 19549
rect 12985 19544 15903 19546
rect 12985 19488 12990 19544
rect 13046 19488 15014 19544
rect 15070 19488 15842 19544
rect 15898 19488 15903 19544
rect 12985 19486 15903 19488
rect 12985 19483 13051 19486
rect 15009 19483 15075 19486
rect 15837 19483 15903 19486
rect 3693 19410 3759 19413
rect 6637 19412 6703 19413
rect 4838 19410 4844 19412
rect 3693 19408 4844 19410
rect 3693 19352 3698 19408
rect 3754 19352 4844 19408
rect 3693 19350 4844 19352
rect 3693 19347 3759 19350
rect 4838 19348 4844 19350
rect 4908 19348 4914 19412
rect 6637 19410 6684 19412
rect 6592 19408 6684 19410
rect 6592 19352 6642 19408
rect 6592 19350 6684 19352
rect 6637 19348 6684 19350
rect 6748 19348 6754 19412
rect 6913 19410 6979 19413
rect 8109 19410 8175 19413
rect 6913 19408 8175 19410
rect 6913 19352 6918 19408
rect 6974 19352 8114 19408
rect 8170 19352 8175 19408
rect 6913 19350 8175 19352
rect 6637 19347 6703 19348
rect 6913 19347 6979 19350
rect 8109 19347 8175 19350
rect 1853 19276 1919 19277
rect 2129 19276 2195 19277
rect 1853 19274 1900 19276
rect 1808 19272 1900 19274
rect 1808 19216 1858 19272
rect 1808 19214 1900 19216
rect 1853 19212 1900 19214
rect 1964 19212 1970 19276
rect 2078 19274 2084 19276
rect 2038 19214 2084 19274
rect 2148 19272 2195 19276
rect 2190 19216 2195 19272
rect 2078 19212 2084 19214
rect 2148 19212 2195 19216
rect 1853 19211 1919 19212
rect 2129 19211 2195 19212
rect 2865 19274 2931 19277
rect 2998 19274 3004 19276
rect 2865 19272 3004 19274
rect 2865 19216 2870 19272
rect 2926 19216 3004 19272
rect 2865 19214 3004 19216
rect 2865 19211 2931 19214
rect 2998 19212 3004 19214
rect 3068 19212 3074 19276
rect 4521 19274 4587 19277
rect 4654 19274 4660 19276
rect 4521 19272 4660 19274
rect 4521 19216 4526 19272
rect 4582 19216 4660 19272
rect 4521 19214 4660 19216
rect 4521 19211 4587 19214
rect 4654 19212 4660 19214
rect 4724 19212 4730 19276
rect 17718 19212 17724 19276
rect 17788 19274 17794 19276
rect 18137 19274 18203 19277
rect 17788 19272 18203 19274
rect 17788 19216 18142 19272
rect 18198 19216 18203 19272
rect 17788 19214 18203 19216
rect 17788 19212 17794 19214
rect 18137 19211 18203 19214
rect 18597 19274 18663 19277
rect 19241 19274 19307 19277
rect 18597 19272 19307 19274
rect 18597 19216 18602 19272
rect 18658 19216 19246 19272
rect 19302 19216 19307 19272
rect 18597 19214 19307 19216
rect 18597 19211 18663 19214
rect 19241 19211 19307 19214
rect 200 19138 800 19168
rect 2814 19138 2820 19140
rect 200 19078 2820 19138
rect 200 19048 800 19078
rect 2814 19076 2820 19078
rect 2884 19076 2890 19140
rect 10041 19138 10107 19141
rect 12341 19138 12407 19141
rect 10041 19136 12407 19138
rect 10041 19080 10046 19136
rect 10102 19080 12346 19136
rect 12402 19080 12407 19136
rect 10041 19078 12407 19080
rect 10041 19075 10107 19078
rect 12341 19075 12407 19078
rect 38285 19138 38351 19141
rect 39200 19138 39800 19168
rect 38285 19136 39800 19138
rect 38285 19080 38290 19136
rect 38346 19080 39800 19136
rect 38285 19078 39800 19080
rect 38285 19075 38351 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 39800 19078
rect 34930 19007 35246 19008
rect 1158 18940 1164 19004
rect 1228 19002 1234 19004
rect 2497 19002 2563 19005
rect 8569 19002 8635 19005
rect 1228 19000 2563 19002
rect 1228 18944 2502 19000
rect 2558 18944 2563 19000
rect 1228 18942 2563 18944
rect 1228 18940 1234 18942
rect 2497 18939 2563 18942
rect 8526 19000 8635 19002
rect 8526 18944 8574 19000
rect 8630 18944 8635 19000
rect 8526 18939 8635 18944
rect 11697 19002 11763 19005
rect 12341 19002 12407 19005
rect 14733 19002 14799 19005
rect 16205 19002 16271 19005
rect 11697 19000 16271 19002
rect 11697 18944 11702 19000
rect 11758 18944 12346 19000
rect 12402 18944 14738 19000
rect 14794 18944 16210 19000
rect 16266 18944 16271 19000
rect 11697 18942 16271 18944
rect 11697 18939 11763 18942
rect 12341 18939 12407 18942
rect 14733 18939 14799 18942
rect 16205 18939 16271 18942
rect 4245 18866 4311 18869
rect 8526 18866 8586 18939
rect 4245 18864 8586 18866
rect 4245 18808 4250 18864
rect 4306 18808 8586 18864
rect 4245 18806 8586 18808
rect 4245 18803 4311 18806
rect 6361 18730 6427 18733
rect 9305 18730 9371 18733
rect 6361 18728 9371 18730
rect 6361 18672 6366 18728
rect 6422 18672 9310 18728
rect 9366 18672 9371 18728
rect 6361 18670 9371 18672
rect 6361 18667 6427 18670
rect 9305 18667 9371 18670
rect 16430 18668 16436 18732
rect 16500 18730 16506 18732
rect 18137 18730 18203 18733
rect 16500 18728 18203 18730
rect 16500 18672 18142 18728
rect 18198 18672 18203 18728
rect 16500 18670 18203 18672
rect 16500 18668 16506 18670
rect 18137 18667 18203 18670
rect 12157 18594 12223 18597
rect 13629 18594 13695 18597
rect 12157 18592 13695 18594
rect 12157 18536 12162 18592
rect 12218 18536 13634 18592
rect 13690 18536 13695 18592
rect 12157 18534 13695 18536
rect 12157 18531 12223 18534
rect 13629 18531 13695 18534
rect 19570 18528 19886 18529
rect 200 18458 800 18488
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 3049 18458 3115 18461
rect 200 18456 3115 18458
rect 200 18400 3054 18456
rect 3110 18400 3115 18456
rect 200 18398 3115 18400
rect 200 18368 800 18398
rect 3049 18395 3115 18398
rect 10041 18458 10107 18461
rect 10869 18458 10935 18461
rect 10041 18456 10935 18458
rect 10041 18400 10046 18456
rect 10102 18400 10874 18456
rect 10930 18400 10935 18456
rect 10041 18398 10935 18400
rect 10041 18395 10107 18398
rect 10869 18395 10935 18398
rect 13537 18458 13603 18461
rect 17033 18458 17099 18461
rect 13537 18456 17099 18458
rect 13537 18400 13542 18456
rect 13598 18400 17038 18456
rect 17094 18400 17099 18456
rect 13537 18398 17099 18400
rect 13537 18395 13603 18398
rect 17033 18395 17099 18398
rect 4654 18260 4660 18324
rect 4724 18322 4730 18324
rect 8661 18322 8727 18325
rect 4724 18320 8727 18322
rect 4724 18264 8666 18320
rect 8722 18264 8727 18320
rect 4724 18262 8727 18264
rect 4724 18260 4730 18262
rect 8661 18259 8727 18262
rect 11094 18260 11100 18324
rect 11164 18322 11170 18324
rect 13077 18322 13143 18325
rect 11164 18320 13143 18322
rect 11164 18264 13082 18320
rect 13138 18264 13143 18320
rect 11164 18262 13143 18264
rect 11164 18260 11170 18262
rect 13077 18259 13143 18262
rect 5257 18186 5323 18189
rect 7046 18186 7052 18188
rect 5257 18184 7052 18186
rect 5257 18128 5262 18184
rect 5318 18128 7052 18184
rect 5257 18126 7052 18128
rect 5257 18123 5323 18126
rect 7046 18124 7052 18126
rect 7116 18124 7122 18188
rect 10041 18186 10107 18189
rect 13629 18186 13695 18189
rect 10041 18184 13695 18186
rect 10041 18128 10046 18184
rect 10102 18128 13634 18184
rect 13690 18128 13695 18184
rect 10041 18126 13695 18128
rect 10041 18123 10107 18126
rect 13629 18123 13695 18126
rect 15285 18186 15351 18189
rect 15745 18186 15811 18189
rect 15285 18184 15811 18186
rect 15285 18128 15290 18184
rect 15346 18128 15750 18184
rect 15806 18128 15811 18184
rect 15285 18126 15811 18128
rect 15285 18123 15351 18126
rect 15745 18123 15811 18126
rect 13486 17988 13492 18052
rect 13556 18050 13562 18052
rect 15101 18050 15167 18053
rect 13556 18048 15167 18050
rect 13556 17992 15106 18048
rect 15162 17992 15167 18048
rect 13556 17990 15167 17992
rect 13556 17988 13562 17990
rect 15101 17987 15167 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 7649 17916 7715 17917
rect 7598 17914 7604 17916
rect 7558 17854 7604 17914
rect 7668 17912 7715 17916
rect 7710 17856 7715 17912
rect 7598 17852 7604 17854
rect 7668 17852 7715 17856
rect 7649 17851 7715 17852
rect 8753 17914 8819 17917
rect 10593 17914 10659 17917
rect 8753 17912 10659 17914
rect 8753 17856 8758 17912
rect 8814 17856 10598 17912
rect 10654 17856 10659 17912
rect 8753 17854 10659 17856
rect 8753 17851 8819 17854
rect 10593 17851 10659 17854
rect 13077 17914 13143 17917
rect 16021 17914 16087 17917
rect 13077 17912 16087 17914
rect 13077 17856 13082 17912
rect 13138 17856 16026 17912
rect 16082 17856 16087 17912
rect 13077 17854 16087 17856
rect 13077 17851 13143 17854
rect 16021 17851 16087 17854
rect 2630 17716 2636 17780
rect 2700 17778 2706 17780
rect 4705 17778 4771 17781
rect 2700 17776 4771 17778
rect 2700 17720 4710 17776
rect 4766 17720 4771 17776
rect 2700 17718 4771 17720
rect 2700 17716 2706 17718
rect 4705 17715 4771 17718
rect 10041 17778 10107 17781
rect 10869 17778 10935 17781
rect 10041 17776 10935 17778
rect 10041 17720 10046 17776
rect 10102 17720 10874 17776
rect 10930 17720 10935 17776
rect 10041 17718 10935 17720
rect 10041 17715 10107 17718
rect 10869 17715 10935 17718
rect 38285 17778 38351 17781
rect 39200 17778 39800 17808
rect 38285 17776 39800 17778
rect 38285 17720 38290 17776
rect 38346 17720 39800 17776
rect 38285 17718 39800 17720
rect 38285 17715 38351 17718
rect 39200 17688 39800 17718
rect 3969 17644 4035 17645
rect 3918 17642 3924 17644
rect 3878 17582 3924 17642
rect 3988 17640 4035 17644
rect 4030 17584 4035 17640
rect 3918 17580 3924 17582
rect 3988 17580 4035 17584
rect 3969 17579 4035 17580
rect 4245 17642 4311 17645
rect 4521 17642 4587 17645
rect 12433 17642 12499 17645
rect 17309 17642 17375 17645
rect 4245 17640 17375 17642
rect 4245 17584 4250 17640
rect 4306 17584 4526 17640
rect 4582 17584 12438 17640
rect 12494 17584 17314 17640
rect 17370 17584 17375 17640
rect 4245 17582 17375 17584
rect 4245 17579 4311 17582
rect 4521 17579 4587 17582
rect 12433 17579 12499 17582
rect 17309 17579 17375 17582
rect 19885 17642 19951 17645
rect 21173 17642 21239 17645
rect 19885 17640 21239 17642
rect 19885 17584 19890 17640
rect 19946 17584 21178 17640
rect 21234 17584 21239 17640
rect 19885 17582 21239 17584
rect 19885 17579 19951 17582
rect 21173 17579 21239 17582
rect 1853 17506 1919 17509
rect 6177 17506 6243 17509
rect 11145 17506 11211 17509
rect 1853 17504 5090 17506
rect 1853 17448 1858 17504
rect 1914 17448 5090 17504
rect 1853 17446 5090 17448
rect 1853 17443 1919 17446
rect 841 17370 907 17373
rect 4797 17370 4863 17373
rect 841 17368 4863 17370
rect 841 17312 846 17368
rect 902 17312 4802 17368
rect 4858 17312 4863 17368
rect 841 17310 4863 17312
rect 5030 17370 5090 17446
rect 6177 17504 11211 17506
rect 6177 17448 6182 17504
rect 6238 17448 11150 17504
rect 11206 17448 11211 17504
rect 6177 17446 11211 17448
rect 6177 17443 6243 17446
rect 11145 17443 11211 17446
rect 16113 17506 16179 17509
rect 16665 17506 16731 17509
rect 16113 17504 16731 17506
rect 16113 17448 16118 17504
rect 16174 17448 16670 17504
rect 16726 17448 16731 17504
rect 16113 17446 16731 17448
rect 16113 17443 16179 17446
rect 16665 17443 16731 17446
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 9121 17370 9187 17373
rect 5030 17368 9187 17370
rect 5030 17312 9126 17368
rect 9182 17312 9187 17368
rect 5030 17310 9187 17312
rect 841 17307 907 17310
rect 4797 17307 4863 17310
rect 9121 17307 9187 17310
rect 10685 17370 10751 17373
rect 11145 17370 11211 17373
rect 10685 17368 11211 17370
rect 10685 17312 10690 17368
rect 10746 17312 11150 17368
rect 11206 17312 11211 17368
rect 10685 17310 11211 17312
rect 10685 17307 10751 17310
rect 11145 17307 11211 17310
rect 13721 17370 13787 17373
rect 17677 17370 17743 17373
rect 13721 17368 17743 17370
rect 13721 17312 13726 17368
rect 13782 17312 17682 17368
rect 17738 17312 17743 17368
rect 13721 17310 17743 17312
rect 13721 17307 13787 17310
rect 17677 17307 17743 17310
rect 7046 17172 7052 17236
rect 7116 17234 7122 17236
rect 12566 17234 12572 17236
rect 7116 17174 12572 17234
rect 7116 17172 7122 17174
rect 12566 17172 12572 17174
rect 12636 17172 12642 17236
rect 13353 17234 13419 17237
rect 17309 17234 17375 17237
rect 13353 17232 17375 17234
rect 13353 17176 13358 17232
rect 13414 17176 17314 17232
rect 17370 17176 17375 17232
rect 13353 17174 17375 17176
rect 13353 17171 13419 17174
rect 17309 17171 17375 17174
rect 200 17098 800 17128
rect 2773 17098 2839 17101
rect 200 17096 2839 17098
rect 200 17040 2778 17096
rect 2834 17040 2839 17096
rect 200 17038 2839 17040
rect 200 17008 800 17038
rect 2773 17035 2839 17038
rect 19333 17098 19399 17101
rect 19701 17098 19767 17101
rect 19333 17096 19767 17098
rect 19333 17040 19338 17096
rect 19394 17040 19706 17096
rect 19762 17040 19767 17096
rect 19333 17038 19767 17040
rect 19333 17035 19399 17038
rect 19701 17035 19767 17038
rect 11881 16962 11947 16965
rect 12341 16962 12407 16965
rect 11881 16960 12407 16962
rect 11881 16904 11886 16960
rect 11942 16904 12346 16960
rect 12402 16904 12407 16960
rect 11881 16902 12407 16904
rect 11881 16899 11947 16902
rect 12341 16899 12407 16902
rect 14273 16962 14339 16965
rect 18965 16962 19031 16965
rect 14273 16960 19031 16962
rect 14273 16904 14278 16960
rect 14334 16904 18970 16960
rect 19026 16904 19031 16960
rect 14273 16902 19031 16904
rect 14273 16899 14339 16902
rect 18965 16899 19031 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 12341 16826 12407 16829
rect 18597 16826 18663 16829
rect 12341 16824 18663 16826
rect 12341 16768 12346 16824
rect 12402 16768 18602 16824
rect 18658 16768 18663 16824
rect 12341 16766 18663 16768
rect 12341 16763 12407 16766
rect 18597 16763 18663 16766
rect 3141 16690 3207 16693
rect 9213 16690 9279 16693
rect 3141 16688 9279 16690
rect 3141 16632 3146 16688
rect 3202 16632 9218 16688
rect 9274 16632 9279 16688
rect 3141 16630 9279 16632
rect 3141 16627 3207 16630
rect 9213 16627 9279 16630
rect 10961 16690 11027 16693
rect 17493 16690 17559 16693
rect 10961 16688 17559 16690
rect 10961 16632 10966 16688
rect 11022 16632 17498 16688
rect 17554 16632 17559 16688
rect 10961 16630 17559 16632
rect 10961 16627 11027 16630
rect 17493 16627 17559 16630
rect 9305 16554 9371 16557
rect 9438 16554 9444 16556
rect 9305 16552 9444 16554
rect 9305 16496 9310 16552
rect 9366 16496 9444 16552
rect 9305 16494 9444 16496
rect 9305 16491 9371 16494
rect 9438 16492 9444 16494
rect 9508 16492 9514 16556
rect 12525 16554 12591 16557
rect 20253 16554 20319 16557
rect 12525 16552 20319 16554
rect 12525 16496 12530 16552
rect 12586 16496 20258 16552
rect 20314 16496 20319 16552
rect 12525 16494 20319 16496
rect 12525 16491 12591 16494
rect 20253 16491 20319 16494
rect 2221 16418 2287 16421
rect 2865 16418 2931 16421
rect 2221 16416 2931 16418
rect 2221 16360 2226 16416
rect 2282 16360 2870 16416
rect 2926 16360 2931 16416
rect 2221 16358 2931 16360
rect 2221 16355 2287 16358
rect 2865 16355 2931 16358
rect 4061 16418 4127 16421
rect 7465 16418 7531 16421
rect 9121 16420 9187 16421
rect 4061 16416 7531 16418
rect 4061 16360 4066 16416
rect 4122 16360 7470 16416
rect 7526 16360 7531 16416
rect 4061 16358 7531 16360
rect 4061 16355 4127 16358
rect 7465 16355 7531 16358
rect 9070 16356 9076 16420
rect 9140 16418 9187 16420
rect 12249 16418 12315 16421
rect 16297 16418 16363 16421
rect 9140 16416 9232 16418
rect 9182 16360 9232 16416
rect 9140 16358 9232 16360
rect 12249 16416 16363 16418
rect 12249 16360 12254 16416
rect 12310 16360 16302 16416
rect 16358 16360 16363 16416
rect 12249 16358 16363 16360
rect 9140 16356 9187 16358
rect 9121 16355 9187 16356
rect 12249 16355 12315 16358
rect 16297 16355 16363 16358
rect 38193 16418 38259 16421
rect 39200 16418 39800 16448
rect 38193 16416 39800 16418
rect 38193 16360 38198 16416
rect 38254 16360 39800 16416
rect 38193 16358 39800 16360
rect 38193 16355 38259 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 39200 16328 39800 16358
rect 19570 16287 19886 16288
rect 3509 16282 3575 16285
rect 5533 16282 5599 16285
rect 3509 16280 5599 16282
rect 3509 16224 3514 16280
rect 3570 16224 5538 16280
rect 5594 16224 5599 16280
rect 3509 16222 5599 16224
rect 3509 16219 3575 16222
rect 5533 16219 5599 16222
rect 13261 16282 13327 16285
rect 15561 16282 15627 16285
rect 13261 16280 15627 16282
rect 13261 16224 13266 16280
rect 13322 16224 15566 16280
rect 15622 16224 15627 16280
rect 13261 16222 15627 16224
rect 13261 16219 13327 16222
rect 15561 16219 15627 16222
rect 5165 16146 5231 16149
rect 5809 16146 5875 16149
rect 5165 16144 5875 16146
rect 5165 16088 5170 16144
rect 5226 16088 5814 16144
rect 5870 16088 5875 16144
rect 5165 16086 5875 16088
rect 5165 16083 5231 16086
rect 5809 16083 5875 16086
rect 7414 16084 7420 16148
rect 7484 16146 7490 16148
rect 15193 16146 15259 16149
rect 7484 16144 15259 16146
rect 7484 16088 15198 16144
rect 15254 16088 15259 16144
rect 7484 16086 15259 16088
rect 7484 16084 7490 16086
rect 15193 16083 15259 16086
rect 3325 16010 3391 16013
rect 8753 16010 8819 16013
rect 3325 16008 8819 16010
rect 3325 15952 3330 16008
rect 3386 15952 8758 16008
rect 8814 15952 8819 16008
rect 3325 15950 8819 15952
rect 3325 15947 3391 15950
rect 8753 15947 8819 15950
rect 9305 16010 9371 16013
rect 16430 16010 16436 16012
rect 9305 16008 16436 16010
rect 9305 15952 9310 16008
rect 9366 15952 16436 16008
rect 9305 15950 16436 15952
rect 9305 15947 9371 15950
rect 16430 15948 16436 15950
rect 16500 15948 16506 16012
rect 14457 15874 14523 15877
rect 15929 15874 15995 15877
rect 14457 15872 15995 15874
rect 14457 15816 14462 15872
rect 14518 15816 15934 15872
rect 15990 15816 15995 15872
rect 14457 15814 15995 15816
rect 14457 15811 14523 15814
rect 15929 15811 15995 15814
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 2773 15738 2839 15741
rect 200 15736 2839 15738
rect 200 15680 2778 15736
rect 2834 15680 2839 15736
rect 200 15678 2839 15680
rect 200 15648 800 15678
rect 2773 15675 2839 15678
rect 8385 15738 8451 15741
rect 8886 15738 8892 15740
rect 8385 15736 8892 15738
rect 8385 15680 8390 15736
rect 8446 15680 8892 15736
rect 8385 15678 8892 15680
rect 8385 15675 8451 15678
rect 8886 15676 8892 15678
rect 8956 15676 8962 15740
rect 9121 15738 9187 15741
rect 9254 15738 9260 15740
rect 9121 15736 9260 15738
rect 9121 15680 9126 15736
rect 9182 15680 9260 15736
rect 9121 15678 9260 15680
rect 9121 15675 9187 15678
rect 9254 15676 9260 15678
rect 9324 15676 9330 15740
rect 10409 15738 10475 15741
rect 12893 15738 12959 15741
rect 15285 15738 15351 15741
rect 10409 15736 15351 15738
rect 10409 15680 10414 15736
rect 10470 15680 12898 15736
rect 12954 15680 15290 15736
rect 15346 15680 15351 15736
rect 10409 15678 15351 15680
rect 10409 15675 10475 15678
rect 12893 15675 12959 15678
rect 15285 15675 15351 15678
rect 38285 15738 38351 15741
rect 39200 15738 39800 15768
rect 38285 15736 39800 15738
rect 38285 15680 38290 15736
rect 38346 15680 39800 15736
rect 38285 15678 39800 15680
rect 38285 15675 38351 15678
rect 39200 15648 39800 15678
rect 3969 15602 4035 15605
rect 5441 15602 5507 15605
rect 3969 15600 5507 15602
rect 3969 15544 3974 15600
rect 4030 15544 5446 15600
rect 5502 15544 5507 15600
rect 3969 15542 5507 15544
rect 3969 15539 4035 15542
rect 5441 15539 5507 15542
rect 6729 15602 6795 15605
rect 12065 15602 12131 15605
rect 6729 15600 12131 15602
rect 6729 15544 6734 15600
rect 6790 15544 12070 15600
rect 12126 15544 12131 15600
rect 6729 15542 12131 15544
rect 6729 15539 6795 15542
rect 12065 15539 12131 15542
rect 20253 15602 20319 15605
rect 20437 15602 20503 15605
rect 20253 15600 20503 15602
rect 20253 15544 20258 15600
rect 20314 15544 20442 15600
rect 20498 15544 20503 15600
rect 20253 15542 20503 15544
rect 20253 15539 20319 15542
rect 20437 15539 20503 15542
rect 12801 15466 12867 15469
rect 13721 15466 13787 15469
rect 15101 15466 15167 15469
rect 12801 15464 15167 15466
rect 12801 15408 12806 15464
rect 12862 15408 13726 15464
rect 13782 15408 15106 15464
rect 15162 15408 15167 15464
rect 12801 15406 15167 15408
rect 12801 15403 12867 15406
rect 13721 15403 13787 15406
rect 15101 15403 15167 15406
rect 16389 15466 16455 15469
rect 22369 15466 22435 15469
rect 16389 15464 22435 15466
rect 16389 15408 16394 15464
rect 16450 15408 22374 15464
rect 22430 15408 22435 15464
rect 16389 15406 22435 15408
rect 16389 15403 16455 15406
rect 22369 15403 22435 15406
rect 4061 15330 4127 15333
rect 7189 15330 7255 15333
rect 4061 15328 7255 15330
rect 4061 15272 4066 15328
rect 4122 15272 7194 15328
rect 7250 15272 7255 15328
rect 4061 15270 7255 15272
rect 4061 15267 4127 15270
rect 7189 15267 7255 15270
rect 11145 15330 11211 15333
rect 13169 15330 13235 15333
rect 11145 15328 13235 15330
rect 11145 15272 11150 15328
rect 11206 15272 13174 15328
rect 13230 15272 13235 15328
rect 11145 15270 13235 15272
rect 11145 15267 11211 15270
rect 13169 15267 13235 15270
rect 16614 15268 16620 15332
rect 16684 15330 16690 15332
rect 17677 15330 17743 15333
rect 16684 15328 17743 15330
rect 16684 15272 17682 15328
rect 17738 15272 17743 15328
rect 16684 15270 17743 15272
rect 16684 15268 16690 15270
rect 17677 15267 17743 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 5533 15196 5599 15197
rect 5533 15194 5580 15196
rect 5488 15192 5580 15194
rect 5488 15136 5538 15192
rect 5488 15134 5580 15136
rect 5533 15132 5580 15134
rect 5644 15132 5650 15196
rect 6545 15194 6611 15197
rect 9489 15194 9555 15197
rect 6545 15192 9555 15194
rect 6545 15136 6550 15192
rect 6606 15136 9494 15192
rect 9550 15136 9555 15192
rect 6545 15134 9555 15136
rect 5533 15131 5599 15132
rect 6545 15131 6611 15134
rect 9489 15131 9555 15134
rect 200 15058 800 15088
rect 3509 15058 3575 15061
rect 200 15056 3575 15058
rect 200 15000 3514 15056
rect 3570 15000 3575 15056
rect 200 14998 3575 15000
rect 200 14968 800 14998
rect 3509 14995 3575 14998
rect 7649 15058 7715 15061
rect 11830 15058 11836 15060
rect 7649 15056 11836 15058
rect 7649 15000 7654 15056
rect 7710 15000 11836 15056
rect 7649 14998 11836 15000
rect 7649 14995 7715 14998
rect 11830 14996 11836 14998
rect 11900 14996 11906 15060
rect 23289 15058 23355 15061
rect 12390 15056 23355 15058
rect 12390 15000 23294 15056
rect 23350 15000 23355 15056
rect 12390 14998 23355 15000
rect 2221 14922 2287 14925
rect 12390 14922 12450 14998
rect 23289 14995 23355 14998
rect 2221 14920 12450 14922
rect 2221 14864 2226 14920
rect 2282 14864 12450 14920
rect 2221 14862 12450 14864
rect 2221 14859 2287 14862
rect 4705 14786 4771 14789
rect 9305 14786 9371 14789
rect 4705 14784 9371 14786
rect 4705 14728 4710 14784
rect 4766 14728 9310 14784
rect 9366 14728 9371 14784
rect 4705 14726 9371 14728
rect 4705 14723 4771 14726
rect 9305 14723 9371 14726
rect 17585 14786 17651 14789
rect 17861 14786 17927 14789
rect 17585 14784 17927 14786
rect 17585 14728 17590 14784
rect 17646 14728 17866 14784
rect 17922 14728 17927 14784
rect 17585 14726 17927 14728
rect 17585 14723 17651 14726
rect 17861 14723 17927 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 5533 14650 5599 14653
rect 10542 14650 10548 14652
rect 5533 14648 10548 14650
rect 5533 14592 5538 14648
rect 5594 14592 10548 14648
rect 5533 14590 10548 14592
rect 5533 14587 5599 14590
rect 10542 14588 10548 14590
rect 10612 14588 10618 14652
rect 14549 14650 14615 14653
rect 16021 14650 16087 14653
rect 14549 14648 16087 14650
rect 14549 14592 14554 14648
rect 14610 14592 16026 14648
rect 16082 14592 16087 14648
rect 14549 14590 16087 14592
rect 14549 14587 14615 14590
rect 16021 14587 16087 14590
rect 7097 14514 7163 14517
rect 7230 14514 7236 14516
rect 7097 14512 7236 14514
rect 7097 14456 7102 14512
rect 7158 14456 7236 14512
rect 7097 14454 7236 14456
rect 7097 14451 7163 14454
rect 7230 14452 7236 14454
rect 7300 14452 7306 14516
rect 9070 14452 9076 14516
rect 9140 14514 9146 14516
rect 9305 14514 9371 14517
rect 9140 14512 9371 14514
rect 9140 14456 9310 14512
rect 9366 14456 9371 14512
rect 9140 14454 9371 14456
rect 9140 14452 9146 14454
rect 9305 14451 9371 14454
rect 2313 14378 2379 14381
rect 9397 14378 9463 14381
rect 2313 14376 9463 14378
rect 2313 14320 2318 14376
rect 2374 14320 9402 14376
rect 9458 14320 9463 14376
rect 2313 14318 9463 14320
rect 2313 14315 2379 14318
rect 9397 14315 9463 14318
rect 38193 14378 38259 14381
rect 39200 14378 39800 14408
rect 38193 14376 39800 14378
rect 38193 14320 38198 14376
rect 38254 14320 39800 14376
rect 38193 14318 39800 14320
rect 38193 14315 38259 14318
rect 39200 14288 39800 14318
rect 4654 14180 4660 14244
rect 4724 14242 4730 14244
rect 5073 14242 5139 14245
rect 4724 14240 5139 14242
rect 4724 14184 5078 14240
rect 5134 14184 5139 14240
rect 4724 14182 5139 14184
rect 4724 14180 4730 14182
rect 5073 14179 5139 14182
rect 11329 14242 11395 14245
rect 11697 14242 11763 14245
rect 18965 14242 19031 14245
rect 11329 14240 19031 14242
rect 11329 14184 11334 14240
rect 11390 14184 11702 14240
rect 11758 14184 18970 14240
rect 19026 14184 19031 14240
rect 11329 14182 19031 14184
rect 11329 14179 11395 14182
rect 11697 14179 11763 14182
rect 18965 14179 19031 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 4613 14106 4679 14109
rect 6862 14106 6868 14108
rect 4613 14104 6868 14106
rect 4613 14048 4618 14104
rect 4674 14048 6868 14104
rect 4613 14046 6868 14048
rect 4613 14043 4679 14046
rect 6862 14044 6868 14046
rect 6932 14044 6938 14108
rect 3969 13970 4035 13973
rect 8017 13970 8083 13973
rect 3969 13968 8083 13970
rect 3969 13912 3974 13968
rect 4030 13912 8022 13968
rect 8078 13912 8083 13968
rect 3969 13910 8083 13912
rect 3969 13907 4035 13910
rect 8017 13907 8083 13910
rect 10685 13970 10751 13973
rect 24669 13970 24735 13973
rect 10685 13968 24735 13970
rect 10685 13912 10690 13968
rect 10746 13912 24674 13968
rect 24730 13912 24735 13968
rect 10685 13910 24735 13912
rect 10685 13907 10751 13910
rect 24669 13907 24735 13910
rect 3693 13834 3759 13837
rect 6637 13834 6703 13837
rect 8845 13834 8911 13837
rect 3693 13832 8911 13834
rect 3693 13776 3698 13832
rect 3754 13776 6642 13832
rect 6698 13776 8850 13832
rect 8906 13776 8911 13832
rect 3693 13774 8911 13776
rect 3693 13771 3759 13774
rect 6637 13771 6703 13774
rect 8845 13771 8911 13774
rect 9949 13834 10015 13837
rect 10317 13834 10383 13837
rect 9949 13832 10383 13834
rect 9949 13776 9954 13832
rect 10010 13776 10322 13832
rect 10378 13776 10383 13832
rect 9949 13774 10383 13776
rect 9949 13771 10015 13774
rect 10317 13771 10383 13774
rect 11830 13772 11836 13836
rect 11900 13834 11906 13836
rect 14273 13834 14339 13837
rect 11900 13832 14339 13834
rect 11900 13776 14278 13832
rect 14334 13776 14339 13832
rect 11900 13774 14339 13776
rect 11900 13772 11906 13774
rect 14273 13771 14339 13774
rect 17677 13834 17743 13837
rect 19517 13834 19583 13837
rect 17677 13832 19583 13834
rect 17677 13776 17682 13832
rect 17738 13776 19522 13832
rect 19578 13776 19583 13832
rect 17677 13774 19583 13776
rect 17677 13771 17743 13774
rect 19517 13771 19583 13774
rect 200 13698 800 13728
rect 2773 13698 2839 13701
rect 200 13696 2839 13698
rect 200 13640 2778 13696
rect 2834 13640 2839 13696
rect 200 13638 2839 13640
rect 200 13608 800 13638
rect 2773 13635 2839 13638
rect 5257 13698 5323 13701
rect 8753 13698 8819 13701
rect 5257 13696 8819 13698
rect 5257 13640 5262 13696
rect 5318 13640 8758 13696
rect 8814 13640 8819 13696
rect 5257 13638 8819 13640
rect 5257 13635 5323 13638
rect 8753 13635 8819 13638
rect 10777 13698 10843 13701
rect 12525 13698 12591 13701
rect 10777 13696 12591 13698
rect 10777 13640 10782 13696
rect 10838 13640 12530 13696
rect 12586 13640 12591 13696
rect 10777 13638 12591 13640
rect 10777 13635 10843 13638
rect 12525 13635 12591 13638
rect 17125 13698 17191 13701
rect 18781 13698 18847 13701
rect 17125 13696 18847 13698
rect 17125 13640 17130 13696
rect 17186 13640 18786 13696
rect 18842 13640 18847 13696
rect 17125 13638 18847 13640
rect 17125 13635 17191 13638
rect 18781 13635 18847 13638
rect 18965 13698 19031 13701
rect 20253 13698 20319 13701
rect 18965 13696 20319 13698
rect 18965 13640 18970 13696
rect 19026 13640 20258 13696
rect 20314 13640 20319 13696
rect 18965 13638 20319 13640
rect 18965 13635 19031 13638
rect 20253 13635 20319 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 12709 13562 12775 13565
rect 19149 13562 19215 13565
rect 12709 13560 19215 13562
rect 12709 13504 12714 13560
rect 12770 13504 19154 13560
rect 19210 13504 19215 13560
rect 12709 13502 19215 13504
rect 12709 13499 12775 13502
rect 19149 13499 19215 13502
rect 19885 13562 19951 13565
rect 23473 13562 23539 13565
rect 19885 13560 23539 13562
rect 19885 13504 19890 13560
rect 19946 13504 23478 13560
rect 23534 13504 23539 13560
rect 19885 13502 23539 13504
rect 19885 13499 19951 13502
rect 23473 13499 23539 13502
rect 974 13364 980 13428
rect 1044 13426 1050 13428
rect 4337 13426 4403 13429
rect 1044 13424 4403 13426
rect 1044 13368 4342 13424
rect 4398 13368 4403 13424
rect 1044 13366 4403 13368
rect 1044 13364 1050 13366
rect 4337 13363 4403 13366
rect 6269 13426 6335 13429
rect 8385 13426 8451 13429
rect 6269 13424 8451 13426
rect 6269 13368 6274 13424
rect 6330 13368 8390 13424
rect 8446 13368 8451 13424
rect 6269 13366 8451 13368
rect 6269 13363 6335 13366
rect 8385 13363 8451 13366
rect 10685 13426 10751 13429
rect 13445 13426 13511 13429
rect 10685 13424 13511 13426
rect 10685 13368 10690 13424
rect 10746 13368 13450 13424
rect 13506 13368 13511 13424
rect 10685 13366 13511 13368
rect 10685 13363 10751 13366
rect 13445 13363 13511 13366
rect 16430 13364 16436 13428
rect 16500 13426 16506 13428
rect 22093 13426 22159 13429
rect 16500 13424 22159 13426
rect 16500 13368 22098 13424
rect 22154 13368 22159 13424
rect 16500 13366 22159 13368
rect 16500 13364 16506 13366
rect 22093 13363 22159 13366
rect 3969 13290 4035 13293
rect 10174 13290 10180 13292
rect 3969 13288 10180 13290
rect 3969 13232 3974 13288
rect 4030 13232 10180 13288
rect 3969 13230 10180 13232
rect 3969 13227 4035 13230
rect 10174 13228 10180 13230
rect 10244 13228 10250 13292
rect 13997 13290 14063 13293
rect 27061 13290 27127 13293
rect 13997 13288 27127 13290
rect 13997 13232 14002 13288
rect 14058 13232 27066 13288
rect 27122 13232 27127 13288
rect 13997 13230 27127 13232
rect 13997 13227 14063 13230
rect 27061 13227 27127 13230
rect 12341 13154 12407 13157
rect 14825 13154 14891 13157
rect 12341 13152 14891 13154
rect 12341 13096 12346 13152
rect 12402 13096 14830 13152
rect 14886 13096 14891 13152
rect 12341 13094 14891 13096
rect 12341 13091 12407 13094
rect 14825 13091 14891 13094
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 17953 13018 18019 13021
rect 19241 13018 19307 13021
rect 17953 13016 19307 13018
rect 17953 12960 17958 13016
rect 18014 12960 19246 13016
rect 19302 12960 19307 13016
rect 17953 12958 19307 12960
rect 17953 12955 18019 12958
rect 19241 12955 19307 12958
rect 38193 13018 38259 13021
rect 39200 13018 39800 13048
rect 38193 13016 39800 13018
rect 38193 12960 38198 13016
rect 38254 12960 39800 13016
rect 38193 12958 39800 12960
rect 38193 12955 38259 12958
rect 39200 12928 39800 12958
rect 10225 12882 10291 12885
rect 12433 12882 12499 12885
rect 13077 12884 13143 12885
rect 13077 12882 13124 12884
rect 10225 12880 12499 12882
rect 10225 12824 10230 12880
rect 10286 12824 12438 12880
rect 12494 12824 12499 12880
rect 10225 12822 12499 12824
rect 13032 12880 13124 12882
rect 13032 12824 13082 12880
rect 13032 12822 13124 12824
rect 10225 12819 10291 12822
rect 12433 12819 12499 12822
rect 13077 12820 13124 12822
rect 13188 12820 13194 12884
rect 17309 12882 17375 12885
rect 18597 12882 18663 12885
rect 17309 12880 18663 12882
rect 17309 12824 17314 12880
rect 17370 12824 18602 12880
rect 18658 12824 18663 12880
rect 17309 12822 18663 12824
rect 13077 12819 13143 12820
rect 17309 12819 17375 12822
rect 18597 12819 18663 12822
rect 3969 12746 4035 12749
rect 4245 12746 4311 12749
rect 3969 12744 4311 12746
rect 3969 12688 3974 12744
rect 4030 12688 4250 12744
rect 4306 12688 4311 12744
rect 3969 12686 4311 12688
rect 3969 12683 4035 12686
rect 4245 12683 4311 12686
rect 5625 12746 5691 12749
rect 5758 12746 5764 12748
rect 5625 12744 5764 12746
rect 5625 12688 5630 12744
rect 5686 12688 5764 12744
rect 5625 12686 5764 12688
rect 5625 12683 5691 12686
rect 5758 12684 5764 12686
rect 5828 12684 5834 12748
rect 13261 12746 13327 12749
rect 13629 12746 13695 12749
rect 13261 12744 13695 12746
rect 13261 12688 13266 12744
rect 13322 12688 13634 12744
rect 13690 12688 13695 12744
rect 13261 12686 13695 12688
rect 13261 12683 13327 12686
rect 13629 12683 13695 12686
rect 17217 12746 17283 12749
rect 17585 12746 17651 12749
rect 38193 12746 38259 12749
rect 17217 12744 17651 12746
rect 17217 12688 17222 12744
rect 17278 12688 17590 12744
rect 17646 12688 17651 12744
rect 17217 12686 17651 12688
rect 17217 12683 17283 12686
rect 17585 12683 17651 12686
rect 22050 12744 38259 12746
rect 22050 12688 38198 12744
rect 38254 12688 38259 12744
rect 22050 12686 38259 12688
rect 13169 12610 13235 12613
rect 20069 12610 20135 12613
rect 20437 12610 20503 12613
rect 13169 12608 13370 12610
rect 13169 12552 13174 12608
rect 13230 12552 13370 12608
rect 13169 12550 13370 12552
rect 13169 12547 13235 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 4981 12474 5047 12477
rect 7557 12474 7623 12477
rect 13169 12476 13235 12477
rect 13118 12474 13124 12476
rect 4981 12472 7623 12474
rect 4981 12416 4986 12472
rect 5042 12416 7562 12472
rect 7618 12416 7623 12472
rect 4981 12414 7623 12416
rect 13078 12414 13124 12474
rect 13188 12472 13235 12476
rect 13230 12416 13235 12472
rect 4981 12411 5047 12414
rect 7557 12411 7623 12414
rect 13118 12412 13124 12414
rect 13188 12412 13235 12416
rect 13310 12474 13370 12550
rect 20069 12608 20503 12610
rect 20069 12552 20074 12608
rect 20130 12552 20442 12608
rect 20498 12552 20503 12608
rect 20069 12550 20503 12552
rect 20069 12547 20135 12550
rect 20437 12547 20503 12550
rect 13537 12474 13603 12477
rect 22050 12474 22110 12686
rect 38193 12683 38259 12686
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 13310 12472 13603 12474
rect 13310 12416 13542 12472
rect 13598 12416 13603 12472
rect 13310 12414 13603 12416
rect 13169 12411 13235 12412
rect 13537 12411 13603 12414
rect 20670 12414 22110 12474
rect 200 12338 800 12368
rect 3141 12340 3207 12341
rect 200 12278 2790 12338
rect 200 12248 800 12278
rect 2730 12202 2790 12278
rect 3141 12336 3188 12340
rect 3252 12338 3258 12340
rect 8201 12338 8267 12341
rect 11329 12338 11395 12341
rect 3141 12280 3146 12336
rect 3141 12276 3188 12280
rect 3252 12278 3298 12338
rect 8201 12336 11395 12338
rect 8201 12280 8206 12336
rect 8262 12280 11334 12336
rect 11390 12280 11395 12336
rect 8201 12278 11395 12280
rect 3252 12276 3258 12278
rect 3141 12275 3207 12276
rect 8201 12275 8267 12278
rect 11329 12275 11395 12278
rect 14641 12338 14707 12341
rect 16573 12338 16639 12341
rect 14641 12336 16639 12338
rect 14641 12280 14646 12336
rect 14702 12280 16578 12336
rect 16634 12280 16639 12336
rect 14641 12278 16639 12280
rect 14641 12275 14707 12278
rect 16573 12275 16639 12278
rect 19425 12338 19491 12341
rect 20110 12338 20116 12340
rect 19425 12336 20116 12338
rect 19425 12280 19430 12336
rect 19486 12280 20116 12336
rect 19425 12278 20116 12280
rect 19425 12275 19491 12278
rect 20110 12276 20116 12278
rect 20180 12338 20186 12340
rect 20670 12338 20730 12414
rect 20180 12278 20730 12338
rect 38101 12338 38167 12341
rect 39200 12338 39800 12368
rect 38101 12336 39800 12338
rect 38101 12280 38106 12336
rect 38162 12280 39800 12336
rect 38101 12278 39800 12280
rect 20180 12276 20186 12278
rect 38101 12275 38167 12278
rect 39200 12248 39800 12278
rect 3693 12202 3759 12205
rect 2730 12200 3759 12202
rect 2730 12144 3698 12200
rect 3754 12144 3759 12200
rect 2730 12142 3759 12144
rect 3693 12139 3759 12142
rect 14549 12202 14615 12205
rect 19977 12202 20043 12205
rect 14549 12200 20043 12202
rect 14549 12144 14554 12200
rect 14610 12144 19982 12200
rect 20038 12144 20043 12200
rect 14549 12142 20043 12144
rect 14549 12139 14615 12142
rect 19977 12139 20043 12142
rect 10961 12066 11027 12069
rect 13261 12066 13327 12069
rect 10961 12064 13327 12066
rect 10961 12008 10966 12064
rect 11022 12008 13266 12064
rect 13322 12008 13327 12064
rect 10961 12006 13327 12008
rect 10961 12003 11027 12006
rect 13261 12003 13327 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 12617 11930 12683 11933
rect 15837 11930 15903 11933
rect 12617 11928 15903 11930
rect 12617 11872 12622 11928
rect 12678 11872 15842 11928
rect 15898 11872 15903 11928
rect 12617 11870 15903 11872
rect 12617 11867 12683 11870
rect 15837 11867 15903 11870
rect 6821 11794 6887 11797
rect 23289 11794 23355 11797
rect 6821 11792 23355 11794
rect 6821 11736 6826 11792
rect 6882 11736 23294 11792
rect 23350 11736 23355 11792
rect 6821 11734 23355 11736
rect 6821 11731 6887 11734
rect 23289 11731 23355 11734
rect 200 11658 800 11688
rect 2773 11658 2839 11661
rect 200 11656 2839 11658
rect 200 11600 2778 11656
rect 2834 11600 2839 11656
rect 200 11598 2839 11600
rect 200 11568 800 11598
rect 2773 11595 2839 11598
rect 3417 11658 3483 11661
rect 6494 11658 6500 11660
rect 3417 11656 6500 11658
rect 3417 11600 3422 11656
rect 3478 11600 6500 11656
rect 3417 11598 6500 11600
rect 3417 11595 3483 11598
rect 6494 11596 6500 11598
rect 6564 11658 6570 11660
rect 8017 11658 8083 11661
rect 6564 11656 8083 11658
rect 6564 11600 8022 11656
rect 8078 11600 8083 11656
rect 6564 11598 8083 11600
rect 6564 11596 6570 11598
rect 8017 11595 8083 11598
rect 9673 11658 9739 11661
rect 12065 11658 12131 11661
rect 9673 11656 12131 11658
rect 9673 11600 9678 11656
rect 9734 11600 12070 11656
rect 12126 11600 12131 11656
rect 9673 11598 12131 11600
rect 9673 11595 9739 11598
rect 12065 11595 12131 11598
rect 12433 11658 12499 11661
rect 12433 11656 15026 11658
rect 12433 11600 12438 11656
rect 12494 11600 15026 11656
rect 12433 11598 15026 11600
rect 12433 11595 12499 11598
rect 6637 11524 6703 11525
rect 6637 11520 6684 11524
rect 6748 11522 6754 11524
rect 8937 11522 9003 11525
rect 11973 11522 12039 11525
rect 6637 11464 6642 11520
rect 6637 11460 6684 11464
rect 6748 11462 6794 11522
rect 8937 11520 12039 11522
rect 8937 11464 8942 11520
rect 8998 11464 11978 11520
rect 12034 11464 12039 11520
rect 8937 11462 12039 11464
rect 6748 11460 6754 11462
rect 6637 11459 6703 11460
rect 8937 11459 9003 11462
rect 11973 11459 12039 11462
rect 12157 11522 12223 11525
rect 12433 11522 12499 11525
rect 12157 11520 12499 11522
rect 12157 11464 12162 11520
rect 12218 11464 12438 11520
rect 12494 11464 12499 11520
rect 12157 11462 12499 11464
rect 14966 11522 15026 11598
rect 15510 11596 15516 11660
rect 15580 11658 15586 11660
rect 15653 11658 15719 11661
rect 15580 11656 15719 11658
rect 15580 11600 15658 11656
rect 15714 11600 15719 11656
rect 15580 11598 15719 11600
rect 15580 11596 15586 11598
rect 15653 11595 15719 11598
rect 17902 11596 17908 11660
rect 17972 11658 17978 11660
rect 22001 11658 22067 11661
rect 23013 11658 23079 11661
rect 17972 11656 23079 11658
rect 17972 11600 22006 11656
rect 22062 11600 23018 11656
rect 23074 11600 23079 11656
rect 17972 11598 23079 11600
rect 17972 11596 17978 11598
rect 22001 11595 22067 11598
rect 23013 11595 23079 11598
rect 17033 11522 17099 11525
rect 14966 11520 17099 11522
rect 14966 11464 17038 11520
rect 17094 11464 17099 11520
rect 14966 11462 17099 11464
rect 12157 11459 12223 11462
rect 12433 11459 12499 11462
rect 17033 11459 17099 11462
rect 19241 11522 19307 11525
rect 21725 11522 21791 11525
rect 19241 11520 21791 11522
rect 19241 11464 19246 11520
rect 19302 11464 21730 11520
rect 21786 11464 21791 11520
rect 19241 11462 21791 11464
rect 19241 11459 19307 11462
rect 21725 11459 21791 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 9765 11386 9831 11389
rect 11421 11386 11487 11389
rect 13813 11386 13879 11389
rect 18229 11386 18295 11389
rect 9765 11384 18295 11386
rect 9765 11328 9770 11384
rect 9826 11328 11426 11384
rect 11482 11328 13818 11384
rect 13874 11328 18234 11384
rect 18290 11328 18295 11384
rect 9765 11326 18295 11328
rect 9765 11323 9831 11326
rect 11421 11323 11487 11326
rect 13813 11323 13879 11326
rect 18229 11323 18295 11326
rect 20253 11386 20319 11389
rect 21909 11386 21975 11389
rect 20253 11384 21975 11386
rect 20253 11328 20258 11384
rect 20314 11328 21914 11384
rect 21970 11328 21975 11384
rect 20253 11326 21975 11328
rect 20253 11323 20319 11326
rect 21909 11323 21975 11326
rect 4889 11250 4955 11253
rect 4662 11248 4955 11250
rect 4662 11192 4894 11248
rect 4950 11192 4955 11248
rect 4662 11190 4955 11192
rect 4662 11117 4722 11190
rect 4889 11187 4955 11190
rect 14089 11250 14155 11253
rect 19425 11250 19491 11253
rect 20621 11250 20687 11253
rect 14089 11248 20687 11250
rect 14089 11192 14094 11248
rect 14150 11192 19430 11248
rect 19486 11192 20626 11248
rect 20682 11192 20687 11248
rect 14089 11190 20687 11192
rect 14089 11187 14155 11190
rect 19425 11187 19491 11190
rect 20621 11187 20687 11190
rect 4613 11112 4722 11117
rect 4613 11056 4618 11112
rect 4674 11056 4722 11112
rect 4613 11054 4722 11056
rect 9305 11114 9371 11117
rect 14641 11114 14707 11117
rect 9305 11112 14707 11114
rect 9305 11056 9310 11112
rect 9366 11056 14646 11112
rect 14702 11056 14707 11112
rect 9305 11054 14707 11056
rect 4613 11051 4679 11054
rect 9305 11051 9371 11054
rect 14641 11051 14707 11054
rect 22001 11114 22067 11117
rect 25129 11114 25195 11117
rect 22001 11112 25195 11114
rect 22001 11056 22006 11112
rect 22062 11056 25134 11112
rect 25190 11056 25195 11112
rect 22001 11054 25195 11056
rect 22001 11051 22067 11054
rect 23384 10981 23444 11054
rect 25129 11051 25195 11054
rect 9673 10978 9739 10981
rect 16941 10978 17007 10981
rect 9673 10976 17007 10978
rect 9673 10920 9678 10976
rect 9734 10920 16946 10976
rect 17002 10920 17007 10976
rect 9673 10918 17007 10920
rect 9673 10915 9739 10918
rect 16941 10915 17007 10918
rect 23381 10976 23447 10981
rect 23381 10920 23386 10976
rect 23442 10920 23447 10976
rect 23381 10915 23447 10920
rect 37181 10978 37247 10981
rect 39200 10978 39800 11008
rect 37181 10976 39800 10978
rect 37181 10920 37186 10976
rect 37242 10920 39800 10976
rect 37181 10918 39800 10920
rect 37181 10915 37247 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 39200 10888 39800 10918
rect 19570 10847 19886 10848
rect 8293 10842 8359 10845
rect 15009 10842 15075 10845
rect 8293 10840 15075 10842
rect 8293 10784 8298 10840
rect 8354 10784 15014 10840
rect 15070 10784 15075 10840
rect 8293 10782 15075 10784
rect 8293 10779 8359 10782
rect 15009 10779 15075 10782
rect 15929 10842 15995 10845
rect 18597 10842 18663 10845
rect 15929 10840 18663 10842
rect 15929 10784 15934 10840
rect 15990 10784 18602 10840
rect 18658 10784 18663 10840
rect 15929 10782 18663 10784
rect 15929 10779 15995 10782
rect 18597 10779 18663 10782
rect 5441 10706 5507 10709
rect 20253 10706 20319 10709
rect 5441 10704 20319 10706
rect 5441 10648 5446 10704
rect 5502 10648 20258 10704
rect 20314 10648 20319 10704
rect 5441 10646 20319 10648
rect 5441 10643 5507 10646
rect 20253 10643 20319 10646
rect 6729 10570 6795 10573
rect 9438 10570 9444 10572
rect 6729 10568 9444 10570
rect 6729 10512 6734 10568
rect 6790 10512 9444 10568
rect 6729 10510 9444 10512
rect 6729 10507 6795 10510
rect 9438 10508 9444 10510
rect 9508 10570 9514 10572
rect 9581 10570 9647 10573
rect 9508 10568 9647 10570
rect 9508 10512 9586 10568
rect 9642 10512 9647 10568
rect 9508 10510 9647 10512
rect 9508 10508 9514 10510
rect 9581 10507 9647 10510
rect 10593 10570 10659 10573
rect 11881 10570 11947 10573
rect 10593 10568 11947 10570
rect 10593 10512 10598 10568
rect 10654 10512 11886 10568
rect 11942 10512 11947 10568
rect 10593 10510 11947 10512
rect 10593 10507 10659 10510
rect 11881 10507 11947 10510
rect 12157 10570 12223 10573
rect 22737 10570 22803 10573
rect 12157 10568 22803 10570
rect 12157 10512 12162 10568
rect 12218 10512 22742 10568
rect 22798 10512 22803 10568
rect 12157 10510 22803 10512
rect 12157 10507 12223 10510
rect 22737 10507 22803 10510
rect 11421 10434 11487 10437
rect 12157 10434 12223 10437
rect 11421 10432 12223 10434
rect 11421 10376 11426 10432
rect 11482 10376 12162 10432
rect 12218 10376 12223 10432
rect 11421 10374 12223 10376
rect 11421 10371 11487 10374
rect 12157 10371 12223 10374
rect 12341 10434 12407 10437
rect 15469 10434 15535 10437
rect 12341 10432 15535 10434
rect 12341 10376 12346 10432
rect 12402 10376 15474 10432
rect 15530 10376 15535 10432
rect 12341 10374 15535 10376
rect 12341 10371 12407 10374
rect 15469 10371 15535 10374
rect 18505 10434 18571 10437
rect 18781 10434 18847 10437
rect 20161 10434 20227 10437
rect 18505 10432 20227 10434
rect 18505 10376 18510 10432
rect 18566 10376 18786 10432
rect 18842 10376 20166 10432
rect 20222 10376 20227 10432
rect 18505 10374 20227 10376
rect 18505 10371 18571 10374
rect 18781 10371 18847 10374
rect 20161 10371 20227 10374
rect 4210 10368 4526 10369
rect 200 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 3785 10298 3851 10301
rect 200 10296 3851 10298
rect 200 10240 3790 10296
rect 3846 10240 3851 10296
rect 200 10238 3851 10240
rect 200 10208 800 10238
rect 3785 10235 3851 10238
rect 16389 10298 16455 10301
rect 18413 10298 18479 10301
rect 16389 10296 18479 10298
rect 16389 10240 16394 10296
rect 16450 10240 18418 10296
rect 18474 10240 18479 10296
rect 16389 10238 18479 10240
rect 16389 10235 16455 10238
rect 18413 10235 18479 10238
rect 15009 10162 15075 10165
rect 23565 10162 23631 10165
rect 15009 10160 23631 10162
rect 15009 10104 15014 10160
rect 15070 10104 23570 10160
rect 23626 10104 23631 10160
rect 15009 10102 23631 10104
rect 15009 10099 15075 10102
rect 23565 10099 23631 10102
rect 12433 10026 12499 10029
rect 15837 10026 15903 10029
rect 12433 10024 15903 10026
rect 12433 9968 12438 10024
rect 12494 9968 15842 10024
rect 15898 9968 15903 10024
rect 12433 9966 15903 9968
rect 12433 9963 12499 9966
rect 15837 9963 15903 9966
rect 16573 10026 16639 10029
rect 23841 10026 23907 10029
rect 16573 10024 23907 10026
rect 16573 9968 16578 10024
rect 16634 9968 23846 10024
rect 23902 9968 23907 10024
rect 16573 9966 23907 9968
rect 16573 9963 16639 9966
rect 23841 9963 23907 9966
rect 4521 9890 4587 9893
rect 5533 9890 5599 9893
rect 4521 9888 5599 9890
rect 4521 9832 4526 9888
rect 4582 9832 5538 9888
rect 5594 9832 5599 9888
rect 4521 9830 5599 9832
rect 4521 9827 4587 9830
rect 5533 9827 5599 9830
rect 11697 9890 11763 9893
rect 12341 9890 12407 9893
rect 14917 9890 14983 9893
rect 18413 9890 18479 9893
rect 11697 9888 18479 9890
rect 11697 9832 11702 9888
rect 11758 9832 12346 9888
rect 12402 9832 14922 9888
rect 14978 9832 18418 9888
rect 18474 9832 18479 9888
rect 11697 9830 18479 9832
rect 11697 9827 11763 9830
rect 12341 9827 12407 9830
rect 14917 9827 14983 9830
rect 18413 9827 18479 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 13997 9754 14063 9757
rect 15193 9754 15259 9757
rect 13997 9752 15259 9754
rect 13997 9696 14002 9752
rect 14058 9696 15198 9752
rect 15254 9696 15259 9752
rect 13997 9694 15259 9696
rect 13997 9691 14063 9694
rect 15193 9691 15259 9694
rect 20805 9754 20871 9757
rect 20805 9752 20914 9754
rect 20805 9696 20810 9752
rect 20866 9696 20914 9752
rect 20805 9691 20914 9696
rect 16297 9618 16363 9621
rect 16430 9618 16436 9620
rect 16297 9616 16436 9618
rect 16297 9560 16302 9616
rect 16358 9560 16436 9616
rect 16297 9558 16436 9560
rect 16297 9555 16363 9558
rect 16430 9556 16436 9558
rect 16500 9556 16506 9620
rect 3417 9482 3483 9485
rect 9581 9482 9647 9485
rect 3417 9480 9647 9482
rect 3417 9424 3422 9480
rect 3478 9424 9586 9480
rect 9642 9424 9647 9480
rect 3417 9422 9647 9424
rect 3417 9419 3483 9422
rect 9581 9419 9647 9422
rect 10961 9482 11027 9485
rect 11421 9482 11487 9485
rect 20854 9482 20914 9691
rect 38193 9618 38259 9621
rect 39200 9618 39800 9648
rect 38193 9616 39800 9618
rect 38193 9560 38198 9616
rect 38254 9560 39800 9616
rect 38193 9558 39800 9560
rect 38193 9555 38259 9558
rect 39200 9528 39800 9558
rect 22645 9482 22711 9485
rect 10961 9480 22711 9482
rect 10961 9424 10966 9480
rect 11022 9424 11426 9480
rect 11482 9424 22650 9480
rect 22706 9424 22711 9480
rect 10961 9422 22711 9424
rect 10961 9419 11027 9422
rect 11421 9419 11487 9422
rect 22645 9419 22711 9422
rect 14917 9346 14983 9349
rect 20161 9346 20227 9349
rect 14917 9344 20227 9346
rect 14917 9288 14922 9344
rect 14978 9288 20166 9344
rect 20222 9288 20227 9344
rect 14917 9286 20227 9288
rect 14917 9283 14983 9286
rect 20161 9283 20227 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 13721 9074 13787 9077
rect 17033 9074 17099 9077
rect 13721 9072 17099 9074
rect 13721 9016 13726 9072
rect 13782 9016 17038 9072
rect 17094 9016 17099 9072
rect 13721 9014 17099 9016
rect 13721 9011 13787 9014
rect 17033 9011 17099 9014
rect 17677 9074 17743 9077
rect 19057 9074 19123 9077
rect 17677 9072 19123 9074
rect 17677 9016 17682 9072
rect 17738 9016 19062 9072
rect 19118 9016 19123 9072
rect 17677 9014 19123 9016
rect 17677 9011 17743 9014
rect 19057 9011 19123 9014
rect 200 8938 800 8968
rect 3969 8938 4035 8941
rect 200 8936 4035 8938
rect 200 8880 3974 8936
rect 4030 8880 4035 8936
rect 200 8878 4035 8880
rect 200 8848 800 8878
rect 3969 8875 4035 8878
rect 9949 8938 10015 8941
rect 22737 8938 22803 8941
rect 9949 8936 22803 8938
rect 9949 8880 9954 8936
rect 10010 8880 22742 8936
rect 22798 8880 22803 8936
rect 9949 8878 22803 8880
rect 9949 8875 10015 8878
rect 22737 8875 22803 8878
rect 14825 8802 14891 8805
rect 15745 8802 15811 8805
rect 14825 8800 15811 8802
rect 14825 8744 14830 8800
rect 14886 8744 15750 8800
rect 15806 8744 15811 8800
rect 14825 8742 15811 8744
rect 14825 8739 14891 8742
rect 15745 8739 15811 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 1577 8666 1643 8669
rect 7097 8668 7163 8669
rect 1710 8666 1716 8668
rect 1577 8664 1716 8666
rect 1577 8608 1582 8664
rect 1638 8608 1716 8664
rect 1577 8606 1716 8608
rect 1577 8603 1643 8606
rect 1710 8604 1716 8606
rect 1780 8604 1786 8668
rect 7046 8604 7052 8668
rect 7116 8666 7163 8668
rect 7116 8664 7208 8666
rect 7158 8608 7208 8664
rect 7116 8606 7208 8608
rect 7116 8604 7163 8606
rect 7097 8603 7163 8604
rect 13629 8530 13695 8533
rect 15469 8530 15535 8533
rect 13629 8528 15535 8530
rect 13629 8472 13634 8528
rect 13690 8472 15474 8528
rect 15530 8472 15535 8528
rect 13629 8470 15535 8472
rect 13629 8467 13695 8470
rect 15469 8467 15535 8470
rect 17125 8530 17191 8533
rect 23381 8530 23447 8533
rect 17125 8528 23447 8530
rect 17125 8472 17130 8528
rect 17186 8472 23386 8528
rect 23442 8472 23447 8528
rect 17125 8470 23447 8472
rect 17125 8467 17191 8470
rect 23381 8467 23447 8470
rect 17217 8394 17283 8397
rect 24577 8394 24643 8397
rect 17217 8392 24643 8394
rect 17217 8336 17222 8392
rect 17278 8336 24582 8392
rect 24638 8336 24643 8392
rect 17217 8334 24643 8336
rect 17217 8331 17283 8334
rect 24577 8331 24643 8334
rect 15101 8258 15167 8261
rect 21725 8258 21791 8261
rect 15101 8256 21791 8258
rect 15101 8200 15106 8256
rect 15162 8200 21730 8256
rect 21786 8200 21791 8256
rect 15101 8198 21791 8200
rect 15101 8195 15167 8198
rect 21725 8195 21791 8198
rect 38101 8258 38167 8261
rect 39200 8258 39800 8288
rect 38101 8256 39800 8258
rect 38101 8200 38106 8256
rect 38162 8200 39800 8256
rect 38101 8198 39800 8200
rect 38101 8195 38167 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 39200 8168 39800 8198
rect 34930 8127 35246 8128
rect 790 8060 796 8124
rect 860 8122 866 8124
rect 3417 8122 3483 8125
rect 860 8120 3483 8122
rect 860 8064 3422 8120
rect 3478 8064 3483 8120
rect 860 8062 3483 8064
rect 860 8060 866 8062
rect 3417 8059 3483 8062
rect 19241 8122 19307 8125
rect 22461 8122 22527 8125
rect 22645 8122 22711 8125
rect 19241 8120 22711 8122
rect 19241 8064 19246 8120
rect 19302 8064 22466 8120
rect 22522 8064 22650 8120
rect 22706 8064 22711 8120
rect 19241 8062 22711 8064
rect 19241 8059 19307 8062
rect 22461 8059 22527 8062
rect 22645 8059 22711 8062
rect 18229 7986 18295 7989
rect 26233 7986 26299 7989
rect 18229 7984 26299 7986
rect 18229 7928 18234 7984
rect 18290 7928 26238 7984
rect 26294 7928 26299 7984
rect 18229 7926 26299 7928
rect 18229 7923 18295 7926
rect 26233 7923 26299 7926
rect 16665 7850 16731 7853
rect 25313 7850 25379 7853
rect 16665 7848 25379 7850
rect 16665 7792 16670 7848
rect 16726 7792 25318 7848
rect 25374 7792 25379 7848
rect 16665 7790 25379 7792
rect 16665 7787 16731 7790
rect 25313 7787 25379 7790
rect 14825 7714 14891 7717
rect 19149 7714 19215 7717
rect 14825 7712 19215 7714
rect 14825 7656 14830 7712
rect 14886 7656 19154 7712
rect 19210 7656 19215 7712
rect 14825 7654 19215 7656
rect 14825 7651 14891 7654
rect 19149 7651 19215 7654
rect 19570 7648 19886 7649
rect 200 7578 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 1393 7578 1459 7581
rect 200 7576 1459 7578
rect 200 7520 1398 7576
rect 1454 7520 1459 7576
rect 200 7518 1459 7520
rect 200 7488 800 7518
rect 1393 7515 1459 7518
rect 9857 7578 9923 7581
rect 19241 7578 19307 7581
rect 9857 7576 19307 7578
rect 9857 7520 9862 7576
rect 9918 7520 19246 7576
rect 19302 7520 19307 7576
rect 9857 7518 19307 7520
rect 9857 7515 9923 7518
rect 19241 7515 19307 7518
rect 37457 7578 37523 7581
rect 39200 7578 39800 7608
rect 37457 7576 39800 7578
rect 37457 7520 37462 7576
rect 37518 7520 39800 7576
rect 37457 7518 39800 7520
rect 37457 7515 37523 7518
rect 39200 7488 39800 7518
rect 10961 7442 11027 7445
rect 21449 7442 21515 7445
rect 10961 7440 21515 7442
rect 10961 7384 10966 7440
rect 11022 7384 21454 7440
rect 21510 7384 21515 7440
rect 10961 7382 21515 7384
rect 10961 7379 11027 7382
rect 21449 7379 21515 7382
rect 1853 7306 1919 7309
rect 17902 7306 17908 7308
rect 1853 7304 17908 7306
rect 1853 7248 1858 7304
rect 1914 7248 17908 7304
rect 1853 7246 17908 7248
rect 1853 7243 1919 7246
rect 17902 7244 17908 7246
rect 17972 7244 17978 7308
rect 10777 7170 10843 7173
rect 18873 7170 18939 7173
rect 10777 7168 18939 7170
rect 10777 7112 10782 7168
rect 10838 7112 18878 7168
rect 18934 7112 18939 7168
rect 10777 7110 18939 7112
rect 10777 7107 10843 7110
rect 18873 7107 18939 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 9673 7034 9739 7037
rect 11145 7034 11211 7037
rect 9673 7032 11211 7034
rect 9673 6976 9678 7032
rect 9734 6976 11150 7032
rect 11206 6976 11211 7032
rect 9673 6974 11211 6976
rect 9673 6971 9739 6974
rect 11145 6971 11211 6974
rect 13445 7034 13511 7037
rect 21173 7034 21239 7037
rect 13445 7032 21239 7034
rect 13445 6976 13450 7032
rect 13506 6976 21178 7032
rect 21234 6976 21239 7032
rect 13445 6974 21239 6976
rect 13445 6971 13511 6974
rect 21173 6971 21239 6974
rect 200 6898 800 6928
rect 1761 6898 1827 6901
rect 200 6896 1827 6898
rect 200 6840 1766 6896
rect 1822 6840 1827 6896
rect 200 6838 1827 6840
rect 200 6808 800 6838
rect 1761 6835 1827 6838
rect 9673 6898 9739 6901
rect 10501 6898 10567 6901
rect 9673 6896 10567 6898
rect 9673 6840 9678 6896
rect 9734 6840 10506 6896
rect 10562 6840 10567 6896
rect 9673 6838 10567 6840
rect 9673 6835 9739 6838
rect 10501 6835 10567 6838
rect 13169 6898 13235 6901
rect 15285 6898 15351 6901
rect 17769 6900 17835 6901
rect 17718 6898 17724 6900
rect 13169 6896 15351 6898
rect 13169 6840 13174 6896
rect 13230 6840 15290 6896
rect 15346 6840 15351 6896
rect 13169 6838 15351 6840
rect 17678 6838 17724 6898
rect 17788 6896 17835 6900
rect 17830 6840 17835 6896
rect 13169 6835 13235 6838
rect 15285 6835 15351 6838
rect 17718 6836 17724 6838
rect 17788 6836 17835 6840
rect 17769 6835 17835 6836
rect 18045 6898 18111 6901
rect 21357 6898 21423 6901
rect 18045 6896 21423 6898
rect 18045 6840 18050 6896
rect 18106 6840 21362 6896
rect 21418 6840 21423 6896
rect 18045 6838 21423 6840
rect 18045 6835 18111 6838
rect 21357 6835 21423 6838
rect 7649 6762 7715 6765
rect 15653 6762 15719 6765
rect 7649 6760 15719 6762
rect 7649 6704 7654 6760
rect 7710 6704 15658 6760
rect 15714 6704 15719 6760
rect 7649 6702 15719 6704
rect 7649 6699 7715 6702
rect 15653 6699 15719 6702
rect 15837 6762 15903 6765
rect 23289 6762 23355 6765
rect 15837 6760 23355 6762
rect 15837 6704 15842 6760
rect 15898 6704 23294 6760
rect 23350 6704 23355 6760
rect 15837 6702 23355 6704
rect 15837 6699 15903 6702
rect 23289 6699 23355 6702
rect 12249 6626 12315 6629
rect 14406 6626 14412 6628
rect 12249 6624 14412 6626
rect 12249 6568 12254 6624
rect 12310 6568 14412 6624
rect 12249 6566 14412 6568
rect 12249 6563 12315 6566
rect 14406 6564 14412 6566
rect 14476 6626 14482 6628
rect 18045 6626 18111 6629
rect 14476 6624 18111 6626
rect 14476 6568 18050 6624
rect 18106 6568 18111 6624
rect 14476 6566 18111 6568
rect 14476 6564 14482 6566
rect 18045 6563 18111 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 16849 6490 16915 6493
rect 18045 6490 18111 6493
rect 16849 6488 18111 6490
rect 16849 6432 16854 6488
rect 16910 6432 18050 6488
rect 18106 6432 18111 6488
rect 16849 6430 18111 6432
rect 16849 6427 16915 6430
rect 18045 6427 18111 6430
rect 15653 6354 15719 6357
rect 20713 6354 20779 6357
rect 15653 6352 20779 6354
rect 15653 6296 15658 6352
rect 15714 6296 20718 6352
rect 20774 6296 20779 6352
rect 15653 6294 20779 6296
rect 15653 6291 15719 6294
rect 20713 6291 20779 6294
rect 16481 6218 16547 6221
rect 30649 6218 30715 6221
rect 16481 6216 30715 6218
rect 16481 6160 16486 6216
rect 16542 6160 30654 6216
rect 30710 6160 30715 6216
rect 16481 6158 30715 6160
rect 16481 6155 16547 6158
rect 30649 6155 30715 6158
rect 38285 6218 38351 6221
rect 39200 6218 39800 6248
rect 38285 6216 39800 6218
rect 38285 6160 38290 6216
rect 38346 6160 39800 6216
rect 38285 6158 39800 6160
rect 38285 6155 38351 6158
rect 39200 6128 39800 6158
rect 15653 6082 15719 6085
rect 22829 6082 22895 6085
rect 15653 6080 22895 6082
rect 15653 6024 15658 6080
rect 15714 6024 22834 6080
rect 22890 6024 22895 6080
rect 15653 6022 22895 6024
rect 15653 6019 15719 6022
rect 22829 6019 22895 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 8661 5946 8727 5949
rect 23289 5946 23355 5949
rect 8661 5944 23355 5946
rect 8661 5888 8666 5944
rect 8722 5888 23294 5944
rect 23350 5888 23355 5944
rect 8661 5886 23355 5888
rect 8661 5883 8727 5886
rect 23289 5883 23355 5886
rect 4061 5810 4127 5813
rect 18045 5810 18111 5813
rect 4061 5808 18111 5810
rect 4061 5752 4066 5808
rect 4122 5752 18050 5808
rect 18106 5752 18111 5808
rect 4061 5750 18111 5752
rect 4061 5747 4127 5750
rect 18045 5747 18111 5750
rect 18689 5810 18755 5813
rect 21817 5810 21883 5813
rect 18689 5808 21883 5810
rect 18689 5752 18694 5808
rect 18750 5752 21822 5808
rect 21878 5752 21883 5808
rect 18689 5750 21883 5752
rect 18689 5747 18755 5750
rect 21817 5747 21883 5750
rect 8385 5674 8451 5677
rect 12617 5674 12683 5677
rect 8385 5672 12683 5674
rect 8385 5616 8390 5672
rect 8446 5616 12622 5672
rect 12678 5616 12683 5672
rect 8385 5614 12683 5616
rect 8385 5611 8451 5614
rect 12617 5611 12683 5614
rect 17401 5674 17467 5677
rect 17861 5674 17927 5677
rect 20897 5674 20963 5677
rect 17401 5672 20963 5674
rect 17401 5616 17406 5672
rect 17462 5616 17866 5672
rect 17922 5616 20902 5672
rect 20958 5616 20963 5672
rect 17401 5614 20963 5616
rect 17401 5611 17467 5614
rect 17861 5611 17927 5614
rect 20897 5611 20963 5614
rect 200 5538 800 5568
rect 1393 5538 1459 5541
rect 200 5536 1459 5538
rect 200 5480 1398 5536
rect 1454 5480 1459 5536
rect 200 5478 1459 5480
rect 200 5448 800 5478
rect 1393 5475 1459 5478
rect 17861 5538 17927 5541
rect 19333 5538 19399 5541
rect 17861 5536 19399 5538
rect 17861 5480 17866 5536
rect 17922 5480 19338 5536
rect 19394 5480 19399 5536
rect 17861 5478 19399 5480
rect 17861 5475 17927 5478
rect 19333 5475 19399 5478
rect 20069 5538 20135 5541
rect 20529 5538 20595 5541
rect 20069 5536 20595 5538
rect 20069 5480 20074 5536
rect 20130 5480 20534 5536
rect 20590 5480 20595 5536
rect 20069 5478 20595 5480
rect 20069 5475 20135 5478
rect 20529 5475 20595 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 9029 5402 9095 5405
rect 11605 5402 11671 5405
rect 9029 5400 11671 5402
rect 9029 5344 9034 5400
rect 9090 5344 11610 5400
rect 11666 5344 11671 5400
rect 9029 5342 11671 5344
rect 9029 5339 9095 5342
rect 11605 5339 11671 5342
rect 13905 5402 13971 5405
rect 18137 5402 18203 5405
rect 13905 5400 18203 5402
rect 13905 5344 13910 5400
rect 13966 5344 18142 5400
rect 18198 5344 18203 5400
rect 13905 5342 18203 5344
rect 13905 5339 13971 5342
rect 18137 5339 18203 5342
rect 19977 5402 20043 5405
rect 20253 5402 20319 5405
rect 19977 5400 20319 5402
rect 19977 5344 19982 5400
rect 20038 5344 20258 5400
rect 20314 5344 20319 5400
rect 19977 5342 20319 5344
rect 19977 5339 20043 5342
rect 20253 5339 20319 5342
rect 20621 5402 20687 5405
rect 21173 5402 21239 5405
rect 20621 5400 21239 5402
rect 20621 5344 20626 5400
rect 20682 5344 21178 5400
rect 21234 5344 21239 5400
rect 20621 5342 21239 5344
rect 20621 5339 20687 5342
rect 21173 5339 21239 5342
rect 6913 5266 6979 5269
rect 21081 5266 21147 5269
rect 6913 5264 21147 5266
rect 6913 5208 6918 5264
rect 6974 5208 21086 5264
rect 21142 5208 21147 5264
rect 6913 5206 21147 5208
rect 6913 5203 6979 5206
rect 21081 5203 21147 5206
rect 15745 5130 15811 5133
rect 17585 5130 17651 5133
rect 15745 5128 17651 5130
rect 15745 5072 15750 5128
rect 15806 5072 17590 5128
rect 17646 5072 17651 5128
rect 15745 5070 17651 5072
rect 15745 5067 15811 5070
rect 17585 5067 17651 5070
rect 18045 5130 18111 5133
rect 23749 5130 23815 5133
rect 18045 5128 23815 5130
rect 18045 5072 18050 5128
rect 18106 5072 23754 5128
rect 23810 5072 23815 5128
rect 18045 5070 23815 5072
rect 18045 5067 18111 5070
rect 23749 5067 23815 5070
rect 13261 4994 13327 4997
rect 22001 4994 22067 4997
rect 13261 4992 22067 4994
rect 13261 4936 13266 4992
rect 13322 4936 22006 4992
rect 22062 4936 22067 4992
rect 13261 4934 22067 4936
rect 13261 4931 13327 4934
rect 22001 4931 22067 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 9305 4858 9371 4861
rect 20529 4858 20595 4861
rect 9305 4856 20595 4858
rect 9305 4800 9310 4856
rect 9366 4800 20534 4856
rect 20590 4800 20595 4856
rect 9305 4798 20595 4800
rect 9305 4795 9371 4798
rect 20529 4795 20595 4798
rect 38193 4858 38259 4861
rect 39200 4858 39800 4888
rect 38193 4856 39800 4858
rect 38193 4800 38198 4856
rect 38254 4800 39800 4856
rect 38193 4798 39800 4800
rect 38193 4795 38259 4798
rect 39200 4768 39800 4798
rect 7741 4722 7807 4725
rect 13813 4722 13879 4725
rect 7741 4720 13879 4722
rect 7741 4664 7746 4720
rect 7802 4664 13818 4720
rect 13874 4664 13879 4720
rect 7741 4662 13879 4664
rect 7741 4659 7807 4662
rect 13813 4659 13879 4662
rect 15837 4722 15903 4725
rect 20713 4722 20779 4725
rect 15837 4720 20779 4722
rect 15837 4664 15842 4720
rect 15898 4664 20718 4720
rect 20774 4664 20779 4720
rect 15837 4662 20779 4664
rect 15837 4659 15903 4662
rect 20713 4659 20779 4662
rect 7925 4586 7991 4589
rect 24669 4586 24735 4589
rect 7925 4584 24735 4586
rect 7925 4528 7930 4584
rect 7986 4528 24674 4584
rect 24730 4528 24735 4584
rect 7925 4526 24735 4528
rect 7925 4523 7991 4526
rect 24669 4523 24735 4526
rect 8109 4450 8175 4453
rect 19241 4450 19307 4453
rect 8109 4448 19307 4450
rect 8109 4392 8114 4448
rect 8170 4392 19246 4448
rect 19302 4392 19307 4448
rect 8109 4390 19307 4392
rect 8109 4387 8175 4390
rect 19241 4387 19307 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 13813 4314 13879 4317
rect 15101 4314 15167 4317
rect 13813 4312 15167 4314
rect 13813 4256 13818 4312
rect 13874 4256 15106 4312
rect 15162 4256 15167 4312
rect 13813 4254 15167 4256
rect 13813 4251 13879 4254
rect 15101 4251 15167 4254
rect 16021 4314 16087 4317
rect 18689 4314 18755 4317
rect 16021 4312 18755 4314
rect 16021 4256 16026 4312
rect 16082 4256 18694 4312
rect 18750 4256 18755 4312
rect 16021 4254 18755 4256
rect 16021 4251 16087 4254
rect 18689 4251 18755 4254
rect 19333 4316 19399 4317
rect 19333 4312 19380 4316
rect 19444 4314 19450 4316
rect 19977 4314 20043 4317
rect 21909 4314 21975 4317
rect 19333 4256 19338 4312
rect 19333 4252 19380 4256
rect 19444 4254 19490 4314
rect 19977 4312 21975 4314
rect 19977 4256 19982 4312
rect 20038 4256 21914 4312
rect 21970 4256 21975 4312
rect 19977 4254 21975 4256
rect 19444 4252 19450 4254
rect 19333 4251 19399 4252
rect 19977 4251 20043 4254
rect 21909 4251 21975 4254
rect 200 4178 800 4208
rect 1669 4178 1735 4181
rect 200 4176 1735 4178
rect 200 4120 1674 4176
rect 1730 4120 1735 4176
rect 200 4118 1735 4120
rect 200 4088 800 4118
rect 1669 4115 1735 4118
rect 9581 4178 9647 4181
rect 24577 4178 24643 4181
rect 9581 4176 24643 4178
rect 9581 4120 9586 4176
rect 9642 4120 24582 4176
rect 24638 4120 24643 4176
rect 9581 4118 24643 4120
rect 9581 4115 9647 4118
rect 24577 4115 24643 4118
rect 38285 4178 38351 4181
rect 39200 4178 39800 4208
rect 38285 4176 39800 4178
rect 38285 4120 38290 4176
rect 38346 4120 39800 4176
rect 38285 4118 39800 4120
rect 38285 4115 38351 4118
rect 39200 4088 39800 4118
rect 8937 4042 9003 4045
rect 12065 4042 12131 4045
rect 8937 4040 12131 4042
rect 8937 3984 8942 4040
rect 8998 3984 12070 4040
rect 12126 3984 12131 4040
rect 8937 3982 12131 3984
rect 8937 3979 9003 3982
rect 12065 3979 12131 3982
rect 13537 4042 13603 4045
rect 21541 4042 21607 4045
rect 13537 4040 21607 4042
rect 13537 3984 13542 4040
rect 13598 3984 21546 4040
rect 21602 3984 21607 4040
rect 13537 3982 21607 3984
rect 13537 3979 13603 3982
rect 21541 3979 21607 3982
rect 11329 3906 11395 3909
rect 12985 3906 13051 3909
rect 11329 3904 13051 3906
rect 11329 3848 11334 3904
rect 11390 3848 12990 3904
rect 13046 3848 13051 3904
rect 11329 3846 13051 3848
rect 11329 3843 11395 3846
rect 12985 3843 13051 3846
rect 15285 3906 15351 3909
rect 23381 3906 23447 3909
rect 15285 3904 23447 3906
rect 15285 3848 15290 3904
rect 15346 3848 23386 3904
rect 23442 3848 23447 3904
rect 15285 3846 23447 3848
rect 15285 3843 15351 3846
rect 23381 3843 23447 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 9397 3770 9463 3773
rect 12249 3770 12315 3773
rect 9397 3768 12315 3770
rect 9397 3712 9402 3768
rect 9458 3712 12254 3768
rect 12310 3712 12315 3768
rect 9397 3710 12315 3712
rect 9397 3707 9463 3710
rect 12249 3707 12315 3710
rect 16573 3770 16639 3773
rect 17217 3770 17283 3773
rect 16573 3768 17283 3770
rect 16573 3712 16578 3768
rect 16634 3712 17222 3768
rect 17278 3712 17283 3768
rect 16573 3710 17283 3712
rect 16573 3707 16639 3710
rect 17217 3707 17283 3710
rect 19333 3770 19399 3773
rect 21173 3770 21239 3773
rect 19333 3768 21239 3770
rect 19333 3712 19338 3768
rect 19394 3712 21178 3768
rect 21234 3712 21239 3768
rect 19333 3710 21239 3712
rect 19333 3707 19399 3710
rect 21173 3707 21239 3710
rect 6637 3634 6703 3637
rect 8385 3634 8451 3637
rect 12157 3634 12223 3637
rect 6637 3632 12223 3634
rect 6637 3576 6642 3632
rect 6698 3576 8390 3632
rect 8446 3576 12162 3632
rect 12218 3576 12223 3632
rect 6637 3574 12223 3576
rect 6637 3571 6703 3574
rect 8385 3571 8451 3574
rect 12157 3571 12223 3574
rect 16389 3634 16455 3637
rect 23381 3634 23447 3637
rect 16389 3632 23447 3634
rect 16389 3576 16394 3632
rect 16450 3576 23386 3632
rect 23442 3576 23447 3632
rect 16389 3574 23447 3576
rect 16389 3571 16455 3574
rect 23381 3571 23447 3574
rect 200 3498 800 3528
rect 4061 3498 4127 3501
rect 200 3496 4127 3498
rect 200 3440 4066 3496
rect 4122 3440 4127 3496
rect 200 3438 4127 3440
rect 200 3408 800 3438
rect 4061 3435 4127 3438
rect 7557 3498 7623 3501
rect 17769 3498 17835 3501
rect 18873 3498 18939 3501
rect 7557 3496 17648 3498
rect 7557 3440 7562 3496
rect 7618 3440 17648 3496
rect 7557 3438 17648 3440
rect 7557 3435 7623 3438
rect 3141 3362 3207 3365
rect 6085 3362 6151 3365
rect 3141 3360 6151 3362
rect 3141 3304 3146 3360
rect 3202 3304 6090 3360
rect 6146 3304 6151 3360
rect 3141 3302 6151 3304
rect 3141 3299 3207 3302
rect 6085 3299 6151 3302
rect 13629 3362 13695 3365
rect 16297 3362 16363 3365
rect 13629 3360 16363 3362
rect 13629 3304 13634 3360
rect 13690 3304 16302 3360
rect 16358 3304 16363 3360
rect 13629 3302 16363 3304
rect 13629 3299 13695 3302
rect 16297 3299 16363 3302
rect 16757 3362 16823 3365
rect 17309 3362 17375 3365
rect 16757 3360 17375 3362
rect 16757 3304 16762 3360
rect 16818 3304 17314 3360
rect 17370 3304 17375 3360
rect 16757 3302 17375 3304
rect 17588 3362 17648 3438
rect 17769 3496 18939 3498
rect 17769 3440 17774 3496
rect 17830 3440 18878 3496
rect 18934 3440 18939 3496
rect 17769 3438 18939 3440
rect 17769 3435 17835 3438
rect 18873 3435 18939 3438
rect 19374 3436 19380 3500
rect 19444 3498 19450 3500
rect 22737 3498 22803 3501
rect 19444 3496 22803 3498
rect 19444 3440 22742 3496
rect 22798 3440 22803 3496
rect 19444 3438 22803 3440
rect 19444 3436 19450 3438
rect 22737 3435 22803 3438
rect 18045 3362 18111 3365
rect 17588 3360 18111 3362
rect 17588 3304 18050 3360
rect 18106 3304 18111 3360
rect 17588 3302 18111 3304
rect 16757 3299 16823 3302
rect 17309 3299 17375 3302
rect 18045 3299 18111 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 16665 3226 16731 3229
rect 19241 3226 19307 3229
rect 16665 3224 19307 3226
rect 16665 3168 16670 3224
rect 16726 3168 19246 3224
rect 19302 3168 19307 3224
rect 16665 3166 19307 3168
rect 16665 3163 16731 3166
rect 19241 3163 19307 3166
rect 4337 3090 4403 3093
rect 7281 3090 7347 3093
rect 4337 3088 7347 3090
rect 4337 3032 4342 3088
rect 4398 3032 7286 3088
rect 7342 3032 7347 3088
rect 4337 3030 7347 3032
rect 4337 3027 4403 3030
rect 7281 3027 7347 3030
rect 14825 3090 14891 3093
rect 17953 3090 18019 3093
rect 14825 3088 18019 3090
rect 14825 3032 14830 3088
rect 14886 3032 17958 3088
rect 18014 3032 18019 3088
rect 14825 3030 18019 3032
rect 14825 3027 14891 3030
rect 17953 3027 18019 3030
rect 18137 3090 18203 3093
rect 18965 3090 19031 3093
rect 22553 3090 22619 3093
rect 18137 3088 22619 3090
rect 18137 3032 18142 3088
rect 18198 3032 18970 3088
rect 19026 3032 22558 3088
rect 22614 3032 22619 3088
rect 18137 3030 22619 3032
rect 18137 3027 18203 3030
rect 18965 3027 19031 3030
rect 22553 3027 22619 3030
rect 4061 2954 4127 2957
rect 20069 2954 20135 2957
rect 4061 2952 20135 2954
rect 4061 2896 4066 2952
rect 4122 2896 20074 2952
rect 20130 2896 20135 2952
rect 4061 2894 20135 2896
rect 4061 2891 4127 2894
rect 20069 2891 20135 2894
rect 5533 2818 5599 2821
rect 14181 2818 14247 2821
rect 5533 2816 14247 2818
rect 5533 2760 5538 2816
rect 5594 2760 14186 2816
rect 14242 2760 14247 2816
rect 5533 2758 14247 2760
rect 5533 2755 5599 2758
rect 14181 2755 14247 2758
rect 15469 2818 15535 2821
rect 24025 2818 24091 2821
rect 15469 2816 24091 2818
rect 15469 2760 15474 2816
rect 15530 2760 24030 2816
rect 24086 2760 24091 2816
rect 15469 2758 24091 2760
rect 15469 2755 15535 2758
rect 24025 2755 24091 2758
rect 38285 2818 38351 2821
rect 39200 2818 39800 2848
rect 38285 2816 39800 2818
rect 38285 2760 38290 2816
rect 38346 2760 39800 2816
rect 38285 2758 39800 2760
rect 38285 2755 38351 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 39200 2728 39800 2758
rect 34930 2687 35246 2688
rect 5257 2682 5323 2685
rect 10869 2684 10935 2685
rect 13445 2684 13511 2685
rect 7414 2682 7420 2684
rect 5257 2680 7420 2682
rect 5257 2624 5262 2680
rect 5318 2624 7420 2680
rect 5257 2622 7420 2624
rect 5257 2619 5323 2622
rect 7414 2620 7420 2622
rect 7484 2620 7490 2684
rect 10869 2680 10916 2684
rect 10980 2682 10986 2684
rect 10869 2624 10874 2680
rect 10869 2620 10916 2624
rect 10980 2622 11026 2682
rect 13445 2680 13492 2684
rect 13556 2682 13562 2684
rect 13445 2624 13450 2680
rect 10980 2620 10986 2622
rect 13445 2620 13492 2624
rect 13556 2622 13602 2682
rect 13556 2620 13562 2622
rect 10869 2619 10935 2620
rect 13445 2619 13511 2620
rect 10501 2546 10567 2549
rect 23381 2546 23447 2549
rect 10501 2544 23447 2546
rect 10501 2488 10506 2544
rect 10562 2488 23386 2544
rect 23442 2488 23447 2544
rect 10501 2486 23447 2488
rect 10501 2483 10567 2486
rect 23381 2483 23447 2486
rect 10961 2410 11027 2413
rect 27153 2410 27219 2413
rect 10961 2408 27219 2410
rect 10961 2352 10966 2408
rect 11022 2352 27158 2408
rect 27214 2352 27219 2408
rect 10961 2350 27219 2352
rect 10961 2347 11027 2350
rect 27153 2347 27219 2350
rect 19570 2208 19886 2209
rect 200 2138 800 2168
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 2497 2138 2563 2141
rect 200 2136 2563 2138
rect 200 2080 2502 2136
rect 2558 2080 2563 2136
rect 200 2078 2563 2080
rect 200 2048 800 2078
rect 2497 2075 2563 2078
rect 2681 2002 2747 2005
rect 26049 2002 26115 2005
rect 2681 2000 26115 2002
rect 2681 1944 2686 2000
rect 2742 1944 26054 2000
rect 26110 1944 26115 2000
rect 2681 1942 26115 1944
rect 2681 1939 2747 1942
rect 26049 1939 26115 1942
rect 2865 1866 2931 1869
rect 23565 1866 23631 1869
rect 2865 1864 23631 1866
rect 2865 1808 2870 1864
rect 2926 1808 23570 1864
rect 23626 1808 23631 1864
rect 2865 1806 23631 1808
rect 2865 1803 2931 1806
rect 23565 1803 23631 1806
rect 10409 1730 10475 1733
rect 22093 1730 22159 1733
rect 10409 1728 22159 1730
rect 10409 1672 10414 1728
rect 10470 1672 22098 1728
rect 22154 1672 22159 1728
rect 10409 1670 22159 1672
rect 10409 1667 10475 1670
rect 22093 1667 22159 1670
rect 36905 1458 36971 1461
rect 39200 1458 39800 1488
rect 36905 1456 39800 1458
rect 36905 1400 36910 1456
rect 36966 1400 39800 1456
rect 36905 1398 39800 1400
rect 36905 1395 36971 1398
rect 39200 1368 39800 1398
rect 200 778 800 808
rect 1669 778 1735 781
rect 200 776 1735 778
rect 200 720 1674 776
rect 1730 720 1735 776
rect 200 718 1735 720
rect 200 688 800 718
rect 1669 715 1735 718
rect 37641 778 37707 781
rect 39200 778 39800 808
rect 37641 776 39800 778
rect 37641 720 37646 776
rect 37702 720 39800 776
rect 37641 718 39800 720
rect 37641 715 37707 718
rect 39200 688 39800 718
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 1900 29004 1964 29068
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 12572 28052 12636 28116
rect 13124 27916 13188 27980
rect 980 27780 1044 27844
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 1716 27644 1780 27708
rect 2084 27704 2148 27708
rect 2084 27648 2098 27704
rect 2098 27648 2148 27704
rect 2084 27644 2148 27648
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 5580 26828 5644 26892
rect 3004 26692 3068 26756
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 5764 26420 5828 26484
rect 1164 26284 1228 26348
rect 4660 26344 4724 26348
rect 4660 26288 4674 26344
rect 4674 26288 4724 26344
rect 4660 26284 4724 26288
rect 10548 26284 10612 26348
rect 2820 26208 2884 26212
rect 2820 26152 2834 26208
rect 2834 26152 2884 26208
rect 2820 26148 2884 26152
rect 16620 26148 16684 26212
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 9260 25196 9324 25260
rect 7236 25120 7300 25124
rect 7236 25064 7250 25120
rect 7250 25064 7300 25120
rect 7236 25060 7300 25064
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 796 24924 860 24988
rect 3924 24984 3988 24988
rect 3924 24928 3938 24984
rect 3938 24928 3988 24984
rect 3924 24924 3988 24928
rect 4844 24924 4908 24988
rect 7052 24984 7116 24988
rect 7052 24928 7066 24984
rect 7066 24928 7116 24984
rect 7052 24924 7116 24928
rect 15516 24924 15580 24988
rect 5948 24788 6012 24852
rect 8892 24788 8956 24852
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 3556 24108 3620 24172
rect 2636 23972 2700 24036
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 3188 23428 3252 23492
rect 3740 23428 3804 23492
rect 7604 23428 7668 23492
rect 10916 23564 10980 23628
rect 11836 23564 11900 23628
rect 9996 23428 10060 23492
rect 10180 23488 10244 23492
rect 10180 23432 10230 23488
rect 10230 23432 10244 23488
rect 10180 23428 10244 23432
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 14412 23020 14476 23084
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 20116 22476 20180 22540
rect 6500 22340 6564 22404
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 11100 22204 11164 22268
rect 3740 21932 3804 21996
rect 6868 21932 6932 21996
rect 5028 21856 5092 21860
rect 5028 21800 5078 21856
rect 5078 21800 5092 21856
rect 5028 21796 5092 21800
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 11100 21524 11164 21588
rect 3924 21388 3988 21452
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 3556 20980 3620 21044
rect 4660 20768 4724 20772
rect 4660 20712 4710 20768
rect 4710 20712 4724 20768
rect 4660 20708 4724 20712
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 5948 20300 6012 20364
rect 9996 20436 10060 20500
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 5028 19620 5092 19684
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 11100 19484 11164 19548
rect 4844 19348 4908 19412
rect 6684 19408 6748 19412
rect 6684 19352 6698 19408
rect 6698 19352 6748 19408
rect 6684 19348 6748 19352
rect 1900 19272 1964 19276
rect 1900 19216 1914 19272
rect 1914 19216 1964 19272
rect 1900 19212 1964 19216
rect 2084 19272 2148 19276
rect 2084 19216 2134 19272
rect 2134 19216 2148 19272
rect 2084 19212 2148 19216
rect 3004 19212 3068 19276
rect 4660 19212 4724 19276
rect 17724 19212 17788 19276
rect 2820 19076 2884 19140
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 1164 18940 1228 19004
rect 16436 18668 16500 18732
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4660 18260 4724 18324
rect 11100 18260 11164 18324
rect 7052 18124 7116 18188
rect 13492 17988 13556 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 7604 17912 7668 17916
rect 7604 17856 7654 17912
rect 7654 17856 7668 17912
rect 7604 17852 7668 17856
rect 2636 17716 2700 17780
rect 3924 17640 3988 17644
rect 3924 17584 3974 17640
rect 3974 17584 3988 17640
rect 3924 17580 3988 17584
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 7052 17172 7116 17236
rect 12572 17172 12636 17236
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 9444 16492 9508 16556
rect 9076 16416 9140 16420
rect 9076 16360 9126 16416
rect 9126 16360 9140 16416
rect 9076 16356 9140 16360
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 7420 16084 7484 16148
rect 16436 15948 16500 16012
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 8892 15676 8956 15740
rect 9260 15676 9324 15740
rect 16620 15268 16684 15332
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 5580 15192 5644 15196
rect 5580 15136 5594 15192
rect 5594 15136 5644 15192
rect 5580 15132 5644 15136
rect 11836 14996 11900 15060
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 10548 14588 10612 14652
rect 7236 14452 7300 14516
rect 9076 14452 9140 14516
rect 4660 14180 4724 14244
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 6868 14044 6932 14108
rect 11836 13772 11900 13836
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 980 13364 1044 13428
rect 16436 13364 16500 13428
rect 10180 13228 10244 13292
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 13124 12880 13188 12884
rect 13124 12824 13138 12880
rect 13138 12824 13188 12880
rect 13124 12820 13188 12824
rect 5764 12684 5828 12748
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 13124 12472 13188 12476
rect 13124 12416 13174 12472
rect 13174 12416 13188 12472
rect 13124 12412 13188 12416
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 3188 12336 3252 12340
rect 3188 12280 3202 12336
rect 3202 12280 3252 12336
rect 3188 12276 3252 12280
rect 20116 12276 20180 12340
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 6500 11596 6564 11660
rect 6684 11520 6748 11524
rect 6684 11464 6698 11520
rect 6698 11464 6748 11520
rect 6684 11460 6748 11464
rect 15516 11596 15580 11660
rect 17908 11596 17972 11660
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 9444 10508 9508 10572
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 16436 9556 16500 9620
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 1716 8604 1780 8668
rect 7052 8664 7116 8668
rect 7052 8608 7102 8664
rect 7102 8608 7116 8664
rect 7052 8604 7116 8608
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 796 8060 860 8124
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 17908 7244 17972 7308
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 17724 6896 17788 6900
rect 17724 6840 17774 6896
rect 17774 6840 17788 6896
rect 17724 6836 17788 6840
rect 14412 6564 14476 6628
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 19380 4312 19444 4316
rect 19380 4256 19394 4312
rect 19394 4256 19444 4312
rect 19380 4252 19444 4256
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19380 3436 19444 3500
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 7420 2620 7484 2684
rect 10916 2680 10980 2684
rect 10916 2624 10930 2680
rect 10930 2624 10980 2680
rect 10916 2620 10980 2624
rect 13492 2680 13556 2684
rect 13492 2624 13506 2680
rect 13506 2624 13556 2680
rect 13492 2620 13556 2624
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 1899 29068 1965 29069
rect 1899 29004 1900 29068
rect 1964 29004 1965 29068
rect 1899 29003 1965 29004
rect 979 27844 1045 27845
rect 979 27780 980 27844
rect 1044 27780 1045 27844
rect 979 27779 1045 27780
rect 795 24988 861 24989
rect 795 24924 796 24988
rect 860 24924 861 24988
rect 795 24923 861 24924
rect 798 8125 858 24923
rect 982 13429 1042 27779
rect 1715 27708 1781 27709
rect 1715 27644 1716 27708
rect 1780 27644 1781 27708
rect 1715 27643 1781 27644
rect 1163 26348 1229 26349
rect 1163 26284 1164 26348
rect 1228 26284 1229 26348
rect 1163 26283 1229 26284
rect 1166 19005 1226 26283
rect 1163 19004 1229 19005
rect 1163 18940 1164 19004
rect 1228 18940 1229 19004
rect 1163 18939 1229 18940
rect 979 13428 1045 13429
rect 979 13364 980 13428
rect 1044 13364 1045 13428
rect 979 13363 1045 13364
rect 1718 8669 1778 27643
rect 1902 19277 1962 29003
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 12571 28116 12637 28117
rect 12571 28052 12572 28116
rect 12636 28052 12637 28116
rect 12571 28051 12637 28052
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 2083 27708 2149 27709
rect 2083 27644 2084 27708
rect 2148 27644 2149 27708
rect 2083 27643 2149 27644
rect 2086 19277 2146 27643
rect 3003 26756 3069 26757
rect 3003 26692 3004 26756
rect 3068 26692 3069 26756
rect 3003 26691 3069 26692
rect 2819 26212 2885 26213
rect 2819 26148 2820 26212
rect 2884 26148 2885 26212
rect 2819 26147 2885 26148
rect 2635 24036 2701 24037
rect 2635 23972 2636 24036
rect 2700 23972 2701 24036
rect 2635 23971 2701 23972
rect 1899 19276 1965 19277
rect 1899 19212 1900 19276
rect 1964 19212 1965 19276
rect 1899 19211 1965 19212
rect 2083 19276 2149 19277
rect 2083 19212 2084 19276
rect 2148 19212 2149 19276
rect 2083 19211 2149 19212
rect 2638 17781 2698 23971
rect 2822 19141 2882 26147
rect 3006 19277 3066 26691
rect 4208 26688 4528 27712
rect 5579 26892 5645 26893
rect 5579 26828 5580 26892
rect 5644 26828 5645 26892
rect 5579 26827 5645 26828
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4659 26348 4725 26349
rect 4659 26284 4660 26348
rect 4724 26284 4725 26348
rect 4659 26283 4725 26284
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 3923 24988 3989 24989
rect 3923 24924 3924 24988
rect 3988 24924 3989 24988
rect 3923 24923 3989 24924
rect 3555 24172 3621 24173
rect 3555 24108 3556 24172
rect 3620 24108 3621 24172
rect 3555 24107 3621 24108
rect 3187 23492 3253 23493
rect 3187 23428 3188 23492
rect 3252 23428 3253 23492
rect 3187 23427 3253 23428
rect 3003 19276 3069 19277
rect 3003 19212 3004 19276
rect 3068 19212 3069 19276
rect 3003 19211 3069 19212
rect 2819 19140 2885 19141
rect 2819 19076 2820 19140
rect 2884 19076 2885 19140
rect 2819 19075 2885 19076
rect 2635 17780 2701 17781
rect 2635 17716 2636 17780
rect 2700 17716 2701 17780
rect 2635 17715 2701 17716
rect 3190 12341 3250 23427
rect 3558 21045 3618 24107
rect 3739 23492 3805 23493
rect 3739 23428 3740 23492
rect 3804 23428 3805 23492
rect 3739 23427 3805 23428
rect 3742 21997 3802 23427
rect 3739 21996 3805 21997
rect 3739 21932 3740 21996
rect 3804 21932 3805 21996
rect 3739 21931 3805 21932
rect 3926 21453 3986 24923
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 3923 21452 3989 21453
rect 3923 21388 3924 21452
rect 3988 21388 3989 21452
rect 3923 21387 3989 21388
rect 3555 21044 3621 21045
rect 3555 20980 3556 21044
rect 3620 20980 3621 21044
rect 3555 20979 3621 20980
rect 3926 17645 3986 21387
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4662 20773 4722 26283
rect 4843 24988 4909 24989
rect 4843 24924 4844 24988
rect 4908 24924 4909 24988
rect 4843 24923 4909 24924
rect 4659 20772 4725 20773
rect 4659 20708 4660 20772
rect 4724 20708 4725 20772
rect 4659 20707 4725 20708
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4846 19413 4906 24923
rect 5027 21860 5093 21861
rect 5027 21796 5028 21860
rect 5092 21796 5093 21860
rect 5027 21795 5093 21796
rect 5030 19685 5090 21795
rect 5027 19684 5093 19685
rect 5027 19620 5028 19684
rect 5092 19620 5093 19684
rect 5027 19619 5093 19620
rect 4843 19412 4909 19413
rect 4843 19348 4844 19412
rect 4908 19348 4909 19412
rect 4843 19347 4909 19348
rect 4659 19276 4725 19277
rect 4659 19212 4660 19276
rect 4724 19212 4725 19276
rect 4659 19211 4725 19212
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4662 18325 4722 19211
rect 4659 18324 4725 18325
rect 4659 18260 4660 18324
rect 4724 18260 4725 18324
rect 4659 18259 4725 18260
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 3923 17644 3989 17645
rect 3923 17580 3924 17644
rect 3988 17580 3989 17644
rect 3923 17579 3989 17580
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4662 14245 4722 18259
rect 5582 15197 5642 26827
rect 5763 26484 5829 26485
rect 5763 26420 5764 26484
rect 5828 26420 5829 26484
rect 5763 26419 5829 26420
rect 5579 15196 5645 15197
rect 5579 15132 5580 15196
rect 5644 15132 5645 15196
rect 5579 15131 5645 15132
rect 4659 14244 4725 14245
rect 4659 14180 4660 14244
rect 4724 14180 4725 14244
rect 4659 14179 4725 14180
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 5766 12749 5826 26419
rect 10547 26348 10613 26349
rect 10547 26284 10548 26348
rect 10612 26284 10613 26348
rect 10547 26283 10613 26284
rect 9259 25260 9325 25261
rect 9259 25196 9260 25260
rect 9324 25196 9325 25260
rect 9259 25195 9325 25196
rect 7235 25124 7301 25125
rect 7235 25060 7236 25124
rect 7300 25060 7301 25124
rect 7235 25059 7301 25060
rect 7051 24988 7117 24989
rect 7051 24924 7052 24988
rect 7116 24924 7117 24988
rect 7051 24923 7117 24924
rect 5947 24852 6013 24853
rect 5947 24788 5948 24852
rect 6012 24788 6013 24852
rect 5947 24787 6013 24788
rect 5950 20365 6010 24787
rect 6499 22404 6565 22405
rect 6499 22340 6500 22404
rect 6564 22340 6565 22404
rect 6499 22339 6565 22340
rect 5947 20364 6013 20365
rect 5947 20300 5948 20364
rect 6012 20300 6013 20364
rect 5947 20299 6013 20300
rect 5763 12748 5829 12749
rect 5763 12684 5764 12748
rect 5828 12684 5829 12748
rect 5763 12683 5829 12684
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 3187 12340 3253 12341
rect 3187 12276 3188 12340
rect 3252 12276 3253 12340
rect 3187 12275 3253 12276
rect 4208 11456 4528 12480
rect 6502 11661 6562 22339
rect 6867 21996 6933 21997
rect 6867 21932 6868 21996
rect 6932 21932 6933 21996
rect 6867 21931 6933 21932
rect 6683 19412 6749 19413
rect 6683 19348 6684 19412
rect 6748 19348 6749 19412
rect 6683 19347 6749 19348
rect 6499 11660 6565 11661
rect 6499 11596 6500 11660
rect 6564 11596 6565 11660
rect 6499 11595 6565 11596
rect 6686 11525 6746 19347
rect 6870 14109 6930 21931
rect 7054 18189 7114 24923
rect 7051 18188 7117 18189
rect 7051 18124 7052 18188
rect 7116 18124 7117 18188
rect 7051 18123 7117 18124
rect 7051 17236 7117 17237
rect 7051 17172 7052 17236
rect 7116 17172 7117 17236
rect 7051 17171 7117 17172
rect 6867 14108 6933 14109
rect 6867 14044 6868 14108
rect 6932 14044 6933 14108
rect 6867 14043 6933 14044
rect 6683 11524 6749 11525
rect 6683 11460 6684 11524
rect 6748 11460 6749 11524
rect 6683 11459 6749 11460
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 1715 8668 1781 8669
rect 1715 8604 1716 8668
rect 1780 8604 1781 8668
rect 1715 8603 1781 8604
rect 4208 8192 4528 9216
rect 7054 8669 7114 17171
rect 7238 14517 7298 25059
rect 8891 24852 8957 24853
rect 8891 24788 8892 24852
rect 8956 24788 8957 24852
rect 8891 24787 8957 24788
rect 7603 23492 7669 23493
rect 7603 23428 7604 23492
rect 7668 23428 7669 23492
rect 7603 23427 7669 23428
rect 7606 17917 7666 23427
rect 7603 17916 7669 17917
rect 7603 17852 7604 17916
rect 7668 17852 7669 17916
rect 7603 17851 7669 17852
rect 7419 16148 7485 16149
rect 7419 16084 7420 16148
rect 7484 16084 7485 16148
rect 7419 16083 7485 16084
rect 7235 14516 7301 14517
rect 7235 14452 7236 14516
rect 7300 14452 7301 14516
rect 7235 14451 7301 14452
rect 7051 8668 7117 8669
rect 7051 8604 7052 8668
rect 7116 8604 7117 8668
rect 7051 8603 7117 8604
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 795 8124 861 8125
rect 795 8060 796 8124
rect 860 8060 861 8124
rect 795 8059 861 8060
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 7422 2685 7482 16083
rect 8894 15741 8954 24787
rect 9075 16420 9141 16421
rect 9075 16356 9076 16420
rect 9140 16356 9141 16420
rect 9075 16355 9141 16356
rect 8891 15740 8957 15741
rect 8891 15676 8892 15740
rect 8956 15676 8957 15740
rect 8891 15675 8957 15676
rect 9078 14517 9138 16355
rect 9262 15741 9322 25195
rect 9995 23492 10061 23493
rect 9995 23428 9996 23492
rect 10060 23428 10061 23492
rect 9995 23427 10061 23428
rect 10179 23492 10245 23493
rect 10179 23428 10180 23492
rect 10244 23428 10245 23492
rect 10179 23427 10245 23428
rect 9998 20501 10058 23427
rect 9995 20500 10061 20501
rect 9995 20436 9996 20500
rect 10060 20436 10061 20500
rect 9995 20435 10061 20436
rect 9443 16556 9509 16557
rect 9443 16492 9444 16556
rect 9508 16492 9509 16556
rect 9443 16491 9509 16492
rect 9259 15740 9325 15741
rect 9259 15676 9260 15740
rect 9324 15676 9325 15740
rect 9259 15675 9325 15676
rect 9075 14516 9141 14517
rect 9075 14452 9076 14516
rect 9140 14452 9141 14516
rect 9075 14451 9141 14452
rect 9446 10573 9506 16491
rect 10182 13293 10242 23427
rect 10550 14653 10610 26283
rect 10915 23628 10981 23629
rect 10915 23564 10916 23628
rect 10980 23564 10981 23628
rect 10915 23563 10981 23564
rect 11835 23628 11901 23629
rect 11835 23564 11836 23628
rect 11900 23564 11901 23628
rect 11835 23563 11901 23564
rect 10547 14652 10613 14653
rect 10547 14588 10548 14652
rect 10612 14588 10613 14652
rect 10547 14587 10613 14588
rect 10179 13292 10245 13293
rect 10179 13228 10180 13292
rect 10244 13228 10245 13292
rect 10179 13227 10245 13228
rect 9443 10572 9509 10573
rect 9443 10508 9444 10572
rect 9508 10508 9509 10572
rect 9443 10507 9509 10508
rect 10918 2685 10978 23563
rect 11099 22268 11165 22269
rect 11099 22204 11100 22268
rect 11164 22204 11165 22268
rect 11099 22203 11165 22204
rect 11102 21589 11162 22203
rect 11099 21588 11165 21589
rect 11099 21524 11100 21588
rect 11164 21524 11165 21588
rect 11099 21523 11165 21524
rect 11099 19548 11165 19549
rect 11099 19484 11100 19548
rect 11164 19484 11165 19548
rect 11099 19483 11165 19484
rect 11102 18325 11162 19483
rect 11099 18324 11165 18325
rect 11099 18260 11100 18324
rect 11164 18260 11165 18324
rect 11099 18259 11165 18260
rect 11838 15061 11898 23563
rect 12574 17237 12634 28051
rect 13123 27980 13189 27981
rect 13123 27916 13124 27980
rect 13188 27916 13189 27980
rect 13123 27915 13189 27916
rect 12571 17236 12637 17237
rect 12571 17172 12572 17236
rect 12636 17172 12637 17236
rect 12571 17171 12637 17172
rect 11835 15060 11901 15061
rect 11835 14996 11836 15060
rect 11900 14996 11901 15060
rect 11835 14995 11901 14996
rect 11838 13837 11898 14995
rect 11835 13836 11901 13837
rect 11835 13772 11836 13836
rect 11900 13772 11901 13836
rect 11835 13771 11901 13772
rect 13126 12885 13186 27915
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 16619 26212 16685 26213
rect 16619 26148 16620 26212
rect 16684 26148 16685 26212
rect 16619 26147 16685 26148
rect 15515 24988 15581 24989
rect 15515 24924 15516 24988
rect 15580 24924 15581 24988
rect 15515 24923 15581 24924
rect 14411 23084 14477 23085
rect 14411 23020 14412 23084
rect 14476 23020 14477 23084
rect 14411 23019 14477 23020
rect 13491 18052 13557 18053
rect 13491 17988 13492 18052
rect 13556 17988 13557 18052
rect 13491 17987 13557 17988
rect 13123 12884 13189 12885
rect 13123 12820 13124 12884
rect 13188 12820 13189 12884
rect 13123 12819 13189 12820
rect 13126 12477 13186 12819
rect 13123 12476 13189 12477
rect 13123 12412 13124 12476
rect 13188 12412 13189 12476
rect 13123 12411 13189 12412
rect 13494 2685 13554 17987
rect 14414 6629 14474 23019
rect 15518 11661 15578 24923
rect 16435 18732 16501 18733
rect 16435 18668 16436 18732
rect 16500 18668 16501 18732
rect 16435 18667 16501 18668
rect 16438 16013 16498 18667
rect 16435 16012 16501 16013
rect 16435 15948 16436 16012
rect 16500 15948 16501 16012
rect 16435 15947 16501 15948
rect 16622 15333 16682 26147
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 20115 22540 20181 22541
rect 20115 22476 20116 22540
rect 20180 22476 20181 22540
rect 20115 22475 20181 22476
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 17723 19276 17789 19277
rect 17723 19212 17724 19276
rect 17788 19212 17789 19276
rect 17723 19211 17789 19212
rect 16619 15332 16685 15333
rect 16619 15268 16620 15332
rect 16684 15268 16685 15332
rect 16619 15267 16685 15268
rect 16435 13428 16501 13429
rect 16435 13364 16436 13428
rect 16500 13364 16501 13428
rect 16435 13363 16501 13364
rect 15515 11660 15581 11661
rect 15515 11596 15516 11660
rect 15580 11596 15581 11660
rect 15515 11595 15581 11596
rect 16438 9621 16498 13363
rect 16435 9620 16501 9621
rect 16435 9556 16436 9620
rect 16500 9556 16501 9620
rect 16435 9555 16501 9556
rect 17726 6901 17786 19211
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 20118 12341 20178 22475
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 20115 12340 20181 12341
rect 20115 12276 20116 12340
rect 20180 12276 20181 12340
rect 20115 12275 20181 12276
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 17907 11660 17973 11661
rect 17907 11596 17908 11660
rect 17972 11596 17973 11660
rect 17907 11595 17973 11596
rect 17910 7309 17970 11595
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 17907 7308 17973 7309
rect 17907 7244 17908 7308
rect 17972 7244 17973 7308
rect 17907 7243 17973 7244
rect 17723 6900 17789 6901
rect 17723 6836 17724 6900
rect 17788 6836 17789 6900
rect 17723 6835 17789 6836
rect 14411 6628 14477 6629
rect 14411 6564 14412 6628
rect 14476 6564 14477 6628
rect 14411 6563 14477 6564
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19379 4316 19445 4317
rect 19379 4252 19380 4316
rect 19444 4252 19445 4316
rect 19379 4251 19445 4252
rect 19382 3501 19442 4251
rect 19379 3500 19445 3501
rect 19379 3436 19380 3500
rect 19444 3436 19445 3500
rect 19379 3435 19445 3436
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 7419 2684 7485 2685
rect 7419 2620 7420 2684
rect 7484 2620 7485 2684
rect 7419 2619 7485 2620
rect 10915 2684 10981 2685
rect 10915 2620 10916 2684
rect 10980 2620 10981 2684
rect 10915 2619 10981 2620
rect 13491 2684 13557 2685
rect 13491 2620 13492 2684
rect 13556 2620 13557 2684
rect 13491 2619 13557 2620
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11592 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform 1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1667941163
transform 1 0 35788 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1667941163
transform 1 0 2116 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1667941163
transform 1 0 35420 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17
timestamp 1667941163
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34
timestamp 1667941163
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41
timestamp 1667941163
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68
timestamp 1667941163
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1667941163
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91
timestamp 1667941163
transform 1 0 9476 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95
timestamp 1667941163
transform 1 0 9844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102
timestamp 1667941163
transform 1 0 10488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1667941163
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119
timestamp 1667941163
transform 1 0 12052 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_130
timestamp 1667941163
transform 1 0 13064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1667941163
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1667941163
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_174
timestamp 1667941163
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1667941163
transform 1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_190
timestamp 1667941163
transform 1 0 18584 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1667941163
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_214
timestamp 1667941163
transform 1 0 20792 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1667941163
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1667941163
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_238
timestamp 1667941163
transform 1 0 23000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245
timestamp 1667941163
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1667941163
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_258
timestamp 1667941163
transform 1 0 24840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_266
timestamp 1667941163
transform 1 0 25576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_274
timestamp 1667941163
transform 1 0 26312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1667941163
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_293
timestamp 1667941163
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1667941163
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1667941163
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_315
timestamp 1667941163
transform 1 0 30084 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_322 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 30728 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1667941163
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1667941163
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_357
timestamp 1667941163
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1667941163
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_371
timestamp 1667941163
transform 1 0 35236 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_379
timestamp 1667941163
transform 1 0 35972 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1667941163
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1667941163
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_20
timestamp 1667941163
transform 1 0 2944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1667941163
transform 1 0 3588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_34
timestamp 1667941163
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_41
timestamp 1667941163
transform 1 0 4876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49
timestamp 1667941163
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1667941163
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_63
timestamp 1667941163
transform 1 0 6900 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_67
timestamp 1667941163
transform 1 0 7268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_74
timestamp 1667941163
transform 1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_81
timestamp 1667941163
transform 1 0 8556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1667941163
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1667941163
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_119
timestamp 1667941163
transform 1 0 12052 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_123
timestamp 1667941163
transform 1 0 12420 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_152
timestamp 1667941163
transform 1 0 15088 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_156
timestamp 1667941163
transform 1 0 15456 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1667941163
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_180
timestamp 1667941163
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1667941163
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_204
timestamp 1667941163
transform 1 0 19872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1667941163
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1667941163
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_230
timestamp 1667941163
transform 1 0 22264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_244
timestamp 1667941163
transform 1 0 23552 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_251
timestamp 1667941163
transform 1 0 24196 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_258
timestamp 1667941163
transform 1 0 24840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_265
timestamp 1667941163
transform 1 0 25484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_272
timestamp 1667941163
transform 1 0 26128 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_286
timestamp 1667941163
transform 1 0 27416 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_298
timestamp 1667941163
transform 1 0 28520 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_310
timestamp 1667941163
transform 1 0 29624 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_322
timestamp 1667941163
transform 1 0 30728 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1667941163
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_357
timestamp 1667941163
transform 1 0 33948 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_369
timestamp 1667941163
transform 1 0 35052 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_381
timestamp 1667941163
transform 1 0 36156 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1667941163
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_398
timestamp 1667941163
transform 1 0 37720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_12
timestamp 1667941163
transform 1 0 2208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_19
timestamp 1667941163
transform 1 0 2852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1667941163
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_33
timestamp 1667941163
transform 1 0 4140 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_37
timestamp 1667941163
transform 1 0 4508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_44
timestamp 1667941163
transform 1 0 5152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_51
timestamp 1667941163
transform 1 0 5796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_58
timestamp 1667941163
transform 1 0 6440 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1667941163
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_92
timestamp 1667941163
transform 1 0 9568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_99
timestamp 1667941163
transform 1 0 10212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_106
timestamp 1667941163
transform 1 0 10856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1667941163
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1667941163
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_163
timestamp 1667941163
transform 1 0 16100 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1667941163
transform 1 0 17664 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_187
timestamp 1667941163
transform 1 0 18308 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1667941163
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_203
timestamp 1667941163
transform 1 0 19780 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_210
timestamp 1667941163
transform 1 0 20424 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_217
timestamp 1667941163
transform 1 0 21068 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_224
timestamp 1667941163
transform 1 0 21712 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_231
timestamp 1667941163
transform 1 0 22356 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_238
timestamp 1667941163
transform 1 0 23000 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1667941163
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1667941163
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_258
timestamp 1667941163
transform 1 0 24840 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_272
timestamp 1667941163
transform 1 0 26128 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_279
timestamp 1667941163
transform 1 0 26772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_291
timestamp 1667941163
transform 1 0 27876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_303
timestamp 1667941163
transform 1 0 28980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_389
timestamp 1667941163
transform 1 0 36892 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_398
timestamp 1667941163
transform 1 0 37720 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_9
timestamp 1667941163
transform 1 0 1932 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_20
timestamp 1667941163
transform 1 0 2944 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_45
timestamp 1667941163
transform 1 0 5244 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1667941163
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1667941163
transform 1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_86
timestamp 1667941163
transform 1 0 9016 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1667941163
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_117
timestamp 1667941163
transform 1 0 11868 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_121
timestamp 1667941163
transform 1 0 12236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_128
timestamp 1667941163
transform 1 0 12880 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_155
timestamp 1667941163
transform 1 0 15364 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1667941163
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_191
timestamp 1667941163
transform 1 0 18676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_200
timestamp 1667941163
transform 1 0 19504 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_207
timestamp 1667941163
transform 1 0 20148 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_214
timestamp 1667941163
transform 1 0 20792 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_221
timestamp 1667941163
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_230
timestamp 1667941163
transform 1 0 22264 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_244
timestamp 1667941163
transform 1 0 23552 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_251
timestamp 1667941163
transform 1 0 24196 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_258
timestamp 1667941163
transform 1 0 24840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_265
timestamp 1667941163
transform 1 0 25484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_272
timestamp 1667941163
transform 1 0 26128 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_401
timestamp 1667941163
transform 1 0 37996 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1667941163
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_34
timestamp 1667941163
transform 1 0 4232 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_43
timestamp 1667941163
transform 1 0 5060 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_50
timestamp 1667941163
transform 1 0 5704 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_113
timestamp 1667941163
transform 1 0 11500 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_117
timestamp 1667941163
transform 1 0 11868 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1667941163
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_163
timestamp 1667941163
transform 1 0 16100 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_176
timestamp 1667941163
transform 1 0 17296 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_184
timestamp 1667941163
transform 1 0 18032 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1667941163
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_207
timestamp 1667941163
transform 1 0 20148 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_214
timestamp 1667941163
transform 1 0 20792 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_228
timestamp 1667941163
transform 1 0 22080 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_235
timestamp 1667941163
transform 1 0 22724 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_242
timestamp 1667941163
transform 1 0 23368 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1667941163
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_258
timestamp 1667941163
transform 1 0 24840 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1667941163
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_397
timestamp 1667941163
transform 1 0 37628 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_402
timestamp 1667941163
transform 1 0 38088 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_406
timestamp 1667941163
transform 1 0 38456 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_15
timestamp 1667941163
transform 1 0 2484 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_23
timestamp 1667941163
transform 1 0 3220 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1667941163
transform 1 0 3588 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1667941163
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1667941163
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_74
timestamp 1667941163
transform 1 0 7912 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_98
timestamp 1667941163
transform 1 0 10120 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_106
timestamp 1667941163
transform 1 0 10856 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1667941163
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_130
timestamp 1667941163
transform 1 0 13064 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_154
timestamp 1667941163
transform 1 0 15272 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1667941163
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_184
timestamp 1667941163
transform 1 0 18032 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_197
timestamp 1667941163
transform 1 0 19228 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_203
timestamp 1667941163
transform 1 0 19780 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_213
timestamp 1667941163
transform 1 0 20700 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1667941163
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_236
timestamp 1667941163
transform 1 0 22816 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_243
timestamp 1667941163
transform 1 0 23460 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_250
timestamp 1667941163
transform 1 0 24104 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_262
timestamp 1667941163
transform 1 0 25208 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_270
timestamp 1667941163
transform 1 0 25944 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1667941163
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_312
timestamp 1667941163
transform 1 0 29808 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_319
timestamp 1667941163
transform 1 0 30452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_331
timestamp 1667941163
transform 1 0 31556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp 1667941163
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_34
timestamp 1667941163
transform 1 0 4232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_68
timestamp 1667941163
transform 1 0 7360 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_75
timestamp 1667941163
transform 1 0 8004 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1667941163
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_163
timestamp 1667941163
transform 1 0 16100 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_180
timestamp 1667941163
transform 1 0 17664 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 1667941163
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_205
timestamp 1667941163
transform 1 0 19964 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_212
timestamp 1667941163
transform 1 0 20608 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_219
timestamp 1667941163
transform 1 0 21252 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_226
timestamp 1667941163
transform 1 0 21896 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_240
timestamp 1667941163
transform 1 0 23184 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_247
timestamp 1667941163
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_270
timestamp 1667941163
transform 1 0 25944 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_282
timestamp 1667941163
transform 1 0 27048 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_294
timestamp 1667941163
transform 1 0 28152 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1667941163
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1667941163
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_401
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1667941163
transform 1 0 1748 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_11
timestamp 1667941163
transform 1 0 2116 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_18
timestamp 1667941163
transform 1 0 2760 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_27
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_35
timestamp 1667941163
transform 1 0 4324 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_39
timestamp 1667941163
transform 1 0 4692 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1667941163
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_79
timestamp 1667941163
transform 1 0 8372 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_83
timestamp 1667941163
transform 1 0 8740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_106
timestamp 1667941163
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_126
timestamp 1667941163
transform 1 0 12696 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_154
timestamp 1667941163
transform 1 0 15272 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1667941163
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_174
timestamp 1667941163
transform 1 0 17112 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_178
timestamp 1667941163
transform 1 0 17480 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_192
timestamp 1667941163
transform 1 0 18768 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_204
timestamp 1667941163
transform 1 0 19872 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_211
timestamp 1667941163
transform 1 0 20516 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_218
timestamp 1667941163
transform 1 0 21160 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_231
timestamp 1667941163
transform 1 0 22356 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_241
timestamp 1667941163
transform 1 0 23276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_253
timestamp 1667941163
transform 1 0 24380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_265
timestamp 1667941163
transform 1 0 25484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_277
timestamp 1667941163
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_323
timestamp 1667941163
transform 1 0 30820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_401
timestamp 1667941163
transform 1 0 37996 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_9
timestamp 1667941163
transform 1 0 1932 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_16
timestamp 1667941163
transform 1 0 2576 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1667941163
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_34
timestamp 1667941163
transform 1 0 4232 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_42
timestamp 1667941163
transform 1 0 4968 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_74
timestamp 1667941163
transform 1 0 7912 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1667941163
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_91
timestamp 1667941163
transform 1 0 9476 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_98
timestamp 1667941163
transform 1 0 10120 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_105
timestamp 1667941163
transform 1 0 10764 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_129
timestamp 1667941163
transform 1 0 12972 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1667941163
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_163
timestamp 1667941163
transform 1 0 16100 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_176
timestamp 1667941163
transform 1 0 17296 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_208
timestamp 1667941163
transform 1 0 20240 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1667941163
transform 1 0 20884 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_222
timestamp 1667941163
transform 1 0 21528 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_229
timestamp 1667941163
transform 1 0 22172 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_236
timestamp 1667941163
transform 1 0 22816 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_243
timestamp 1667941163
transform 1 0 23460 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1667941163
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1667941163
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1667941163
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1667941163
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_9
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_17
timestamp 1667941163
transform 1 0 2668 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_38
timestamp 1667941163
transform 1 0 4600 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_50
timestamp 1667941163
transform 1 0 5704 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1667941163
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_80
timestamp 1667941163
transform 1 0 8464 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_104
timestamp 1667941163
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_136
timestamp 1667941163
transform 1 0 13616 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_160
timestamp 1667941163
transform 1 0 15824 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_188
timestamp 1667941163
transform 1 0 18400 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_205
timestamp 1667941163
transform 1 0 19964 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_213
timestamp 1667941163
transform 1 0 20700 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1667941163
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_235
timestamp 1667941163
transform 1 0 22724 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_242
timestamp 1667941163
transform 1 0 23368 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_261
timestamp 1667941163
transform 1 0 25116 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_267
timestamp 1667941163
transform 1 0 25668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1667941163
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_286
timestamp 1667941163
transform 1 0 27416 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_298
timestamp 1667941163
transform 1 0 28520 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_310
timestamp 1667941163
transform 1 0 29624 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_322
timestamp 1667941163
transform 1 0 30728 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp 1667941163
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1667941163
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_35
timestamp 1667941163
transform 1 0 4324 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_47
timestamp 1667941163
transform 1 0 5428 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_51
timestamp 1667941163
transform 1 0 5796 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_55
timestamp 1667941163
transform 1 0 6164 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_64
timestamp 1667941163
transform 1 0 6992 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_76
timestamp 1667941163
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1667941163
transform 1 0 9476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_112
timestamp 1667941163
transform 1 0 11408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_116
timestamp 1667941163
transform 1 0 11776 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1667941163
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_163
timestamp 1667941163
transform 1 0 16100 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_180
timestamp 1667941163
transform 1 0 17664 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_184
timestamp 1667941163
transform 1 0 18032 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1667941163
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_202
timestamp 1667941163
transform 1 0 19688 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_219
timestamp 1667941163
transform 1 0 21252 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_236
timestamp 1667941163
transform 1 0 22816 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_243
timestamp 1667941163
transform 1 0 23460 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1667941163
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_258
timestamp 1667941163
transform 1 0 24840 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_270
timestamp 1667941163
transform 1 0 25944 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_282
timestamp 1667941163
transform 1 0 27048 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_294
timestamp 1667941163
transform 1 0 28152 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1667941163
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_314
timestamp 1667941163
transform 1 0 29992 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_326
timestamp 1667941163
transform 1 0 31096 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_338
timestamp 1667941163
transform 1 0 32200 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_350
timestamp 1667941163
transform 1 0 33304 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp 1667941163
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1667941163
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_8
timestamp 1667941163
transform 1 0 1840 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_32
timestamp 1667941163
transform 1 0 4048 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_39
timestamp 1667941163
transform 1 0 4692 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_46
timestamp 1667941163
transform 1 0 5336 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1667941163
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_62
timestamp 1667941163
transform 1 0 6808 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_86
timestamp 1667941163
transform 1 0 9016 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1667941163
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_135
timestamp 1667941163
transform 1 0 13524 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_159
timestamp 1667941163
transform 1 0 15732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1667941163
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_180
timestamp 1667941163
transform 1 0 17664 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_190
timestamp 1667941163
transform 1 0 18584 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_196
timestamp 1667941163
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_210
timestamp 1667941163
transform 1 0 20424 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_219
timestamp 1667941163
transform 1 0 21252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1667941163
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_230
timestamp 1667941163
transform 1 0 22264 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1667941163
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_251
timestamp 1667941163
transform 1 0 24196 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_258
timestamp 1667941163
transform 1 0 24840 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_265
timestamp 1667941163
transform 1 0 25484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp 1667941163
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_12
timestamp 1667941163
transform 1 0 2208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_19
timestamp 1667941163
transform 1 0 2852 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1667941163
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_42
timestamp 1667941163
transform 1 0 4968 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_49
timestamp 1667941163
transform 1 0 5612 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_57
timestamp 1667941163
transform 1 0 6348 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_62
timestamp 1667941163
transform 1 0 6808 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_70
timestamp 1667941163
transform 1 0 7544 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1667941163
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_92
timestamp 1667941163
transform 1 0 9568 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_117
timestamp 1667941163
transform 1 0 11868 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_123
timestamp 1667941163
transform 1 0 12420 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_127
timestamp 1667941163
transform 1 0 12788 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 1667941163
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_163
timestamp 1667941163
transform 1 0 16100 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_180
timestamp 1667941163
transform 1 0 17664 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_193
timestamp 1667941163
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_201
timestamp 1667941163
transform 1 0 19596 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_205
timestamp 1667941163
transform 1 0 19964 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_213
timestamp 1667941163
transform 1 0 20700 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_224
timestamp 1667941163
transform 1 0 21712 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_231
timestamp 1667941163
transform 1 0 22356 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_238
timestamp 1667941163
transform 1 0 23000 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_258
timestamp 1667941163
transform 1 0 24840 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_270
timestamp 1667941163
transform 1 0 25944 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_282
timestamp 1667941163
transform 1 0 27048 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_294
timestamp 1667941163
transform 1 0 28152 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1667941163
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_401
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_26
timestamp 1667941163
transform 1 0 3496 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1667941163
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_74
timestamp 1667941163
transform 1 0 7912 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_78
timestamp 1667941163
transform 1 0 8280 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_82
timestamp 1667941163
transform 1 0 8648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1667941163
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_126
timestamp 1667941163
transform 1 0 12696 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_130
timestamp 1667941163
transform 1 0 13064 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_134
timestamp 1667941163
transform 1 0 13432 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_159
timestamp 1667941163
transform 1 0 15732 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1667941163
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_175
timestamp 1667941163
transform 1 0 17204 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_179
timestamp 1667941163
transform 1 0 17572 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_188
timestamp 1667941163
transform 1 0 18400 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_199
timestamp 1667941163
transform 1 0 19412 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_206
timestamp 1667941163
transform 1 0 20056 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_212
timestamp 1667941163
transform 1 0 20608 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1667941163
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_230
timestamp 1667941163
transform 1 0 22264 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_241
timestamp 1667941163
transform 1 0 23276 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_245
timestamp 1667941163
transform 1 0 23644 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_252
timestamp 1667941163
transform 1 0 24288 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_271
timestamp 1667941163
transform 1 0 26036 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_316
timestamp 1667941163
transform 1 0 30176 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_328
timestamp 1667941163
transform 1 0 31280 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_12
timestamp 1667941163
transform 1 0 2208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_19
timestamp 1667941163
transform 1 0 2852 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1667941163
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_51
timestamp 1667941163
transform 1 0 5796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_57
timestamp 1667941163
transform 1 0 6348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_78
timestamp 1667941163
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1667941163
transform 1 0 9476 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_95
timestamp 1667941163
transform 1 0 9844 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_102
timestamp 1667941163
transform 1 0 10488 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_129
timestamp 1667941163
transform 1 0 12972 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1667941163
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_164
timestamp 1667941163
transform 1 0 16192 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_179
timestamp 1667941163
transform 1 0 17572 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1667941163
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1667941163
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_212
timestamp 1667941163
transform 1 0 20608 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_225
timestamp 1667941163
transform 1 0 21804 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_229
timestamp 1667941163
transform 1 0 22172 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_238
timestamp 1667941163
transform 1 0 23000 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1667941163
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1667941163
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_259
timestamp 1667941163
transform 1 0 24932 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_263
timestamp 1667941163
transform 1 0 25300 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_275
timestamp 1667941163
transform 1 0 26404 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_287
timestamp 1667941163
transform 1 0 27508 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_299
timestamp 1667941163
transform 1 0 28612 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_314
timestamp 1667941163
transform 1 0 29992 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_326
timestamp 1667941163
transform 1 0 31096 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_338
timestamp 1667941163
transform 1 0 32200 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_350
timestamp 1667941163
transform 1 0 33304 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_362
timestamp 1667941163
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_405
timestamp 1667941163
transform 1 0 38364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1667941163
transform 1 0 1748 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_11
timestamp 1667941163
transform 1 0 2116 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_18
timestamp 1667941163
transform 1 0 2760 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_25
timestamp 1667941163
transform 1 0 3404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_49
timestamp 1667941163
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1667941163
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1667941163
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_125
timestamp 1667941163
transform 1 0 12604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_152
timestamp 1667941163
transform 1 0 15088 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_156
timestamp 1667941163
transform 1 0 15456 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1667941163
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_179
timestamp 1667941163
transform 1 0 17572 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1667941163
transform 1 0 19136 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1667941163
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1667941163
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_230
timestamp 1667941163
transform 1 0 22264 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_237
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_246
timestamp 1667941163
transform 1 0 23736 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_257
timestamp 1667941163
transform 1 0 24748 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_269
timestamp 1667941163
transform 1 0 25852 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_277
timestamp 1667941163
transform 1 0 26588 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1667941163
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1667941163
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1667941163
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1667941163
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_25
timestamp 1667941163
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_55
timestamp 1667941163
transform 1 0 6164 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1667941163
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_90
timestamp 1667941163
transform 1 0 9384 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_114
timestamp 1667941163
transform 1 0 11592 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1667941163
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_164
timestamp 1667941163
transform 1 0 16192 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_181
timestamp 1667941163
transform 1 0 17756 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_191
timestamp 1667941163
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_208
timestamp 1667941163
transform 1 0 20240 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1667941163
transform 1 0 20884 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_222
timestamp 1667941163
transform 1 0 21528 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_229
timestamp 1667941163
transform 1 0 22172 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_236
timestamp 1667941163
transform 1 0 22816 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_243
timestamp 1667941163
transform 1 0 23460 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_274
timestamp 1667941163
transform 1 0 26312 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_286
timestamp 1667941163
transform 1 0 27416 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_298
timestamp 1667941163
transform 1 0 28520 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1667941163
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_405
timestamp 1667941163
transform 1 0 38364 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1667941163
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_30
timestamp 1667941163
transform 1 0 3864 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1667941163
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_62
timestamp 1667941163
transform 1 0 6808 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_86
timestamp 1667941163
transform 1 0 9016 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1667941163
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1667941163
transform 1 0 11960 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_125
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_152
timestamp 1667941163
transform 1 0 15088 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_156
timestamp 1667941163
transform 1 0 15456 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1667941163
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_180
timestamp 1667941163
transform 1 0 17664 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_190
timestamp 1667941163
transform 1 0 18584 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_200
timestamp 1667941163
transform 1 0 19504 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_208
timestamp 1667941163
transform 1 0 20240 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_213
timestamp 1667941163
transform 1 0 20700 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1667941163
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_240
timestamp 1667941163
transform 1 0 23184 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_247
timestamp 1667941163
transform 1 0 23828 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_259
timestamp 1667941163
transform 1 0 24932 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_271
timestamp 1667941163
transform 1 0 26036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1667941163
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1667941163
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1667941163
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1667941163
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1667941163
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_42
timestamp 1667941163
transform 1 0 4968 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_69
timestamp 1667941163
transform 1 0 7452 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_76
timestamp 1667941163
transform 1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_90
timestamp 1667941163
transform 1 0 9384 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_114
timestamp 1667941163
transform 1 0 11592 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1667941163
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_163
timestamp 1667941163
transform 1 0 16100 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_176
timestamp 1667941163
transform 1 0 17296 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1667941163
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1667941163
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_202
timestamp 1667941163
transform 1 0 19688 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_210
timestamp 1667941163
transform 1 0 20424 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_224
timestamp 1667941163
transform 1 0 21712 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_231
timestamp 1667941163
transform 1 0 22356 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_243
timestamp 1667941163
transform 1 0 23460 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1667941163
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_257
timestamp 1667941163
transform 1 0 24748 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_266
timestamp 1667941163
transform 1 0 25576 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_278
timestamp 1667941163
transform 1 0 26680 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_283
timestamp 1667941163
transform 1 0 27140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_295
timestamp 1667941163
transform 1 0 28244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1667941163
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1667941163
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1667941163
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1667941163
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_26
timestamp 1667941163
transform 1 0 3496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 1667941163
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_63
timestamp 1667941163
transform 1 0 6900 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_90
timestamp 1667941163
transform 1 0 9384 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_94
timestamp 1667941163
transform 1 0 9752 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_106
timestamp 1667941163
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_118
timestamp 1667941163
transform 1 0 11960 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_124
timestamp 1667941163
transform 1 0 12512 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_128
timestamp 1667941163
transform 1 0 12880 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp 1667941163
transform 1 0 15180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1667941163
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_180
timestamp 1667941163
transform 1 0 17664 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_197
timestamp 1667941163
transform 1 0 19228 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_210
timestamp 1667941163
transform 1 0 20424 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1667941163
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1667941163
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_232
timestamp 1667941163
transform 1 0 22448 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_244
timestamp 1667941163
transform 1 0 23552 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_256
timestamp 1667941163
transform 1 0 24656 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_268
timestamp 1667941163
transform 1 0 25760 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_290
timestamp 1667941163
transform 1 0 27784 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_297
timestamp 1667941163
transform 1 0 28428 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_309
timestamp 1667941163
transform 1 0 29532 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_321
timestamp 1667941163
transform 1 0 30636 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_333
timestamp 1667941163
transform 1 0 31740 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1667941163
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_78
timestamp 1667941163
transform 1 0 8280 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_111
timestamp 1667941163
transform 1 0 11316 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1667941163
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_156
timestamp 1667941163
transform 1 0 15456 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_171
timestamp 1667941163
transform 1 0 16836 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_186
timestamp 1667941163
transform 1 0 18216 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1667941163
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_208
timestamp 1667941163
transform 1 0 20240 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_215
timestamp 1667941163
transform 1 0 20884 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_227
timestamp 1667941163
transform 1 0 21988 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_231
timestamp 1667941163
transform 1 0 22356 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_243
timestamp 1667941163
transform 1 0 23460 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1667941163
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_265
timestamp 1667941163
transform 1 0 25484 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_279
timestamp 1667941163
transform 1 0 26772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_291
timestamp 1667941163
transform 1 0 27876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1667941163
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_357
timestamp 1667941163
transform 1 0 33948 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1667941163
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_405
timestamp 1667941163
transform 1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_9
timestamp 1667941163
transform 1 0 1932 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_13
timestamp 1667941163
transform 1 0 2300 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_39
timestamp 1667941163
transform 1 0 4692 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_46
timestamp 1667941163
transform 1 0 5336 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1667941163
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_63
timestamp 1667941163
transform 1 0 6900 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_70
timestamp 1667941163
transform 1 0 7544 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_77
timestamp 1667941163
transform 1 0 8188 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_102
timestamp 1667941163
transform 1 0 10488 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_109
timestamp 1667941163
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_117
timestamp 1667941163
transform 1 0 11868 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_139
timestamp 1667941163
transform 1 0 13892 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_145
timestamp 1667941163
transform 1 0 14444 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_159
timestamp 1667941163
transform 1 0 15732 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1667941163
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_175
timestamp 1667941163
transform 1 0 17204 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_188
timestamp 1667941163
transform 1 0 18400 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_198
timestamp 1667941163
transform 1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_205
timestamp 1667941163
transform 1 0 19964 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1667941163
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_230
timestamp 1667941163
transform 1 0 22264 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_242
timestamp 1667941163
transform 1 0 23368 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_254
timestamp 1667941163
transform 1 0 24472 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_266
timestamp 1667941163
transform 1 0 25576 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1667941163
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1667941163
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1667941163
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1667941163
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_25
timestamp 1667941163
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_42
timestamp 1667941163
transform 1 0 4968 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_50
timestamp 1667941163
transform 1 0 5704 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_57
timestamp 1667941163
transform 1 0 6348 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1667941163
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_107
timestamp 1667941163
transform 1 0 10948 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_114
timestamp 1667941163
transform 1 0 11592 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_133
timestamp 1667941163
transform 1 0 13340 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1667941163
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1667941163
transform 1 0 16100 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_167
timestamp 1667941163
transform 1 0 16468 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_176
timestamp 1667941163
transform 1 0 17296 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1667941163
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1667941163
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_202
timestamp 1667941163
transform 1 0 19688 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_210
timestamp 1667941163
transform 1 0 20424 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1667941163
transform 1 0 20884 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_222
timestamp 1667941163
transform 1 0 21528 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_229
timestamp 1667941163
transform 1 0 22172 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_241
timestamp 1667941163
transform 1 0 23276 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_249
timestamp 1667941163
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_257
timestamp 1667941163
transform 1 0 24748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_266
timestamp 1667941163
transform 1 0 25576 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_278
timestamp 1667941163
transform 1 0 26680 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_285
timestamp 1667941163
transform 1 0 27324 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_297
timestamp 1667941163
transform 1 0 28428 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_305
timestamp 1667941163
transform 1 0 29164 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1667941163
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1667941163
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1667941163
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_405
timestamp 1667941163
transform 1 0 38364 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_25
timestamp 1667941163
transform 1 0 3404 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_49
timestamp 1667941163
transform 1 0 5612 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_61
timestamp 1667941163
transform 1 0 6716 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_82
timestamp 1667941163
transform 1 0 8648 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_107
timestamp 1667941163
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_119
timestamp 1667941163
transform 1 0 12052 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_140
timestamp 1667941163
transform 1 0 13984 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_148
timestamp 1667941163
transform 1 0 14720 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_152
timestamp 1667941163
transform 1 0 15088 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_159
timestamp 1667941163
transform 1 0 15732 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1667941163
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_184
timestamp 1667941163
transform 1 0 18032 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_194
timestamp 1667941163
transform 1 0 18952 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_201
timestamp 1667941163
transform 1 0 19596 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_208
timestamp 1667941163
transform 1 0 20240 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_215
timestamp 1667941163
transform 1 0 20884 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1667941163
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_230
timestamp 1667941163
transform 1 0 22264 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_242
timestamp 1667941163
transform 1 0 23368 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_254
timestamp 1667941163
transform 1 0 24472 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_266
timestamp 1667941163
transform 1 0 25576 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_270
timestamp 1667941163
transform 1 0 25944 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1667941163
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_289
timestamp 1667941163
transform 1 0 27692 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1667941163
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1667941163
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1667941163
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1667941163
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_25
timestamp 1667941163
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1667941163
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_90
timestamp 1667941163
transform 1 0 9384 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_124
timestamp 1667941163
transform 1 0 12512 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_131
timestamp 1667941163
transform 1 0 13156 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1667941163
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_148
timestamp 1667941163
transform 1 0 14720 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_165
timestamp 1667941163
transform 1 0 16284 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_169
timestamp 1667941163
transform 1 0 16652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_176
timestamp 1667941163
transform 1 0 17296 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_184
timestamp 1667941163
transform 1 0 18032 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1667941163
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_202
timestamp 1667941163
transform 1 0 19688 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_209
timestamp 1667941163
transform 1 0 20332 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_215
timestamp 1667941163
transform 1 0 20884 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1667941163
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_236
timestamp 1667941163
transform 1 0 22816 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1667941163
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1667941163
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_277
timestamp 1667941163
transform 1 0 26588 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_285
timestamp 1667941163
transform 1 0 27324 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_291
timestamp 1667941163
transform 1 0 27876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_303
timestamp 1667941163
transform 1 0 28980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1667941163
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_314
timestamp 1667941163
transform 1 0 29992 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_326
timestamp 1667941163
transform 1 0 31096 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_338
timestamp 1667941163
transform 1 0 32200 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_350
timestamp 1667941163
transform 1 0 33304 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1667941163
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_30
timestamp 1667941163
transform 1 0 3864 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1667941163
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_62
timestamp 1667941163
transform 1 0 6808 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_89
timestamp 1667941163
transform 1 0 9292 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_96
timestamp 1667941163
transform 1 0 9936 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_103
timestamp 1667941163
transform 1 0 10580 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1667941163
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1667941163
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_131
timestamp 1667941163
transform 1 0 13156 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_156
timestamp 1667941163
transform 1 0 15456 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_162
timestamp 1667941163
transform 1 0 16008 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1667941163
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_177
timestamp 1667941163
transform 1 0 17388 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_194
timestamp 1667941163
transform 1 0 18952 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_201
timestamp 1667941163
transform 1 0 19596 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_208
timestamp 1667941163
transform 1 0 20240 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_212
timestamp 1667941163
transform 1 0 20608 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_216
timestamp 1667941163
transform 1 0 20976 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_240
timestamp 1667941163
transform 1 0 23184 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_252
timestamp 1667941163
transform 1 0 24288 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_264
timestamp 1667941163
transform 1 0 25392 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1667941163
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_286
timestamp 1667941163
transform 1 0 27416 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_290
timestamp 1667941163
transform 1 0 27784 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_294
timestamp 1667941163
transform 1 0 28152 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_301
timestamp 1667941163
transform 1 0 28796 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_313
timestamp 1667941163
transform 1 0 29900 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_325
timestamp 1667941163
transform 1 0 31004 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_333
timestamp 1667941163
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1667941163
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_401
timestamp 1667941163
transform 1 0 37996 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1667941163
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_34
timestamp 1667941163
transform 1 0 4232 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_58
timestamp 1667941163
transform 1 0 6440 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1667941163
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_98
timestamp 1667941163
transform 1 0 10120 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_125
timestamp 1667941163
transform 1 0 12604 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_133
timestamp 1667941163
transform 1 0 13340 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1667941163
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_163
timestamp 1667941163
transform 1 0 16100 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_174
timestamp 1667941163
transform 1 0 17112 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_181
timestamp 1667941163
transform 1 0 17756 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_189
timestamp 1667941163
transform 1 0 18492 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1667941163
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_212
timestamp 1667941163
transform 1 0 20608 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_224
timestamp 1667941163
transform 1 0 21712 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_235
timestamp 1667941163
transform 1 0 22724 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_247
timestamp 1667941163
transform 1 0 23828 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1667941163
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_263
timestamp 1667941163
transform 1 0 25300 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_275
timestamp 1667941163
transform 1 0 26404 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_287
timestamp 1667941163
transform 1 0 27508 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_299
timestamp 1667941163
transform 1 0 28612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1667941163
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_405
timestamp 1667941163
transform 1 0 38364 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_29
timestamp 1667941163
transform 1 0 3772 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_33
timestamp 1667941163
transform 1 0 4140 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1667941163
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_80
timestamp 1667941163
transform 1 0 8464 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp 1667941163
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_117
timestamp 1667941163
transform 1 0 11868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_139
timestamp 1667941163
transform 1 0 13892 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_163
timestamp 1667941163
transform 1 0 16100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1667941163
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_176
timestamp 1667941163
transform 1 0 17296 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_183
timestamp 1667941163
transform 1 0 17940 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_190
timestamp 1667941163
transform 1 0 18584 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_203
timestamp 1667941163
transform 1 0 19780 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_210
timestamp 1667941163
transform 1 0 20424 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1667941163
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_240
timestamp 1667941163
transform 1 0 23184 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_252
timestamp 1667941163
transform 1 0 24288 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_258
timestamp 1667941163
transform 1 0 24840 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_262
timestamp 1667941163
transform 1 0 25208 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_274
timestamp 1667941163
transform 1 0 26312 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_291
timestamp 1667941163
transform 1 0 27876 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_298
timestamp 1667941163
transform 1 0 28520 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_310
timestamp 1667941163
transform 1 0 29624 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_322
timestamp 1667941163
transform 1 0 30728 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1667941163
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_25
timestamp 1667941163
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_51
timestamp 1667941163
transform 1 0 5796 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_58
timestamp 1667941163
transform 1 0 6440 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1667941163
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_112
timestamp 1667941163
transform 1 0 11408 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1667941163
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_146
timestamp 1667941163
transform 1 0 14536 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_159
timestamp 1667941163
transform 1 0 15732 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_172
timestamp 1667941163
transform 1 0 16928 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_179
timestamp 1667941163
transform 1 0 17572 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_186
timestamp 1667941163
transform 1 0 18216 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1667941163
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_212
timestamp 1667941163
transform 1 0 20608 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_224
timestamp 1667941163
transform 1 0 21712 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_230
timestamp 1667941163
transform 1 0 22264 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_240
timestamp 1667941163
transform 1 0 23184 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1667941163
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_289
timestamp 1667941163
transform 1 0 27692 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_294
timestamp 1667941163
transform 1 0 28152 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 1667941163
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_317
timestamp 1667941163
transform 1 0 30268 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_323
timestamp 1667941163
transform 1 0 30820 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_335
timestamp 1667941163
transform 1 0 31924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_347
timestamp 1667941163
transform 1 0 33028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_359
timestamp 1667941163
transform 1 0 34132 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_7
timestamp 1667941163
transform 1 0 1748 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_12
timestamp 1667941163
transform 1 0 2208 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_25
timestamp 1667941163
transform 1 0 3404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_29
timestamp 1667941163
transform 1 0 3772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_39
timestamp 1667941163
transform 1 0 4692 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1667941163
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_68
timestamp 1667941163
transform 1 0 7360 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_72
timestamp 1667941163
transform 1 0 7728 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_94
timestamp 1667941163
transform 1 0 9752 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_100
timestamp 1667941163
transform 1 0 10304 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1667941163
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_129
timestamp 1667941163
transform 1 0 12972 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_146
timestamp 1667941163
transform 1 0 14536 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_154
timestamp 1667941163
transform 1 0 15272 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1667941163
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1667941163
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_174
timestamp 1667941163
transform 1 0 17112 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1667941163
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1667941163
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_205
timestamp 1667941163
transform 1 0 19964 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_209
timestamp 1667941163
transform 1 0 20332 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_213
timestamp 1667941163
transform 1 0 20700 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_221
timestamp 1667941163
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_240
timestamp 1667941163
transform 1 0 23184 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_244
timestamp 1667941163
transform 1 0 23552 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_254
timestamp 1667941163
transform 1 0 24472 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1667941163
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1667941163
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1667941163
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_291
timestamp 1667941163
transform 1 0 27876 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_303
timestamp 1667941163
transform 1 0 28980 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_315
timestamp 1667941163
transform 1 0 30084 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_327
timestamp 1667941163
transform 1 0 31188 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_333
timestamp 1667941163
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_401
timestamp 1667941163
transform 1 0 37996 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_20
timestamp 1667941163
transform 1 0 2944 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_33
timestamp 1667941163
transform 1 0 4140 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_37
timestamp 1667941163
transform 1 0 4508 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_50
timestamp 1667941163
transform 1 0 5704 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_57
timestamp 1667941163
transform 1 0 6348 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_74
timestamp 1667941163
transform 1 0 7912 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_78
timestamp 1667941163
transform 1 0 8280 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1667941163
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_107
timestamp 1667941163
transform 1 0 10948 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_111
timestamp 1667941163
transform 1 0 11316 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_121
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1667941163
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_147
timestamp 1667941163
transform 1 0 14628 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_153
timestamp 1667941163
transform 1 0 15180 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_163
timestamp 1667941163
transform 1 0 16100 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_171
timestamp 1667941163
transform 1 0 16836 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_175
timestamp 1667941163
transform 1 0 17204 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_183
timestamp 1667941163
transform 1 0 17940 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1667941163
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1667941163
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1667941163
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_224
timestamp 1667941163
transform 1 0 21712 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_236
timestamp 1667941163
transform 1 0 22816 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_240
timestamp 1667941163
transform 1 0 23184 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1667941163
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_264
timestamp 1667941163
transform 1 0 25392 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_276
timestamp 1667941163
transform 1 0 26496 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_282
timestamp 1667941163
transform 1 0 27048 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_294
timestamp 1667941163
transform 1 0 28152 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1667941163
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1667941163
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_398
timestamp 1667941163
transform 1 0 37720 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_405
timestamp 1667941163
transform 1 0 38364 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_9
timestamp 1667941163
transform 1 0 1932 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_30
timestamp 1667941163
transform 1 0 3864 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_41
timestamp 1667941163
transform 1 0 4876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1667941163
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_62
timestamp 1667941163
transform 1 0 6808 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_79
timestamp 1667941163
transform 1 0 8372 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_103
timestamp 1667941163
transform 1 0 10580 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1667941163
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_124
timestamp 1667941163
transform 1 0 12512 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_130
timestamp 1667941163
transform 1 0 13064 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_134
timestamp 1667941163
transform 1 0 13432 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_151
timestamp 1667941163
transform 1 0 14996 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1667941163
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_180
timestamp 1667941163
transform 1 0 17664 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_199
timestamp 1667941163
transform 1 0 19412 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_206
timestamp 1667941163
transform 1 0 20056 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_218
timestamp 1667941163
transform 1 0 21160 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1667941163
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_249
timestamp 1667941163
transform 1 0 24012 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_253
timestamp 1667941163
transform 1 0 24380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_260
timestamp 1667941163
transform 1 0 25024 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_267
timestamp 1667941163
transform 1 0 25668 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_274
timestamp 1667941163
transform 1 0 26312 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1667941163
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1667941163
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1667941163
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1667941163
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_390
timestamp 1667941163
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_402
timestamp 1667941163
transform 1 0 38088 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_406
timestamp 1667941163
transform 1 0 38456 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_19
timestamp 1667941163
transform 1 0 2852 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1667941163
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_44
timestamp 1667941163
transform 1 0 5152 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_52
timestamp 1667941163
transform 1 0 5888 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_56
timestamp 1667941163
transform 1 0 6256 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_69
timestamp 1667941163
transform 1 0 7452 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1667941163
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_90
timestamp 1667941163
transform 1 0 9384 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_107
timestamp 1667941163
transform 1 0 10948 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_124
timestamp 1667941163
transform 1 0 12512 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_137
timestamp 1667941163
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_152
timestamp 1667941163
transform 1 0 15088 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_159
timestamp 1667941163
transform 1 0 15732 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_166
timestamp 1667941163
transform 1 0 16376 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_173
timestamp 1667941163
transform 1 0 17020 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_188
timestamp 1667941163
transform 1 0 18400 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_208
timestamp 1667941163
transform 1 0 20240 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_214
timestamp 1667941163
transform 1 0 20792 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_228
timestamp 1667941163
transform 1 0 22080 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_240
timestamp 1667941163
transform 1 0 23184 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_264
timestamp 1667941163
transform 1 0 25392 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_273
timestamp 1667941163
transform 1 0 26220 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_285
timestamp 1667941163
transform 1 0 27324 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_297
timestamp 1667941163
transform 1 0 28428 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_305
timestamp 1667941163
transform 1 0 29164 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_392
timestamp 1667941163
transform 1 0 37168 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_18
timestamp 1667941163
transform 1 0 2760 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_31
timestamp 1667941163
transform 1 0 3956 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_37
timestamp 1667941163
transform 1 0 4508 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_41
timestamp 1667941163
transform 1 0 4876 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1667941163
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_61
timestamp 1667941163
transform 1 0 6716 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_71
timestamp 1667941163
transform 1 0 7636 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_84
timestamp 1667941163
transform 1 0 8832 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_101
timestamp 1667941163
transform 1 0 10396 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1667941163
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_125
timestamp 1667941163
transform 1 0 12604 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_133
timestamp 1667941163
transform 1 0 13340 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_142
timestamp 1667941163
transform 1 0 14168 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_150
timestamp 1667941163
transform 1 0 14904 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1667941163
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_188
timestamp 1667941163
transform 1 0 18400 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_195
timestamp 1667941163
transform 1 0 19044 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_212
timestamp 1667941163
transform 1 0 20608 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_219
timestamp 1667941163
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1667941163
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_230
timestamp 1667941163
transform 1 0 22264 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_242
timestamp 1667941163
transform 1 0 23368 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_254
timestamp 1667941163
transform 1 0 24472 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_266
timestamp 1667941163
transform 1 0 25576 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1667941163
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_287
timestamp 1667941163
transform 1 0 27508 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_291
timestamp 1667941163
transform 1 0 27876 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_303
timestamp 1667941163
transform 1 0 28980 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_315
timestamp 1667941163
transform 1 0 30084 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_327
timestamp 1667941163
transform 1 0 31188 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_369
timestamp 1667941163
transform 1 0 35052 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_397
timestamp 1667941163
transform 1 0 37628 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_401
timestamp 1667941163
transform 1 0 37996 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_9
timestamp 1667941163
transform 1 0 1932 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_22
timestamp 1667941163
transform 1 0 3128 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_40
timestamp 1667941163
transform 1 0 4784 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_57
timestamp 1667941163
transform 1 0 6348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_61
timestamp 1667941163
transform 1 0 6716 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_74
timestamp 1667941163
transform 1 0 7912 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_78
timestamp 1667941163
transform 1 0 8280 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1667941163
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_89
timestamp 1667941163
transform 1 0 9292 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_93
timestamp 1667941163
transform 1 0 9660 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_110
timestamp 1667941163
transform 1 0 11224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_127
timestamp 1667941163
transform 1 0 12788 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1667941163
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_151
timestamp 1667941163
transform 1 0 14996 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_158
timestamp 1667941163
transform 1 0 15640 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_166
timestamp 1667941163
transform 1 0 16376 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_171
timestamp 1667941163
transform 1 0 16836 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_178
timestamp 1667941163
transform 1 0 17480 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_190
timestamp 1667941163
transform 1 0 18584 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_207
timestamp 1667941163
transform 1 0 20148 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_221
timestamp 1667941163
transform 1 0 21436 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_237
timestamp 1667941163
transform 1 0 22908 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_249
timestamp 1667941163
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_274
timestamp 1667941163
transform 1 0 26312 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_286
timestamp 1667941163
transform 1 0 27416 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_298
timestamp 1667941163
transform 1 0 28520 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_306
timestamp 1667941163
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_327
timestamp 1667941163
transform 1 0 31188 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_331
timestamp 1667941163
transform 1 0 31556 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_343
timestamp 1667941163
transform 1 0 32660 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_355
timestamp 1667941163
transform 1 0 33764 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_393
timestamp 1667941163
transform 1 0 37260 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_397
timestamp 1667941163
transform 1 0 37628 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_405
timestamp 1667941163
transform 1 0 38364 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_15
timestamp 1667941163
transform 1 0 2484 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_32
timestamp 1667941163
transform 1 0 4048 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_45
timestamp 1667941163
transform 1 0 5244 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1667941163
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_72
timestamp 1667941163
transform 1 0 7728 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_80
timestamp 1667941163
transform 1 0 8464 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_90
timestamp 1667941163
transform 1 0 9384 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_103
timestamp 1667941163
transform 1 0 10580 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1667941163
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_119
timestamp 1667941163
transform 1 0 12052 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_126
timestamp 1667941163
transform 1 0 12696 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_133
timestamp 1667941163
transform 1 0 13340 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_140
timestamp 1667941163
transform 1 0 13984 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_144
timestamp 1667941163
transform 1 0 14352 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_154
timestamp 1667941163
transform 1 0 15272 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1667941163
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1667941163
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_190
timestamp 1667941163
transform 1 0 18584 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_202
timestamp 1667941163
transform 1 0 19688 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_214
timestamp 1667941163
transform 1 0 20792 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1667941163
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_240
timestamp 1667941163
transform 1 0 23184 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_248
timestamp 1667941163
transform 1 0 23920 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_257
timestamp 1667941163
transform 1 0 24748 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_266
timestamp 1667941163
transform 1 0 25576 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1667941163
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_289
timestamp 1667941163
transform 1 0 27692 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_299
timestamp 1667941163
transform 1 0 28612 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_303
timestamp 1667941163
transform 1 0 28980 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_315
timestamp 1667941163
transform 1 0 30084 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_327
timestamp 1667941163
transform 1 0 31188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_342
timestamp 1667941163
transform 1 0 32568 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_354
timestamp 1667941163
transform 1 0 33672 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_366
timestamp 1667941163
transform 1 0 34776 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_378
timestamp 1667941163
transform 1 0 35880 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_390
timestamp 1667941163
transform 1 0 36984 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_9
timestamp 1667941163
transform 1 0 1932 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_22
timestamp 1667941163
transform 1 0 3128 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_33
timestamp 1667941163
transform 1 0 4140 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_37
timestamp 1667941163
transform 1 0 4508 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_50
timestamp 1667941163
transform 1 0 5704 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_58
timestamp 1667941163
transform 1 0 6440 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_69
timestamp 1667941163
transform 1 0 7452 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_77
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1667941163
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_98
timestamp 1667941163
transform 1 0 10120 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_102
timestamp 1667941163
transform 1 0 10488 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_116
timestamp 1667941163
transform 1 0 11776 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_120
timestamp 1667941163
transform 1 0 12144 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_134
timestamp 1667941163
transform 1 0 13432 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_145
timestamp 1667941163
transform 1 0 14444 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_149
timestamp 1667941163
transform 1 0 14812 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_156
timestamp 1667941163
transform 1 0 15456 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_168
timestamp 1667941163
transform 1 0 16560 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_180
timestamp 1667941163
transform 1 0 17664 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1667941163
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1667941163
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_221
timestamp 1667941163
transform 1 0 21436 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_225
timestamp 1667941163
transform 1 0 21804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_229
timestamp 1667941163
transform 1 0 22172 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_237
timestamp 1667941163
transform 1 0 22908 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_243
timestamp 1667941163
transform 1 0 23460 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1667941163
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1667941163
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_397
timestamp 1667941163
transform 1 0 37628 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_402
timestamp 1667941163
transform 1 0 38088 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_406
timestamp 1667941163
transform 1 0 38456 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_14
timestamp 1667941163
transform 1 0 2392 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_27
timestamp 1667941163
transform 1 0 3588 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_35
timestamp 1667941163
transform 1 0 4324 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_40
timestamp 1667941163
transform 1 0 4784 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_47
timestamp 1667941163
transform 1 0 5428 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1667941163
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_64
timestamp 1667941163
transform 1 0 6992 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_89
timestamp 1667941163
transform 1 0 9292 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1667941163
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_119
timestamp 1667941163
transform 1 0 12052 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_129
timestamp 1667941163
transform 1 0 12972 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_140
timestamp 1667941163
transform 1 0 13984 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_152
timestamp 1667941163
transform 1 0 15088 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1667941163
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_181
timestamp 1667941163
transform 1 0 17756 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_185
timestamp 1667941163
transform 1 0 18124 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_202
timestamp 1667941163
transform 1 0 19688 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_214
timestamp 1667941163
transform 1 0 20792 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_221
timestamp 1667941163
transform 1 0 21436 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_240
timestamp 1667941163
transform 1 0 23184 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_244
timestamp 1667941163
transform 1 0 23552 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_248
timestamp 1667941163
transform 1 0 23920 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_254
timestamp 1667941163
transform 1 0 24472 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_258
timestamp 1667941163
transform 1 0 24840 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_270
timestamp 1667941163
transform 1 0 25944 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1667941163
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1667941163
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1667941163
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_36
timestamp 1667941163
transform 1 0 4416 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_43
timestamp 1667941163
transform 1 0 5060 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_55
timestamp 1667941163
transform 1 0 6164 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_63
timestamp 1667941163
transform 1 0 6900 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_68
timestamp 1667941163
transform 1 0 7360 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_75
timestamp 1667941163
transform 1 0 8004 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1667941163
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_89
timestamp 1667941163
transform 1 0 9292 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_103
timestamp 1667941163
transform 1 0 10580 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_107
timestamp 1667941163
transform 1 0 10948 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_111
timestamp 1667941163
transform 1 0 11316 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_115
timestamp 1667941163
transform 1 0 11684 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_119
timestamp 1667941163
transform 1 0 12052 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1667941163
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_152
timestamp 1667941163
transform 1 0 15088 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_159
timestamp 1667941163
transform 1 0 15732 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_171
timestamp 1667941163
transform 1 0 16836 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_183
timestamp 1667941163
transform 1 0 17940 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_190
timestamp 1667941163
transform 1 0 18584 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1667941163
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1667941163
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1667941163
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1667941163
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1667941163
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_258
timestamp 1667941163
transform 1 0 24840 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_283
timestamp 1667941163
transform 1 0 27140 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_287
timestamp 1667941163
transform 1 0 27508 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_299
timestamp 1667941163
transform 1 0 28612 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_9
timestamp 1667941163
transform 1 0 1932 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_15
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_19
timestamp 1667941163
transform 1 0 2852 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_26
timestamp 1667941163
transform 1 0 3496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_33
timestamp 1667941163
transform 1 0 4140 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_40
timestamp 1667941163
transform 1 0 4784 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_47
timestamp 1667941163
transform 1 0 5428 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1667941163
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_62
timestamp 1667941163
transform 1 0 6808 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_71
timestamp 1667941163
transform 1 0 7636 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_85
timestamp 1667941163
transform 1 0 8924 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_97
timestamp 1667941163
transform 1 0 10028 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_101
timestamp 1667941163
transform 1 0 10396 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1667941163
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1667941163
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_118
timestamp 1667941163
transform 1 0 11960 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_130
timestamp 1667941163
transform 1 0 13064 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_135
timestamp 1667941163
transform 1 0 13524 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_142
timestamp 1667941163
transform 1 0 14168 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_149
timestamp 1667941163
transform 1 0 14812 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_153
timestamp 1667941163
transform 1 0 15180 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_163
timestamp 1667941163
transform 1 0 16100 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1667941163
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_186
timestamp 1667941163
transform 1 0 18216 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1667941163
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1667941163
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1667941163
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_230
timestamp 1667941163
transform 1 0 22264 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_238
timestamp 1667941163
transform 1 0 23000 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_249
timestamp 1667941163
transform 1 0 24012 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_253
timestamp 1667941163
transform 1 0 24380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_257
timestamp 1667941163
transform 1 0 24748 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_269
timestamp 1667941163
transform 1 0 25852 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1667941163
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1667941163
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1667941163
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_346
timestamp 1667941163
transform 1 0 32936 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_358
timestamp 1667941163
transform 1 0 34040 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_370
timestamp 1667941163
transform 1 0 35144 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_382
timestamp 1667941163
transform 1 0 36248 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_390
timestamp 1667941163
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_9
timestamp 1667941163
transform 1 0 1932 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_18
timestamp 1667941163
transform 1 0 2760 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_25
timestamp 1667941163
transform 1 0 3404 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1667941163
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_48
timestamp 1667941163
transform 1 0 5520 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_55
timestamp 1667941163
transform 1 0 6164 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_72
timestamp 1667941163
transform 1 0 7728 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_80
timestamp 1667941163
transform 1 0 8464 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_90
timestamp 1667941163
transform 1 0 9384 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_96
timestamp 1667941163
transform 1 0 9936 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_100
timestamp 1667941163
transform 1 0 10304 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_111
timestamp 1667941163
transform 1 0 11316 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_123
timestamp 1667941163
transform 1 0 12420 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_135
timestamp 1667941163
transform 1 0 13524 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1667941163
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_152
timestamp 1667941163
transform 1 0 15088 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_161
timestamp 1667941163
transform 1 0 15916 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_174
timestamp 1667941163
transform 1 0 17112 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_181
timestamp 1667941163
transform 1 0 17756 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1667941163
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_202
timestamp 1667941163
transform 1 0 19688 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_211
timestamp 1667941163
transform 1 0 20516 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_223
timestamp 1667941163
transform 1 0 21620 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_235
timestamp 1667941163
transform 1 0 22724 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1667941163
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1667941163
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1667941163
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_328
timestamp 1667941163
transform 1 0 31280 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_340
timestamp 1667941163
transform 1 0 32384 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_352
timestamp 1667941163
transform 1 0 33488 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1667941163
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_10
timestamp 1667941163
transform 1 0 2024 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_14
timestamp 1667941163
transform 1 0 2392 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_18
timestamp 1667941163
transform 1 0 2760 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_27
timestamp 1667941163
transform 1 0 3588 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_34
timestamp 1667941163
transform 1 0 4232 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_41
timestamp 1667941163
transform 1 0 4876 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_48
timestamp 1667941163
transform 1 0 5520 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_63
timestamp 1667941163
transform 1 0 6900 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_67
timestamp 1667941163
transform 1 0 7268 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_83
timestamp 1667941163
transform 1 0 8740 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_90
timestamp 1667941163
transform 1 0 9384 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_94
timestamp 1667941163
transform 1 0 9752 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_98
timestamp 1667941163
transform 1 0 10120 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1667941163
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_131
timestamp 1667941163
transform 1 0 13156 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_145
timestamp 1667941163
transform 1 0 14444 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_160
timestamp 1667941163
transform 1 0 15824 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_174
timestamp 1667941163
transform 1 0 17112 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_180
timestamp 1667941163
transform 1 0 17664 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_194
timestamp 1667941163
transform 1 0 18952 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_206
timestamp 1667941163
transform 1 0 20056 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_218
timestamp 1667941163
transform 1 0 21160 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1667941163
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1667941163
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1667941163
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1667941163
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1667941163
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1667941163
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1667941163
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_9
timestamp 1667941163
transform 1 0 1932 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_16
timestamp 1667941163
transform 1 0 2576 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_23
timestamp 1667941163
transform 1 0 3220 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_40
timestamp 1667941163
transform 1 0 4784 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_49
timestamp 1667941163
transform 1 0 5612 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_61
timestamp 1667941163
transform 1 0 6716 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_68
timestamp 1667941163
transform 1 0 7360 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_79
timestamp 1667941163
transform 1 0 8372 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_90
timestamp 1667941163
transform 1 0 9384 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_102
timestamp 1667941163
transform 1 0 10488 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_107
timestamp 1667941163
transform 1 0 10948 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_119
timestamp 1667941163
transform 1 0 12052 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_124
timestamp 1667941163
transform 1 0 12512 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_137
timestamp 1667941163
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_146
timestamp 1667941163
transform 1 0 14536 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_153
timestamp 1667941163
transform 1 0 15180 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_160
timestamp 1667941163
transform 1 0 15824 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_173
timestamp 1667941163
transform 1 0 17020 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_185
timestamp 1667941163
transform 1 0 18124 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1667941163
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_208
timestamp 1667941163
transform 1 0 20240 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_220
timestamp 1667941163
transform 1 0 21344 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_224
timestamp 1667941163
transform 1 0 21712 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_236
timestamp 1667941163
transform 1 0 22816 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1667941163
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1667941163
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1667941163
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_316
timestamp 1667941163
transform 1 0 30176 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_328
timestamp 1667941163
transform 1 0 31280 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_340
timestamp 1667941163
transform 1 0 32384 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_352
timestamp 1667941163
transform 1 0 33488 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_401
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_14
timestamp 1667941163
transform 1 0 2392 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_22
timestamp 1667941163
transform 1 0 3128 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_26
timestamp 1667941163
transform 1 0 3496 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_32
timestamp 1667941163
transform 1 0 4048 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_36
timestamp 1667941163
transform 1 0 4416 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_43
timestamp 1667941163
transform 1 0 5060 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1667941163
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_62
timestamp 1667941163
transform 1 0 6808 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_70
timestamp 1667941163
transform 1 0 7544 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_75
timestamp 1667941163
transform 1 0 8004 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_87
timestamp 1667941163
transform 1 0 9108 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_101
timestamp 1667941163
transform 1 0 10396 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp 1667941163
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_125
timestamp 1667941163
transform 1 0 12604 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_136
timestamp 1667941163
transform 1 0 13616 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_143
timestamp 1667941163
transform 1 0 14260 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_150
timestamp 1667941163
transform 1 0 14904 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_157
timestamp 1667941163
transform 1 0 15548 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_165
timestamp 1667941163
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_174
timestamp 1667941163
transform 1 0 17112 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_189
timestamp 1667941163
transform 1 0 18492 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_201
timestamp 1667941163
transform 1 0 19596 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_213
timestamp 1667941163
transform 1 0 20700 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_221
timestamp 1667941163
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1667941163
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1667941163
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1667941163
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1667941163
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_7
timestamp 1667941163
transform 1 0 1748 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_11
timestamp 1667941163
transform 1 0 2116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_18
timestamp 1667941163
transform 1 0 2760 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_25
timestamp 1667941163
transform 1 0 3404 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_35
timestamp 1667941163
transform 1 0 4324 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_43
timestamp 1667941163
transform 1 0 5060 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_47
timestamp 1667941163
transform 1 0 5428 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_54
timestamp 1667941163
transform 1 0 6072 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_62
timestamp 1667941163
transform 1 0 6808 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_66
timestamp 1667941163
transform 1 0 7176 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_70
timestamp 1667941163
transform 1 0 7544 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_79
timestamp 1667941163
transform 1 0 8372 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_117
timestamp 1667941163
transform 1 0 11868 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_127
timestamp 1667941163
transform 1 0 12788 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_134
timestamp 1667941163
transform 1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_147
timestamp 1667941163
transform 1 0 14628 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_159
timestamp 1667941163
transform 1 0 15732 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_164
timestamp 1667941163
transform 1 0 16192 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_171
timestamp 1667941163
transform 1 0 16836 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_179
timestamp 1667941163
transform 1 0 17572 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_184
timestamp 1667941163
transform 1 0 18032 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_209
timestamp 1667941163
transform 1 0 20332 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_224
timestamp 1667941163
transform 1 0 21712 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_236
timestamp 1667941163
transform 1 0 22816 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1667941163
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1667941163
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1667941163
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1667941163
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_401
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_405
timestamp 1667941163
transform 1 0 38364 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_7
timestamp 1667941163
transform 1 0 1748 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_11
timestamp 1667941163
transform 1 0 2116 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_18
timestamp 1667941163
transform 1 0 2760 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_25
timestamp 1667941163
transform 1 0 3404 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_32
timestamp 1667941163
transform 1 0 4048 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_39
timestamp 1667941163
transform 1 0 4692 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_43
timestamp 1667941163
transform 1 0 5060 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_47
timestamp 1667941163
transform 1 0 5428 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_68
timestamp 1667941163
transform 1 0 7360 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_80
timestamp 1667941163
transform 1 0 8464 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_92
timestamp 1667941163
transform 1 0 9568 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_104
timestamp 1667941163
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_120
timestamp 1667941163
transform 1 0 12144 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_133
timestamp 1667941163
transform 1 0 13340 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_145
timestamp 1667941163
transform 1 0 14444 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_157
timestamp 1667941163
transform 1 0 15548 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_165
timestamp 1667941163
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_180
timestamp 1667941163
transform 1 0 17664 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_200
timestamp 1667941163
transform 1 0 19504 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_212
timestamp 1667941163
transform 1 0 20608 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1667941163
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_398
timestamp 1667941163
transform 1 0 37720 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_406
timestamp 1667941163
transform 1 0 38456 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_7
timestamp 1667941163
transform 1 0 1748 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_11
timestamp 1667941163
transform 1 0 2116 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_18
timestamp 1667941163
transform 1 0 2760 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_25
timestamp 1667941163
transform 1 0 3404 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_34
timestamp 1667941163
transform 1 0 4232 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_46
timestamp 1667941163
transform 1 0 5336 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_58
timestamp 1667941163
transform 1 0 6440 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_70
timestamp 1667941163
transform 1 0 7544 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_75
timestamp 1667941163
transform 1 0 8004 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_93
timestamp 1667941163
transform 1 0 9660 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1667941163
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_121
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_130
timestamp 1667941163
transform 1 0 13064 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1667941163
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1667941163
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_165
timestamp 1667941163
transform 1 0 16284 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_171
timestamp 1667941163
transform 1 0 16836 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_180
timestamp 1667941163
transform 1 0 17664 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_187
timestamp 1667941163
transform 1 0 18308 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1667941163
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_202
timestamp 1667941163
transform 1 0 19688 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_214
timestamp 1667941163
transform 1 0 20792 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_226
timestamp 1667941163
transform 1 0 21896 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_231
timestamp 1667941163
transform 1 0 22356 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_243
timestamp 1667941163
transform 1 0 23460 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1667941163
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_393
timestamp 1667941163
transform 1 0 37260 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_397
timestamp 1667941163
transform 1 0 37628 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_405
timestamp 1667941163
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_12
timestamp 1667941163
transform 1 0 2208 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_19
timestamp 1667941163
transform 1 0 2852 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_26
timestamp 1667941163
transform 1 0 3496 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_33
timestamp 1667941163
transform 1 0 4140 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_45
timestamp 1667941163
transform 1 0 5244 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_49
timestamp 1667941163
transform 1 0 5612 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_53
timestamp 1667941163
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_75
timestamp 1667941163
transform 1 0 8004 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_79
timestamp 1667941163
transform 1 0 8372 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_86
timestamp 1667941163
transform 1 0 9016 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_98
timestamp 1667941163
transform 1 0 10120 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_109
timestamp 1667941163
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_128
timestamp 1667941163
transform 1 0 12880 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_140
timestamp 1667941163
transform 1 0 13984 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_152
timestamp 1667941163
transform 1 0 15088 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1667941163
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_175
timestamp 1667941163
transform 1 0 17204 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_179
timestamp 1667941163
transform 1 0 17572 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_183
timestamp 1667941163
transform 1 0 17940 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_198
timestamp 1667941163
transform 1 0 19320 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_210
timestamp 1667941163
transform 1 0 20424 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_218
timestamp 1667941163
transform 1 0 21160 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1667941163
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1667941163
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1667941163
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1667941163
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1667941163
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1667941163
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_7
timestamp 1667941163
transform 1 0 1748 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_11
timestamp 1667941163
transform 1 0 2116 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_18
timestamp 1667941163
transform 1 0 2760 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_26
timestamp 1667941163
transform 1 0 3496 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1667941163
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1667941163
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_161
timestamp 1667941163
transform 1 0 15916 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_167
timestamp 1667941163
transform 1 0 16468 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_179
timestamp 1667941163
transform 1 0 17572 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_191
timestamp 1667941163
transform 1 0 18676 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1667941163
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1667941163
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1667941163
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1667941163
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1667941163
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1667941163
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_8
timestamp 1667941163
transform 1 0 1840 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_20
timestamp 1667941163
transform 1 0 2944 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_32
timestamp 1667941163
transform 1 0 4048 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_44
timestamp 1667941163
transform 1 0 5152 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_75
timestamp 1667941163
transform 1 0 8004 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_79
timestamp 1667941163
transform 1 0 8372 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_91
timestamp 1667941163
transform 1 0 9476 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_103
timestamp 1667941163
transform 1 0 10580 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_118
timestamp 1667941163
transform 1 0 11960 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_130
timestamp 1667941163
transform 1 0 13064 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_142
timestamp 1667941163
transform 1 0 14168 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_154
timestamp 1667941163
transform 1 0 15272 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1667941163
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_174
timestamp 1667941163
transform 1 0 17112 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1667941163
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1667941163
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1667941163
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_8
timestamp 1667941163
transform 1 0 1840 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_20
timestamp 1667941163
transform 1 0 2944 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_44
timestamp 1667941163
transform 1 0 5152 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_56
timestamp 1667941163
transform 1 0 6256 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_68
timestamp 1667941163
transform 1 0 7360 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_80
timestamp 1667941163
transform 1 0 8464 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_90
timestamp 1667941163
transform 1 0 9384 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_102
timestamp 1667941163
transform 1 0 10488 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_117
timestamp 1667941163
transform 1 0 11868 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_129
timestamp 1667941163
transform 1 0 12972 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_137
timestamp 1667941163
transform 1 0 13708 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_177
timestamp 1667941163
transform 1 0 17388 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_183
timestamp 1667941163
transform 1 0 17940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1667941163
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1667941163
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1667941163
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1667941163
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_277
timestamp 1667941163
transform 1 0 26588 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_288
timestamp 1667941163
transform 1 0 27600 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_300
timestamp 1667941163
transform 1 0 28704 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_405
timestamp 1667941163
transform 1 0 38364 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_9
timestamp 1667941163
transform 1 0 1932 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_21
timestamp 1667941163
transform 1 0 3036 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_33
timestamp 1667941163
transform 1 0 4140 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_38
timestamp 1667941163
transform 1 0 4600 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_50
timestamp 1667941163
transform 1 0 5704 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1667941163
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1667941163
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1667941163
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1667941163
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1667941163
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1667941163
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1667941163
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1667941163
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1667941163
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1667941163
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1667941163
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1667941163
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1667941163
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1667941163
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1667941163
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1667941163
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_34
timestamp 1667941163
transform 1 0 4232 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_46
timestamp 1667941163
transform 1 0 5336 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_50
timestamp 1667941163
transform 1 0 5704 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_54
timestamp 1667941163
transform 1 0 6072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_61
timestamp 1667941163
transform 1 0 6716 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_68
timestamp 1667941163
transform 1 0 7360 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_76
timestamp 1667941163
transform 1 0 8096 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_81
timestamp 1667941163
transform 1 0 8556 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_96
timestamp 1667941163
transform 1 0 9936 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_108
timestamp 1667941163
transform 1 0 11040 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_120
timestamp 1667941163
transform 1 0 12144 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_131
timestamp 1667941163
transform 1 0 13156 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1667941163
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1667941163
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1667941163
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_269
timestamp 1667941163
transform 1 0 25852 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_273
timestamp 1667941163
transform 1 0 26220 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_285
timestamp 1667941163
transform 1 0 27324 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_291
timestamp 1667941163
transform 1 0 27876 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_295
timestamp 1667941163
transform 1 0 28244 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_389
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_405
timestamp 1667941163
transform 1 0 38364 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1667941163
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1667941163
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1667941163
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1667941163
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1667941163
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_309
timestamp 1667941163
transform 1 0 29532 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_321
timestamp 1667941163
transform 1 0 30636 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_333
timestamp 1667941163
transform 1 0 31740 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1667941163
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1667941163
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1667941163
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_217
timestamp 1667941163
transform 1 0 21068 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_223
timestamp 1667941163
transform 1 0 21620 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_235
timestamp 1667941163
transform 1 0 22724 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_247
timestamp 1667941163
transform 1 0 23828 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_258
timestamp 1667941163
transform 1 0 24840 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_270
timestamp 1667941163
transform 1 0 25944 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_282
timestamp 1667941163
transform 1 0 27048 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_290
timestamp 1667941163
transform 1 0 27784 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_295
timestamp 1667941163
transform 1 0 28244 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_9
timestamp 1667941163
transform 1 0 1932 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_13
timestamp 1667941163
transform 1 0 2300 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_25
timestamp 1667941163
transform 1 0 3404 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_37
timestamp 1667941163
transform 1 0 4508 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_49
timestamp 1667941163
transform 1 0 5612 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1667941163
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_85
timestamp 1667941163
transform 1 0 8924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_89
timestamp 1667941163
transform 1 0 9292 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_101
timestamp 1667941163
transform 1 0 10396 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_106
timestamp 1667941163
transform 1 0 10856 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_55_216
timestamp 1667941163
transform 1 0 20976 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_246
timestamp 1667941163
transform 1 0 23736 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_258
timestamp 1667941163
transform 1 0 24840 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_270
timestamp 1667941163
transform 1 0 25944 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 1667941163
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1667941163
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_91
timestamp 1667941163
transform 1 0 9476 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_95
timestamp 1667941163
transform 1 0 9844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_107
timestamp 1667941163
transform 1 0 10948 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_111
timestamp 1667941163
transform 1 0 11316 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_123
timestamp 1667941163
transform 1 0 12420 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_135
timestamp 1667941163
transform 1 0 13524 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_56_298
timestamp 1667941163
transform 1 0 28520 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_306
timestamp 1667941163
transform 1 0 29256 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_352
timestamp 1667941163
transform 1 0 33488 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_405
timestamp 1667941163
transform 1 0 38364 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_9
timestamp 1667941163
transform 1 0 1932 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_21
timestamp 1667941163
transform 1 0 3036 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_33
timestamp 1667941163
transform 1 0 4140 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_45
timestamp 1667941163
transform 1 0 5244 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_53
timestamp 1667941163
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_84
timestamp 1667941163
transform 1 0 8832 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_96
timestamp 1667941163
transform 1 0 9936 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_108
timestamp 1667941163
transform 1 0 11040 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_230
timestamp 1667941163
transform 1 0 22264 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_242
timestamp 1667941163
transform 1 0 23368 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 1667941163
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1667941163
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_27
timestamp 1667941163
transform 1 0 3588 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_38
timestamp 1667941163
transform 1 0 4600 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_50
timestamp 1667941163
transform 1 0 5704 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_8
timestamp 1667941163
transform 1 0 1840 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_20
timestamp 1667941163
transform 1 0 2944 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_25
timestamp 1667941163
transform 1 0 3404 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_202
timestamp 1667941163
transform 1 0 19688 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_214
timestamp 1667941163
transform 1 0 20792 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_226
timestamp 1667941163
transform 1 0 21896 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_238
timestamp 1667941163
transform 1 0 23000 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1667941163
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_401
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_405
timestamp 1667941163
transform 1 0 38364 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1667941163
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1667941163
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1667941163
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1667941163
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_8
timestamp 1667941163
transform 1 0 1840 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_20
timestamp 1667941163
transform 1 0 2944 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_201
timestamp 1667941163
transform 1 0 19596 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_205
timestamp 1667941163
transform 1 0 19964 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_217
timestamp 1667941163
transform 1 0 21068 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_229
timestamp 1667941163
transform 1 0 22172 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_241
timestamp 1667941163
transform 1 0 23276 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_249
timestamp 1667941163
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_397
timestamp 1667941163
transform 1 0 37628 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_16
timestamp 1667941163
transform 1 0 2576 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_23
timestamp 1667941163
transform 1 0 3220 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_35
timestamp 1667941163
transform 1 0 4324 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_47
timestamp 1667941163
transform 1 0 5428 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1667941163
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_91
timestamp 1667941163
transform 1 0 9476 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_103
timestamp 1667941163
transform 1 0 10580 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_137
timestamp 1667941163
transform 1 0 13708 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_144
timestamp 1667941163
transform 1 0 14352 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_148
timestamp 1667941163
transform 1 0 14720 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_152
timestamp 1667941163
transform 1 0 15088 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_164
timestamp 1667941163
transform 1 0 16192 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_175
timestamp 1667941163
transform 1 0 17204 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_179
timestamp 1667941163
transform 1 0 17572 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_183
timestamp 1667941163
transform 1 0 17940 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_195
timestamp 1667941163
transform 1 0 19044 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_207
timestamp 1667941163
transform 1 0 20148 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_219
timestamp 1667941163
transform 1 0 21252 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_230
timestamp 1667941163
transform 1 0 22264 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_238
timestamp 1667941163
transform 1 0 23000 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_251
timestamp 1667941163
transform 1 0 24196 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_263
timestamp 1667941163
transform 1 0 25300 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_275
timestamp 1667941163
transform 1 0 26404 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1667941163
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_286
timestamp 1667941163
transform 1 0 27416 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_298
timestamp 1667941163
transform 1 0 28520 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_310
timestamp 1667941163
transform 1 0 29624 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_322
timestamp 1667941163
transform 1 0 30728 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_334
timestamp 1667941163
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_373
timestamp 1667941163
transform 1 0 35420 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_377
timestamp 1667941163
transform 1 0 35788 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_385
timestamp 1667941163
transform 1 0 36524 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1667941163
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_9
timestamp 1667941163
transform 1 0 1932 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_20
timestamp 1667941163
transform 1 0 2944 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_35
timestamp 1667941163
transform 1 0 4324 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_42
timestamp 1667941163
transform 1 0 4968 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_50
timestamp 1667941163
transform 1 0 5704 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_54
timestamp 1667941163
transform 1 0 6072 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_62
timestamp 1667941163
transform 1 0 6808 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_70
timestamp 1667941163
transform 1 0 7544 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1667941163
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1667941163
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_93
timestamp 1667941163
transform 1 0 9660 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_98
timestamp 1667941163
transform 1 0 10120 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_110
timestamp 1667941163
transform 1 0 11224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_119
timestamp 1667941163
transform 1 0 12052 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_126
timestamp 1667941163
transform 1 0 12696 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_134
timestamp 1667941163
transform 1 0 13432 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1667941163
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_147
timestamp 1667941163
transform 1 0 14628 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_155
timestamp 1667941163
transform 1 0 15364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_161
timestamp 1667941163
transform 1 0 15916 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 1667941163
transform 1 0 16468 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_177
timestamp 1667941163
transform 1 0 17388 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_182
timestamp 1667941163
transform 1 0 17848 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_194
timestamp 1667941163
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_205
timestamp 1667941163
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_210
timestamp 1667941163
transform 1 0 20424 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1667941163
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_237
timestamp 1667941163
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 1667941163
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_259
timestamp 1667941163
transform 1 0 24932 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_266
timestamp 1667941163
transform 1 0 25576 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_278
timestamp 1667941163
transform 1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_287
timestamp 1667941163
transform 1 0 27508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_295
timestamp 1667941163
transform 1 0 28244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_302
timestamp 1667941163
transform 1 0 28888 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_314
timestamp 1667941163
transform 1 0 29992 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_322
timestamp 1667941163
transform 1 0 30728 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_328
timestamp 1667941163
transform 1 0 31280 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_343
timestamp 1667941163
transform 1 0 32660 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_351
timestamp 1667941163
transform 1 0 33396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1667941163
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_371
timestamp 1667941163
transform 1 0 35236 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_375
timestamp 1667941163
transform 1 0 35604 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_379
timestamp 1667941163
transform 1 0 35972 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_385
timestamp 1667941163
transform 1 0 36524 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_391
timestamp 1667941163
transform 1 0 37076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_399
timestamp 1667941163
transform 1 0 37812 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0383_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4508 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0384_
timestamp 1667941163
transform 1 0 9936 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0385_
timestamp 1667941163
transform 1 0 16100 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0386_
timestamp 1667941163
transform 1 0 19688 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0387_
timestamp 1667941163
transform 1 0 7728 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0388_
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0389_
timestamp 1667941163
transform 1 0 8372 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0390_
timestamp 1667941163
transform 1 0 21160 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0391_
timestamp 1667941163
transform 1 0 21436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0392_
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0393_
timestamp 1667941163
transform 1 0 6624 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0394_
timestamp 1667941163
transform 1 0 16100 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0395_
timestamp 1667941163
transform 1 0 5796 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0396_
timestamp 1667941163
transform 1 0 12880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0397_
timestamp 1667941163
transform 1 0 24564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0398_
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0399_
timestamp 1667941163
transform 1 0 24840 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0400_
timestamp 1667941163
transform 1 0 4508 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0401_
timestamp 1667941163
transform 1 0 4140 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0402_
timestamp 1667941163
transform 1 0 2576 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0403_
timestamp 1667941163
transform 1 0 9108 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0404_
timestamp 1667941163
transform 1 0 13524 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0405_
timestamp 1667941163
transform 1 0 23460 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0406_
timestamp 1667941163
transform 1 0 15180 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0407_
timestamp 1667941163
transform 1 0 23368 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0408_
timestamp 1667941163
transform 1 0 27140 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0409_
timestamp 1667941163
transform 1 0 24472 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0410_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 25208 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0411_
timestamp 1667941163
transform 1 0 24564 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0412_
timestamp 1667941163
transform 1 0 28244 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0413_
timestamp 1667941163
transform 1 0 27876 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0414_
timestamp 1667941163
transform 1 0 26772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0415_
timestamp 1667941163
transform 1 0 27784 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0416_
timestamp 1667941163
transform 1 0 27600 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0417_
timestamp 1667941163
transform 1 0 11868 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0418_
timestamp 1667941163
transform 1 0 16192 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0419_
timestamp 1667941163
transform 1 0 11592 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0420_
timestamp 1667941163
transform 1 0 11684 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0421_
timestamp 1667941163
transform 1 0 13156 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0422_
timestamp 1667941163
transform 1 0 12788 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0423_
timestamp 1667941163
transform 1 0 18032 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0424_
timestamp 1667941163
transform 1 0 17664 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0425_
timestamp 1667941163
transform 1 0 17480 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0426_
timestamp 1667941163
transform 1 0 26864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0427_
timestamp 1667941163
transform 1 0 25300 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0428_
timestamp 1667941163
transform 1 0 21896 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0429_
timestamp 1667941163
transform 1 0 21988 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0430_
timestamp 1667941163
transform 1 0 28152 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0431_
timestamp 1667941163
transform 1 0 27508 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0432_
timestamp 1667941163
transform 1 0 27048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0433_
timestamp 1667941163
transform 1 0 27600 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0434_
timestamp 1667941163
transform 1 0 27784 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0435_
timestamp 1667941163
transform 1 0 5612 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0436_
timestamp 1667941163
transform 1 0 5796 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0437_
timestamp 1667941163
transform 1 0 10672 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0438_
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0439_
timestamp 1667941163
transform 1 0 5336 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0440_
timestamp 1667941163
transform 1 0 9108 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0441_
timestamp 1667941163
transform 1 0 15456 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0442_
timestamp 1667941163
transform 1 0 16836 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0443_
timestamp 1667941163
transform 1 0 14904 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0444_
timestamp 1667941163
transform 1 0 17664 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0445_
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0446_
timestamp 1667941163
transform 1 0 9752 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0447_
timestamp 1667941163
transform 1 0 9844 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0448_
timestamp 1667941163
transform 1 0 18676 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0449_
timestamp 1667941163
transform 1 0 19044 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0450_
timestamp 1667941163
transform 1 0 24104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0451_
timestamp 1667941163
transform 1 0 8372 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0452_
timestamp 1667941163
transform 1 0 9384 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0453_
timestamp 1667941163
transform 1 0 15640 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0454_
timestamp 1667941163
transform 1 0 26036 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0455_
timestamp 1667941163
transform 1 0 25392 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0456_
timestamp 1667941163
transform 1 0 15548 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0457_
timestamp 1667941163
transform 1 0 13708 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0458_
timestamp 1667941163
transform 1 0 13064 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0459_
timestamp 1667941163
transform 1 0 13524 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0460_
timestamp 1667941163
transform 1 0 15916 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0461_
timestamp 1667941163
transform 1 0 16560 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0462_
timestamp 1667941163
transform 1 0 13984 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0463_
timestamp 1667941163
transform 1 0 21252 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0464_
timestamp 1667941163
transform 1 0 21988 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0465_
timestamp 1667941163
transform 1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0466_
timestamp 1667941163
transform 1 0 13340 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0467_
timestamp 1667941163
transform 1 0 15272 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0468_
timestamp 1667941163
transform 1 0 7728 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0469_
timestamp 1667941163
transform 1 0 11684 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0470_
timestamp 1667941163
transform 1 0 13892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0471_
timestamp 1667941163
transform 1 0 15640 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0472_
timestamp 1667941163
transform 1 0 8096 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0473_
timestamp 1667941163
transform 1 0 8740 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0474_
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0475_
timestamp 1667941163
transform 1 0 20608 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0476_
timestamp 1667941163
transform 1 0 19320 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0477_
timestamp 1667941163
transform 1 0 18676 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0478_
timestamp 1667941163
transform 1 0 24564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0479_
timestamp 1667941163
transform 1 0 23736 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0480_
timestamp 1667941163
transform 1 0 22632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0481_
timestamp 1667941163
transform 1 0 10212 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0482_
timestamp 1667941163
transform 1 0 19964 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0483_
timestamp 1667941163
transform 1 0 19412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0484_
timestamp 1667941163
transform 1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0485_
timestamp 1667941163
transform 1 0 3956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0486_
timestamp 1667941163
transform 1 0 1840 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0487_
timestamp 1667941163
transform 1 0 12420 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0488_
timestamp 1667941163
transform 1 0 3220 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0489_
timestamp 1667941163
transform 1 0 3220 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1667941163
transform 1 0 2116 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0492_
timestamp 1667941163
transform 1 0 17296 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0493_
timestamp 1667941163
transform 1 0 2300 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0494_
timestamp 1667941163
transform 1 0 8372 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0495_
timestamp 1667941163
transform 1 0 18124 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1667941163
transform 1 0 9108 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1667941163
transform 1 0 9568 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0498_
timestamp 1667941163
transform 1 0 3128 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0499_
timestamp 1667941163
transform 1 0 8372 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0500_
timestamp 1667941163
transform 1 0 18768 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0501_
timestamp 1667941163
transform 1 0 20976 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502_
timestamp 1667941163
transform 1 0 2484 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1667941163
transform 1 0 7912 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0504_
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0505_
timestamp 1667941163
transform 1 0 4416 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0506_
timestamp 1667941163
transform 1 0 2484 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0507_
timestamp 1667941163
transform 1 0 1840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0508_
timestamp 1667941163
transform 1 0 13524 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0509_
timestamp 1667941163
transform 1 0 20424 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0510_
timestamp 1667941163
transform 1 0 18308 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0511_
timestamp 1667941163
transform 1 0 20608 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0512_
timestamp 1667941163
transform 1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0513_
timestamp 1667941163
transform 1 0 23092 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1667941163
transform 1 0 20516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0515_
timestamp 1667941163
transform 1 0 23184 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0516_
timestamp 1667941163
transform 1 0 20976 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0517_
timestamp 1667941163
transform 1 0 20884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0518_
timestamp 1667941163
transform 1 0 19228 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0519_
timestamp 1667941163
transform 1 0 21988 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp 1667941163
transform 1 0 20148 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0521_
timestamp 1667941163
transform 1 0 22080 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0522_
timestamp 1667941163
transform 1 0 19136 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0523_
timestamp 1667941163
transform 1 0 19412 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0524_
timestamp 1667941163
transform 1 0 23368 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0525_
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0526_
timestamp 1667941163
transform 1 0 10304 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0527_
timestamp 1667941163
transform 1 0 5796 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0528_
timestamp 1667941163
transform 1 0 14536 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1667941163
transform 1 0 16836 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0530_
timestamp 1667941163
transform 1 0 21160 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0531_
timestamp 1667941163
transform 1 0 4232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1667941163
transform 1 0 10488 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1667941163
transform 1 0 6532 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0534_
timestamp 1667941163
transform 1 0 18308 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0535_
timestamp 1667941163
transform 1 0 11040 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0536_
timestamp 1667941163
transform 1 0 19320 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0537_
timestamp 1667941163
transform 1 0 23920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1667941163
transform 1 0 20700 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0539_
timestamp 1667941163
transform 1 0 22908 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0540_
timestamp 1667941163
transform 1 0 19780 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0541_
timestamp 1667941163
transform 1 0 23828 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0542_
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0543_
timestamp 1667941163
transform 1 0 19872 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0544_
timestamp 1667941163
transform 1 0 21988 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0545_
timestamp 1667941163
transform 1 0 22632 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0546_
timestamp 1667941163
transform 1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1667941163
transform 1 0 19688 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0548_
timestamp 1667941163
transform 1 0 23276 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0549_
timestamp 1667941163
transform 1 0 11040 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1667941163
transform 1 0 15456 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0551_
timestamp 1667941163
transform 1 0 18676 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0552_
timestamp 1667941163
transform 1 0 21436 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0553_
timestamp 1667941163
transform 1 0 11776 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0554_
timestamp 1667941163
transform 1 0 6716 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0555_
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1667941163
transform 1 0 10488 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0557_
timestamp 1667941163
transform 1 0 14628 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0558_
timestamp 1667941163
transform 1 0 19964 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0559_
timestamp 1667941163
transform 1 0 20608 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0560_
timestamp 1667941163
transform 1 0 14444 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0561_
timestamp 1667941163
transform 1 0 16100 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0562_
timestamp 1667941163
transform 1 0 8372 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0563_
timestamp 1667941163
transform 1 0 11776 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0564_
timestamp 1667941163
transform 1 0 17204 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1667941163
transform 1 0 21988 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0566_
timestamp 1667941163
transform 1 0 18032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0567_
timestamp 1667941163
transform 1 0 19780 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0568_
timestamp 1667941163
transform 1 0 24564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0569_
timestamp 1667941163
transform 1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0570_
timestamp 1667941163
transform 1 0 13156 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1667941163
transform 1 0 16928 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0572_
timestamp 1667941163
transform 1 0 22448 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0573_
timestamp 1667941163
transform 1 0 21252 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0574_
timestamp 1667941163
transform 1 0 6440 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0575_
timestamp 1667941163
transform 1 0 24564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0576_
timestamp 1667941163
transform 1 0 25208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 1667941163
transform 1 0 20976 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0578_
timestamp 1667941163
transform 1 0 20792 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0579_
timestamp 1667941163
transform 1 0 19964 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0580_
timestamp 1667941163
transform 1 0 20240 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0581_
timestamp 1667941163
transform 1 0 16100 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0582_
timestamp 1667941163
transform 1 0 21988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1667941163
transform 1 0 23368 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0584_
timestamp 1667941163
transform 1 0 21988 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0585_
timestamp 1667941163
transform 1 0 7268 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0586_
timestamp 1667941163
transform 1 0 17480 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0587_
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1667941163
transform 1 0 5704 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0589_
timestamp 1667941163
transform 1 0 6532 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0590_
timestamp 1667941163
transform 1 0 22724 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1667941163
transform 1 0 13156 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0592_
timestamp 1667941163
transform 1 0 15456 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0593_
timestamp 1667941163
transform 1 0 20148 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0594_
timestamp 1667941163
transform 1 0 17848 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0595_
timestamp 1667941163
transform 1 0 14536 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1667941163
transform 1 0 6900 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0597_
timestamp 1667941163
transform 1 0 9108 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0598_
timestamp 1667941163
transform 1 0 3220 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0599_
timestamp 1667941163
transform 1 0 13248 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0600_
timestamp 1667941163
transform 1 0 3772 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1667941163
transform 1 0 20056 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0602_
timestamp 1667941163
transform 1 0 3128 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0603_
timestamp 1667941163
transform 1 0 4600 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0604_
timestamp 1667941163
transform 1 0 20424 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0605_
timestamp 1667941163
transform 1 0 10948 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0606_
timestamp 1667941163
transform 1 0 6532 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1667941163
transform 1 0 5152 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0608_
timestamp 1667941163
transform 1 0 8280 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 1667941163
transform 1 0 2576 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1667941163
transform 1 0 24564 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0611_
timestamp 1667941163
transform 1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0612_
timestamp 1667941163
transform 1 0 4324 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0613_
timestamp 1667941163
transform 1 0 23460 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 1667941163
transform 1 0 31280 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0615_
timestamp 1667941163
transform 1 0 31464 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0617_
timestamp 1667941163
transform 1 0 12788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0618_
timestamp 1667941163
transform 1 0 31004 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1667941163
transform 1 0 9568 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 1667941163
transform 1 0 19412 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 1667941163
transform 1 0 20700 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1667941163
transform 1 0 27140 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 1667941163
transform 1 0 7728 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0624_
timestamp 1667941163
transform 1 0 12880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1667941163
transform 1 0 29256 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 1667941163
transform 1 0 2484 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 1667941163
transform 1 0 36708 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1667941163
transform 1 0 10948 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 1667941163
transform 1 0 4048 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0630_
timestamp 1667941163
transform 1 0 29716 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1667941163
transform 1 0 25392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1667941163
transform 1 0 20792 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1667941163
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 1667941163
transform 1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0635_
timestamp 1667941163
transform 1 0 27968 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0636_
timestamp 1667941163
transform 1 0 5796 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1667941163
transform 1 0 29716 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1667941163
transform 1 0 6532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0639_
timestamp 1667941163
transform 1 0 3128 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1667941163
transform 1 0 3956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1667941163
transform 1 0 25668 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0642_
timestamp 1667941163
transform 1 0 22724 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1667941163
transform 1 0 25208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0644_
timestamp 1667941163
transform 1 0 37444 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1667941163
transform 1 0 21436 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1667941163
transform 1 0 23736 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1667941163
transform 1 0 26036 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0648_
timestamp 1667941163
transform 1 0 21620 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0649_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1564 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1667941163
transform 1 0 17480 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0651_
timestamp 1667941163
transform 1 0 10856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1667941163
transform 1 0 9660 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0653_
timestamp 1667941163
transform 1 0 5704 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0654_
timestamp 1667941163
transform 1 0 28704 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1667941163
transform 1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1667941163
transform 1 0 16560 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1667941163
transform 1 0 21344 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 1667941163
transform 1 0 1840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1667941163
transform 1 0 17020 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0660_
timestamp 1667941163
transform 1 0 22080 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0661_
timestamp 1667941163
transform 1 0 1840 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0662_
timestamp 1667941163
transform 1 0 5244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0663_
timestamp 1667941163
transform 1 0 22080 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1667941163
transform 1 0 19412 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1667941163
transform 1 0 23092 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0666_
timestamp 1667941163
transform 1 0 23552 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1667941163
transform 1 0 6164 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1667941163
transform 1 0 8096 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 1667941163
transform 1 0 14352 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 1667941163
transform 1 0 27232 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0671_
timestamp 1667941163
transform 1 0 11040 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1667941163
transform 1 0 29716 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1667941163
transform 1 0 19412 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1667941163
transform 1 0 21252 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1667941163
transform 1 0 15364 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1667941163
transform 1 0 10948 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0678_
timestamp 1667941163
transform 1 0 4232 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1667941163
transform 1 0 4232 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0680_
timestamp 1667941163
transform 1 0 27324 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1667941163
transform 1 0 7728 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1667941163
transform 1 0 7084 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1667941163
transform 1 0 18216 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1667941163
transform 1 0 26036 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1667941163
transform 1 0 4784 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1667941163
transform 1 0 23644 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1667941163
transform 1 0 22080 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1667941163
transform 1 0 7360 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1667941163
transform 1 0 6440 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1667941163
transform 1 0 20240 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1667941163
transform 1 0 21988 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1667941163
transform 1 0 27876 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1667941163
transform 1 0 28244 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1667941163
transform 1 0 18492 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1667941163
transform 1 0 24932 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1667941163
transform 1 0 14076 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1667941163
transform 1 0 1932 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1667941163
transform 1 0 9108 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1667941163
transform 1 0 29900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1667941163
transform 1 0 29532 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1667941163
transform 1 0 3956 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0703_
timestamp 1667941163
transform 1 0 19412 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform 1 0 30544 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1667941163
transform 1 0 27968 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1667941163
transform 1 0 5152 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0707_
timestamp 1667941163
transform 1 0 1840 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1667941163
transform 1 0 21252 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0710_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16836 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _0711_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16836 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1667941163
transform 1 0 1932 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1667941163
transform 1 0 1840 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1667941163
transform 1 0 1840 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1667941163
transform 1 0 6532 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1667941163
transform 1 0 5244 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1667941163
transform 1 0 1932 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1667941163
transform 1 0 3128 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1667941163
transform 1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1667941163
transform 1 0 6716 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0722_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17204 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1667941163
transform 1 0 4416 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1667941163
transform 1 0 5888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1667941163
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1667941163
transform 1 0 11960 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1667941163
transform 1 0 6532 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1667941163
transform 1 0 3220 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1667941163
transform 1 0 21068 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1667941163
transform 1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1667941163
transform 1 0 23184 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1667941163
transform 1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0733_
timestamp 1667941163
transform 1 0 18952 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1667941163
transform 1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1667941163
transform 1 0 12144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1667941163
transform 1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1667941163
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1667941163
transform 1 0 22080 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1667941163
transform 1 0 23828 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1667941163
transform 1 0 11684 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1667941163
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1667941163
transform 1 0 16928 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0744_
timestamp 1667941163
transform 1 0 18400 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1667941163
transform 1 0 17664 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1667941163
transform 1 0 12328 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1667941163
transform 1 0 6532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1667941163
transform 1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform 1 0 3864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1667941163
transform 1 0 6072 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1667941163
transform 1 0 17940 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1667941163
transform 1 0 17480 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1667941163
transform 1 0 10948 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1667941163
transform 1 0 5336 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0755_
timestamp 1667941163
transform 1 0 19412 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1667941163
transform 1 0 9292 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1667941163
transform 1 0 9568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1667941163
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1667941163
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1667941163
transform 1 0 25208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1667941163
transform 1 0 23276 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1667941163
transform 1 0 20516 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1667941163
transform 1 0 23920 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1667941163
transform 1 0 23276 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0766_
timestamp 1667941163
transform 1 0 18032 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1667941163
transform 1 0 11960 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1667941163
transform 1 0 9108 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1667941163
transform 1 0 9752 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1667941163
transform 1 0 14352 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1667941163
transform 1 0 22632 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1667941163
transform 1 0 21804 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1667941163
transform 1 0 24564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1667941163
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1667941163
transform 1 0 27140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1667941163
transform 1 0 4600 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0777_
timestamp 1667941163
transform 1 0 18124 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1667941163
transform 1 0 6992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1667941163
transform 1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1667941163
transform 1 0 25208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1667941163
transform 1 0 26496 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1667941163
transform 1 0 18032 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1667941163
transform 1 0 23552 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1667941163
transform 1 0 7636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1667941163
transform 1 0 6072 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1667941163
transform 1 0 3956 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0788_
timestamp 1667941163
transform 1 0 18768 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1667941163
transform 1 0 7820 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1667941163
transform 1 0 5152 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1667941163
transform 1 0 4416 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1667941163
transform 1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1667941163
transform 1 0 4784 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1667941163
transform 1 0 4600 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1667941163
transform 1 0 11316 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1667941163
transform 1 0 11684 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1667941163
transform 1 0 11684 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1667941163
transform 1 0 8740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0799_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16836 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1667941163
transform 1 0 3956 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1667941163
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1667941163
transform 1 0 3220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1667941163
transform 1 0 4600 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1667941163
transform 1 0 4140 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0806_
timestamp 1667941163
transform 1 0 4784 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1667941163
transform 1 0 3956 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 23184 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1667941163
transform 1 0 5428 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0810_
timestamp 1667941163
transform 1 0 16744 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1667941163
transform 1 0 3956 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1667941163
transform 1 0 13156 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1667941163
transform 1 0 15640 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1667941163
transform 1 0 4600 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1667941163
transform 1 0 5244 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1667941163
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1667941163
transform 1 0 16836 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1667941163
transform 1 0 3312 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1667941163
transform 1 0 5060 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1667941163
transform 1 0 16744 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0821_
timestamp 1667941163
transform 1 0 17940 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1667941163
transform 1 0 10948 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1667941163
transform 1 0 9292 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1667941163
transform 1 0 12512 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1667941163
transform 1 0 6532 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1667941163
transform 1 0 12328 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1667941163
transform 1 0 16100 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1667941163
transform 1 0 14260 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1667941163
transform 1 0 8372 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1667941163
transform 1 0 23184 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0832_
timestamp 1667941163
transform 1 0 18032 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1667941163
transform 1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1667941163
transform 1 0 18584 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1667941163
transform 1 0 19412 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1667941163
transform 1 0 22540 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1667941163
transform 1 0 23368 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1667941163
transform 1 0 10212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1667941163
transform 1 0 24564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1667941163
transform 1 0 24564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1667941163
transform 1 0 8280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1667941163
transform 1 0 23920 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _0843_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1564 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0844_
timestamp 1667941163
transform 1 0 1932 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0845_
timestamp 1667941163
transform 1 0 4140 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0846_
timestamp 1667941163
transform 1 0 4232 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0847_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9016 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0848_
timestamp 1667941163
transform 1 0 6532 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0849_
timestamp 1667941163
transform 1 0 1564 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0850_
timestamp 1667941163
transform 1 0 4048 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0851_
timestamp 1667941163
transform 1 0 6624 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0852_
timestamp 1667941163
transform 1 0 6440 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0853_
timestamp 1667941163
transform 1 0 4232 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0854_
timestamp 1667941163
transform 1 0 4324 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0855_
timestamp 1667941163
transform 1 0 9476 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0856_
timestamp 1667941163
transform 1 0 5520 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0857_
timestamp 1667941163
transform 1 0 6348 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0858_
timestamp 1667941163
transform 1 0 7820 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0859_
timestamp 1667941163
transform 1 0 14260 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0860_
timestamp 1667941163
transform 1 0 11960 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0861_
timestamp 1667941163
transform 1 0 14260 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0862_
timestamp 1667941163
transform 1 0 13984 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0863_
timestamp 1667941163
transform 1 0 11684 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0864_
timestamp 1667941163
transform 1 0 9384 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0865_
timestamp 1667941163
transform 1 0 13800 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0866_
timestamp 1667941163
transform 1 0 9936 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0867_
timestamp 1667941163
transform 1 0 11960 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0868_
timestamp 1667941163
transform 1 0 8280 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0869_
timestamp 1667941163
transform 1 0 8832 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0870_
timestamp 1667941163
transform 1 0 6716 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0871_
timestamp 1667941163
transform 1 0 11960 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0872_
timestamp 1667941163
transform 1 0 14260 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0873_
timestamp 1667941163
transform 1 0 11776 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0874_
timestamp 1667941163
transform 1 0 11960 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0875_
timestamp 1667941163
transform 1 0 1564 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0876_
timestamp 1667941163
transform 1 0 2852 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0877_
timestamp 1667941163
transform 1 0 6808 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0878_
timestamp 1667941163
transform 1 0 9108 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0879_
timestamp 1667941163
transform 1 0 10580 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0880_
timestamp 1667941163
transform 1 0 10672 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0881_
timestamp 1667941163
transform 1 0 14260 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0882_
timestamp 1667941163
transform 1 0 6716 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0883_
timestamp 1667941163
transform 1 0 8924 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0884_
timestamp 1667941163
transform 1 0 9660 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0885_
timestamp 1667941163
transform 1 0 11500 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0886_
timestamp 1667941163
transform 1 0 9292 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0887_
timestamp 1667941163
transform 1 0 14260 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0888_
timestamp 1667941163
transform 1 0 11684 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0889_
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0890_
timestamp 1667941163
transform 1 0 9016 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0891_
timestamp 1667941163
transform 1 0 6532 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0892_
timestamp 1667941163
transform 1 0 3956 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0893_
timestamp 1667941163
transform 1 0 5244 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0894_
timestamp 1667941163
transform 1 0 7176 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0895_
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0896_
timestamp 1667941163
transform 1 0 13524 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0897_
timestamp 1667941163
transform 1 0 9752 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0898_
timestamp 1667941163
transform 1 0 9016 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0899_
timestamp 1667941163
transform 1 0 13432 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0900_
timestamp 1667941163
transform 1 0 14260 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0901_
timestamp 1667941163
transform 1 0 14260 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0902_
timestamp 1667941163
transform 1 0 9384 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0903_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13248 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0904_
timestamp 1667941163
transform 1 0 13156 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0905_
timestamp 1667941163
transform 1 0 14260 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0906_
timestamp 1667941163
transform 1 0 16836 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0907_
timestamp 1667941163
transform 1 0 13892 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0908_
timestamp 1667941163
transform 1 0 14260 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0909_
timestamp 1667941163
transform 1 0 14260 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0910_
timestamp 1667941163
transform 1 0 13432 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0911_
timestamp 1667941163
transform 1 0 3772 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0912_
timestamp 1667941163
transform 1 0 6716 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0913_
timestamp 1667941163
transform 1 0 2024 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0914_
timestamp 1667941163
transform 1 0 1564 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0915_
timestamp 1667941163
transform 1 0 2024 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0916_
timestamp 1667941163
transform 1 0 2760 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0917_
timestamp 1667941163
transform 1 0 1564 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0918_
timestamp 1667941163
transform 1 0 4232 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0919_
timestamp 1667941163
transform 1 0 1564 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0920_
timestamp 1667941163
transform 1 0 9752 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0921_
timestamp 1667941163
transform 1 0 14260 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0922_
timestamp 1667941163
transform 1 0 9384 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0923_
timestamp 1667941163
transform 1 0 1656 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0924_
timestamp 1667941163
transform 1 0 2208 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0925_
timestamp 1667941163
transform 1 0 3864 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0926_
timestamp 1667941163
transform 1 0 4600 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0927_
timestamp 1667941163
transform 1 0 3956 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0928_
timestamp 1667941163
transform 1 0 1564 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0929_
timestamp 1667941163
transform 1 0 1656 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0930_
timestamp 1667941163
transform 1 0 1564 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0931_
timestamp 1667941163
transform 1 0 11960 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0932_
timestamp 1667941163
transform 1 0 3312 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0933_
timestamp 1667941163
transform 1 0 6808 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0934_
timestamp 1667941163
transform 1 0 14260 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0935_
timestamp 1667941163
transform 1 0 12144 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0936_
timestamp 1667941163
transform 1 0 8740 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0937_
timestamp 1667941163
transform 1 0 9108 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0938_
timestamp 1667941163
transform 1 0 6808 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0939_
timestamp 1667941163
transform 1 0 11960 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0940_
timestamp 1667941163
transform 1 0 1564 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0941_
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0942_
timestamp 1667941163
transform 1 0 13248 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0943_
timestamp 1667941163
transform 1 0 1564 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0944_
timestamp 1667941163
transform 1 0 8832 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0945_
timestamp 1667941163
transform 1 0 9568 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0946_
timestamp 1667941163
transform 1 0 10856 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0947_
timestamp 1667941163
transform 1 0 9476 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0948_
timestamp 1667941163
transform 1 0 12972 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0949_
timestamp 1667941163
transform 1 0 14260 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0950_
timestamp 1667941163
transform 1 0 11684 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0951_
timestamp 1667941163
transform 1 0 3956 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0952_
timestamp 1667941163
transform 1 0 4232 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0953_
timestamp 1667941163
transform 1 0 3772 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0954_
timestamp 1667941163
transform 1 0 7176 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0955_
timestamp 1667941163
transform 1 0 6532 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0956_
timestamp 1667941163
transform 1 0 12972 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0957_
timestamp 1667941163
transform 1 0 1564 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0958_
timestamp 1667941163
transform 1 0 6808 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0959_
timestamp 1667941163
transform 1 0 7176 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0960_
timestamp 1667941163
transform 1 0 6072 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0961_
timestamp 1667941163
transform 1 0 5244 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0962_
timestamp 1667941163
transform 1 0 11224 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_1  _0988_
timestamp 1667941163
transform 1 0 29900 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0989_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21068 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0990_
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0991_
timestamp 1667941163
transform 1 0 23092 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0992_
timestamp 1667941163
transform 1 0 8096 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0993_
timestamp 1667941163
transform 1 0 3128 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1667941163
transform 1 0 24564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0995_
timestamp 1667941163
transform 1 0 16468 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0996_
timestamp 1667941163
transform 1 0 37812 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0997_
timestamp 1667941163
transform 1 0 16836 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1667941163
transform 1 0 37720 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0999_
timestamp 1667941163
transform 1 0 22080 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1667941163
transform 1 0 28520 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1001_
timestamp 1667941163
transform 1 0 24472 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1002_
timestamp 1667941163
transform 1 0 19688 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 1667941163
transform 1 0 27140 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1667941163
transform 1 0 16100 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1005_
timestamp 1667941163
transform 1 0 35144 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1667941163
transform 1 0 14812 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1007_
timestamp 1667941163
transform 1 0 22816 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1008_
timestamp 1667941163
transform 1 0 32660 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1667941163
transform 1 0 16100 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1011_
timestamp 1667941163
transform 1 0 8924 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1667941163
transform 1 0 9108 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1667941163
transform 1 0 23828 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1667941163
transform 1 0 4508 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1015_
timestamp 1667941163
transform 1 0 17572 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1667941163
transform 1 0 37812 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1667941163
transform 1 0 32292 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1667941163
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1019_
timestamp 1667941163
transform 1 0 17664 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1020_
timestamp 1667941163
transform 1 0 14904 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1021_
timestamp 1667941163
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1667941163
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1023_
timestamp 1667941163
transform 1 0 37352 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 1667941163
transform 1 0 25944 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1667941163
transform 1 0 9016 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1667941163
transform 1 0 33212 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1027_
timestamp 1667941163
transform 1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1028_
timestamp 1667941163
transform 1 0 37444 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1667941163
transform 1 0 37812 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1030_
timestamp 1667941163
transform 1 0 30452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1667941163
transform 1 0 34132 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1032_
timestamp 1667941163
transform 1 0 5888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1667941163
transform 1 0 30176 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1667941163
transform 1 0 37720 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1035_
timestamp 1667941163
transform 1 0 5152 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1036_
timestamp 1667941163
transform 1 0 21988 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1037_
timestamp 1667941163
transform 1 0 10580 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1038_
timestamp 1667941163
transform 1 0 4324 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1667941163
transform 1 0 21988 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1040_
timestamp 1667941163
transform 1 0 3312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1667941163
transform 1 0 1748 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1042_
timestamp 1667941163
transform 1 0 2300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1043_
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1044_
timestamp 1667941163
transform 1 0 37352 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1045_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5244 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1046_
timestamp 1667941163
transform 1 0 5244 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1047__142 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6992 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1047_
timestamp 1667941163
transform 1 0 6900 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1048_
timestamp 1667941163
transform 1 0 14444 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1049_
timestamp 1667941163
transform 1 0 19412 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1050_
timestamp 1667941163
transform 1 0 6808 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1051_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1564 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1052_
timestamp 1667941163
transform 1 0 16560 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1053_
timestamp 1667941163
transform 1 0 2668 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1054_
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1055_
timestamp 1667941163
transform 1 0 6624 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1056_
timestamp 1667941163
transform 1 0 17020 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1057_
timestamp 1667941163
transform 1 0 15088 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1058_
timestamp 1667941163
transform 1 0 21988 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1059_
timestamp 1667941163
transform 1 0 19228 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1059__143
timestamp 1667941163
transform 1 0 20608 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1060_
timestamp 1667941163
transform 1 0 9384 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1061_
timestamp 1667941163
transform 1 0 21988 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1062_
timestamp 1667941163
transform 1 0 18492 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1063_
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1064_
timestamp 1667941163
transform 1 0 3864 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1065_
timestamp 1667941163
transform 1 0 6624 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1066_
timestamp 1667941163
transform 1 0 7176 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1067_
timestamp 1667941163
transform 1 0 19412 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1068_
timestamp 1667941163
transform 1 0 15272 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1069_
timestamp 1667941163
transform 1 0 19412 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1070_
timestamp 1667941163
transform 1 0 21988 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1071__144
timestamp 1667941163
transform 1 0 20608 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1071_
timestamp 1667941163
transform 1 0 20332 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1072_
timestamp 1667941163
transform 1 0 19412 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1073_
timestamp 1667941163
transform 1 0 15548 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1074_
timestamp 1667941163
transform 1 0 19596 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1075_
timestamp 1667941163
transform 1 0 21988 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1076_
timestamp 1667941163
transform 1 0 16468 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1077_
timestamp 1667941163
transform 1 0 21620 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1078_
timestamp 1667941163
transform 1 0 17940 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1079_
timestamp 1667941163
transform 1 0 16836 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1080_
timestamp 1667941163
transform 1 0 9752 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1081_
timestamp 1667941163
transform 1 0 16468 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1082_
timestamp 1667941163
transform 1 0 21988 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1083__145
timestamp 1667941163
transform 1 0 22264 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1083_
timestamp 1667941163
transform 1 0 17572 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1084_
timestamp 1667941163
transform 1 0 20516 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1085_
timestamp 1667941163
transform 1 0 13340 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1086_
timestamp 1667941163
transform 1 0 13800 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1087_
timestamp 1667941163
transform 1 0 19412 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1088_
timestamp 1667941163
transform 1 0 17388 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1089_
timestamp 1667941163
transform 1 0 12420 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1090_
timestamp 1667941163
transform 1 0 16836 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1091_
timestamp 1667941163
transform 1 0 14260 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1092_
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1093_
timestamp 1667941163
transform 1 0 11592 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1094_
timestamp 1667941163
transform 1 0 1656 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1095__146
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1095_
timestamp 1667941163
transform 1 0 7360 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1096_
timestamp 1667941163
transform 1 0 14536 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1097_
timestamp 1667941163
transform 1 0 18032 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1098_
timestamp 1667941163
transform 1 0 20516 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1099_
timestamp 1667941163
transform 1 0 12236 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1100_
timestamp 1667941163
transform 1 0 21988 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1101_
timestamp 1667941163
transform 1 0 17756 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1102_
timestamp 1667941163
transform 1 0 10580 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1103_
timestamp 1667941163
transform 1 0 13248 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1104_
timestamp 1667941163
transform 1 0 14996 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1105_
timestamp 1667941163
transform 1 0 16468 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1106_
timestamp 1667941163
transform 1 0 18676 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1107__147
timestamp 1667941163
transform 1 0 21988 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1107_
timestamp 1667941163
transform 1 0 20056 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1108_
timestamp 1667941163
transform 1 0 18124 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1109_
timestamp 1667941163
transform 1 0 17572 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1110_
timestamp 1667941163
transform 1 0 16468 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1111_
timestamp 1667941163
transform 1 0 18768 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1112_
timestamp 1667941163
transform 1 0 18216 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1113_
timestamp 1667941163
transform 1 0 16468 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1114_
timestamp 1667941163
transform 1 0 17204 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1115_
timestamp 1667941163
transform 1 0 19412 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1116_
timestamp 1667941163
transform 1 0 20884 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1117_
timestamp 1667941163
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1118_
timestamp 1667941163
transform 1 0 20240 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1119__148
timestamp 1667941163
transform 1 0 5520 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1119_
timestamp 1667941163
transform 1 0 15548 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1120_
timestamp 1667941163
transform 1 0 17756 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1121_
timestamp 1667941163
transform 1 0 10028 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1122_
timestamp 1667941163
transform 1 0 18768 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1123_
timestamp 1667941163
transform 1 0 15272 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1124_
timestamp 1667941163
transform 1 0 14260 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1125_
timestamp 1667941163
transform 1 0 8556 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1126_
timestamp 1667941163
transform 1 0 16468 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1127_
timestamp 1667941163
transform 1 0 9200 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1128_
timestamp 1667941163
transform 1 0 11408 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1129_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22264 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1129__149
timestamp 1667941163
transform 1 0 22632 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1130_
timestamp 1667941163
transform 1 0 21988 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1131_
timestamp 1667941163
transform 1 0 22448 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1132_
timestamp 1667941163
transform 1 0 18124 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1133_
timestamp 1667941163
transform 1 0 17664 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1134_
timestamp 1667941163
transform 1 0 15640 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1135_
timestamp 1667941163
transform 1 0 18032 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1136_
timestamp 1667941163
transform 1 0 17664 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1137_
timestamp 1667941163
transform 1 0 19872 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1138_
timestamp 1667941163
transform 1 0 20884 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1139_
timestamp 1667941163
transform 1 0 19136 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1140_
timestamp 1667941163
transform 1 0 16836 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1141_
timestamp 1667941163
transform 1 0 24840 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1141__150
timestamp 1667941163
transform 1 0 25024 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1142_
timestamp 1667941163
transform 1 0 15548 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1143_
timestamp 1667941163
transform 1 0 19780 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1144_
timestamp 1667941163
transform 1 0 21620 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1145_
timestamp 1667941163
transform 1 0 18952 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1146_
timestamp 1667941163
transform 1 0 6532 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1147__151
timestamp 1667941163
transform 1 0 3956 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1147_
timestamp 1667941163
transform 1 0 2116 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1148_
timestamp 1667941163
transform 1 0 2576 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1149_
timestamp 1667941163
transform 1 0 11684 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1150_
timestamp 1667941163
transform 1 0 4416 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1151_
timestamp 1667941163
transform 1 0 12880 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1152_
timestamp 1667941163
transform 1 0 20700 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1153_
timestamp 1667941163
transform 1 0 9752 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1154__152
timestamp 1667941163
transform 1 0 2944 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1154_
timestamp 1667941163
transform 1 0 2760 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1155_
timestamp 1667941163
transform 1 0 16836 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1156_
timestamp 1667941163
transform 1 0 8004 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1157_
timestamp 1667941163
transform 1 0 19412 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1158_
timestamp 1667941163
transform 1 0 9292 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1159_
timestamp 1667941163
transform 1 0 16836 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1160_
timestamp 1667941163
transform 1 0 1656 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1161_
timestamp 1667941163
transform 1 0 1564 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1162__153
timestamp 1667941163
transform 1 0 3128 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1162_
timestamp 1667941163
transform 1 0 2300 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1163_
timestamp 1667941163
transform 1 0 3956 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1164_
timestamp 1667941163
transform 1 0 3128 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1165_
timestamp 1667941163
transform 1 0 14904 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1166_
timestamp 1667941163
transform 1 0 1656 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1167_
timestamp 1667941163
transform 1 0 11776 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1168__154
timestamp 1667941163
transform 1 0 6164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1168_
timestamp 1667941163
transform 1 0 16836 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1169_
timestamp 1667941163
transform 1 0 16560 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1170_
timestamp 1667941163
transform 1 0 18400 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1171_
timestamp 1667941163
transform 1 0 16836 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1172__155
timestamp 1667941163
transform 1 0 20976 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1172_
timestamp 1667941163
transform 1 0 20792 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1173_
timestamp 1667941163
transform 1 0 16100 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1174_
timestamp 1667941163
transform 1 0 21988 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1175_
timestamp 1667941163
transform 1 0 20700 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1176__156
timestamp 1667941163
transform 1 0 8096 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1176_
timestamp 1667941163
transform 1 0 8004 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1177_
timestamp 1667941163
transform 1 0 16284 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1178_
timestamp 1667941163
transform 1 0 7636 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1179_
timestamp 1667941163
transform 1 0 12144 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1180__157
timestamp 1667941163
transform 1 0 12236 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1180_
timestamp 1667941163
transform 1 0 12880 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1181_
timestamp 1667941163
transform 1 0 17664 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1182_
timestamp 1667941163
transform 1 0 12696 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1183_
timestamp 1667941163
transform 1 0 19412 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1184__158
timestamp 1667941163
transform 1 0 16836 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1184_
timestamp 1667941163
transform 1 0 16192 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1185_
timestamp 1667941163
transform 1 0 13432 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1186_
timestamp 1667941163
transform 1 0 14996 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1187_
timestamp 1667941163
transform 1 0 14260 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1188__159
timestamp 1667941163
transform 1 0 24748 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1188_
timestamp 1667941163
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1189_
timestamp 1667941163
transform 1 0 7820 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1190_
timestamp 1667941163
transform 1 0 23276 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1191_
timestamp 1667941163
transform 1 0 10396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1192__160
timestamp 1667941163
transform 1 0 17756 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1192_
timestamp 1667941163
transform 1 0 17664 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1193_
timestamp 1667941163
transform 1 0 9292 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1194_
timestamp 1667941163
transform 1 0 16836 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1195_
timestamp 1667941163
transform 1 0 10396 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1196_
timestamp 1667941163
transform 1 0 8188 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1197__161
timestamp 1667941163
transform 1 0 14260 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1197_
timestamp 1667941163
transform 1 0 14260 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1198_
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1199_
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1200_
timestamp 1667941163
transform 1 0 15364 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1201_
timestamp 1667941163
transform 1 0 5428 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1202_
timestamp 1667941163
transform 1 0 26036 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1203__162
timestamp 1667941163
transform 1 0 25668 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1203_
timestamp 1667941163
transform 1 0 25944 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1204_
timestamp 1667941163
transform 1 0 22172 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1205_
timestamp 1667941163
transform 1 0 24840 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1206_
timestamp 1667941163
transform 1 0 24840 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1207_
timestamp 1667941163
transform 1 0 24012 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1208_
timestamp 1667941163
transform 1 0 12512 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1209_
timestamp 1667941163
transform 1 0 16836 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1209__163
timestamp 1667941163
transform 1 0 16928 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1210_
timestamp 1667941163
transform 1 0 10396 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1211_
timestamp 1667941163
transform 1 0 11960 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1212_
timestamp 1667941163
transform 1 0 18768 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1213_
timestamp 1667941163
transform 1 0 16928 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1214_
timestamp 1667941163
transform 1 0 27140 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1215__164
timestamp 1667941163
transform 1 0 25944 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1215_
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1216_
timestamp 1667941163
transform 1 0 22448 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1217_
timestamp 1667941163
transform 1 0 24564 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1218_
timestamp 1667941163
transform 1 0 27140 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1219_
timestamp 1667941163
transform 1 0 23276 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1220_
timestamp 1667941163
transform 1 0 12604 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1221_
timestamp 1667941163
transform 1 0 3956 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1222_
timestamp 1667941163
transform 1 0 5152 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1223__165
timestamp 1667941163
transform 1 0 2484 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1223_
timestamp 1667941163
transform 1 0 2300 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1224_
timestamp 1667941163
transform 1 0 20700 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1225_
timestamp 1667941163
transform 1 0 14260 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1226_
timestamp 1667941163
transform 1 0 23644 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1227_
timestamp 1667941163
transform 1 0 11684 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1228_
timestamp 1667941163
transform 1 0 11776 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1229_
timestamp 1667941163
transform 1 0 3220 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1230_
timestamp 1667941163
transform 1 0 20976 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1231_
timestamp 1667941163
transform 1 0 24564 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1232_
timestamp 1667941163
transform 1 0 17664 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1233_
timestamp 1667941163
transform 1 0 18124 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1234_
timestamp 1667941163
transform 1 0 20056 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1235__166
timestamp 1667941163
transform 1 0 22448 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1235_
timestamp 1667941163
transform 1 0 19412 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1236_
timestamp 1667941163
transform 1 0 6532 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1237_
timestamp 1667941163
transform 1 0 17204 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1238_
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1239_
timestamp 1667941163
transform 1 0 18032 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1240_
timestamp 1667941163
transform 1 0 16468 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1241_
timestamp 1667941163
transform 1 0 15640 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1242_
timestamp 1667941163
transform 1 0 6716 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1243_
timestamp 1667941163
transform 1 0 19504 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8924 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk
timestamp 1667941163
transform 1 0 5060 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1667941163
transform 1 0 6900 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1667941163
transform 1 0 3956 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1667941163
transform 1 0 7636 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1667941163
transform 1 0 11684 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1667941163
transform 1 0 12052 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1667941163
transform 1 0 11684 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1667941163
transform 1 0 16560 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1667941163
transform 1 0 3956 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1667941163
transform 1 0 6900 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1667941163
transform 1 0 3956 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1667941163
transform 1 0 5060 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1667941163
transform 1 0 9844 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1667941163
transform 1 0 15824 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1667941163
transform 1 0 9108 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1667941163
transform 1 0 12144 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 1564 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 5796 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 3956 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 23368 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1667941163
transform 1 0 3220 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37444 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1667941163
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1667941163
transform 1 0 25300 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1667941163
transform 1 0 37996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1667941163
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1667941163
transform 1 0 37996 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1667941163
transform 1 0 1564 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1667941163
transform 1 0 1564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1667941163
transform 1 0 12420 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1667941163
transform 1 0 37444 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1667941163
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1667941163
transform 1 0 4692 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1667941163
transform 1 0 36156 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1667941163
transform 1 0 37444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1667941163
transform 1 0 1564 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1667941163
transform 1 0 21160 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1667941163
transform 1 0 37444 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1667941163
transform 1 0 37996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1667941163
transform 1 0 1564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1667941163
transform 1 0 38088 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1667941163
transform 1 0 1564 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1667941163
transform 1 0 1564 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1667941163
transform 1 0 37996 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1667941163
transform 1 0 36708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1667941163
transform 1 0 18584 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1667941163
transform 1 0 31004 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1667941163
transform 1 0 37996 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1667941163
transform 1 0 23276 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1667941163
transform 1 0 2668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1667941163
transform 1 0 1564 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1667941163
transform 1 0 1564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1667941163
transform 1 0 32292 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1667941163
transform 1 0 37444 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1667941163
transform 1 0 5336 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp 1667941163
transform 1 0 37444 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1667941163
transform 1 0 36708 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1667941163
transform 1 0 2944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1667941163
transform 1 0 38088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1667941163
transform 1 0 38088 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1667941163
transform 1 0 3864 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1667941163
transform 1 0 2668 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1667941163
transform 1 0 37444 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1667941163
transform 1 0 5796 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1667941163
transform 1 0 2944 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1667941163
transform 1 0 38088 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1667941163
transform 1 0 7636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1667941163
transform 1 0 2576 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1667941163
transform 1 0 25208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1667941163
transform 1 0 38088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1667941163
transform 1 0 13524 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1667941163
transform 1 0 30452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1667941163
transform 1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1667941163
transform 1 0 1564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1667941163
transform 1 0 38088 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1667941163
transform 1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1667941163
transform 1 0 4600 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1667941163
transform 1 0 5060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1667941163
transform 1 0 21988 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1667941163
transform 1 0 35512 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1667941163
transform 1 0 38088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1667941163
transform 1 0 2300 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1667941163
transform 1 0 2576 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1667941163
transform 1 0 3220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1667941163
transform 1 0 2576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1667941163
transform 1 0 38088 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1667941163
transform 1 0 22632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1667941163
transform 1 0 28612 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1667941163
transform 1 0 1564 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1667941163
transform 1 0 6532 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1667941163
transform 1 0 27784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1667941163
transform 1 0 7176 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1667941163
transform 1 0 1564 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1667941163
transform 1 0 38088 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform 1 0 1564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 15548 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform 1 0 37996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 33028 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform 1 0 3956 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform 1 0 10856 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1667941163
transform 1 0 1564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1667941163
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1667941163
transform 1 0 13432 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1667941163
transform 1 0 33580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1667941163
transform 1 0 7820 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1667941163
transform 1 0 37996 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1667941163
transform 1 0 16836 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1667941163
transform 1 0 11684 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1667941163
transform 1 0 1564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1667941163
transform 1 0 1564 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1667941163
transform 1 0 18216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1667941163
transform 1 0 1564 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1667941163
transform 1 0 34868 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1667941163
transform 1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1667941163
transform 1 0 37996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1667941163
transform 1 0 37996 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1667941163
transform 1 0 27876 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1667941163
transform 1 0 37260 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1667941163
transform 1 0 17480 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1667941163
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1667941163
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1667941163
transform 1 0 14260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1667941163
transform 1 0 9108 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1667941163
transform 1 0 37996 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1667941163
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1667941163
transform 1 0 1564 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1667941163
transform 1 0 1564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1667941163
transform 1 0 37996 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1667941163
transform 1 0 37996 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1667941163
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1667941163
transform 1 0 1564 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1667941163
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1667941163
transform 1 0 6532 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1667941163
transform 1 0 3036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1667941163
transform 1 0 25944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1667941163
transform 1 0 9752 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1667941163
transform 1 0 1564 0 -1 30464
box -38 -48 406 592
<< labels >>
flabel metal3 s 200 28568 800 28688 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 0 nsew signal input
flabel metal2 s 5814 39200 5870 39800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 1 nsew signal input
flabel metal2 s 12898 200 12954 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 2 nsew signal input
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 3 nsew signal input
flabel metal3 s 200 26528 800 26648 0 FreeSans 480 0 0 0 ccff_head
port 4 nsew signal input
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 ccff_tail
port 5 nsew signal tristate
flabel metal3 s 39200 30608 39800 30728 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal2 s 25134 39200 25190 39800 0 FreeSans 224 90 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 39200 8168 39800 8288 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal3 s 200 688 800 808 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal3 s 39200 35368 39800 35488 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 200 19048 800 19168 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal2 s 26422 39200 26478 39800 0 FreeSans 224 90 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 200 23128 800 23248 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal2 s 12254 39200 12310 39800 0 FreeSans 224 90 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal3 s 39200 10888 39800 11008 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 16 nsew signal input
flabel metal2 s 28354 200 28410 800 0 FreeSans 224 90 0 0 chanx_left_in[2]
port 17 nsew signal input
flabel metal2 s 4526 39200 4582 39800 0 FreeSans 224 90 0 0 chanx_left_in[3]
port 18 nsew signal input
flabel metal2 s 36082 39200 36138 39800 0 FreeSans 224 90 0 0 chanx_left_in[4]
port 19 nsew signal input
flabel metal2 s 37370 39200 37426 39800 0 FreeSans 224 90 0 0 chanx_left_in[5]
port 20 nsew signal input
flabel metal3 s 200 5448 800 5568 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 21 nsew signal input
flabel metal2 s 20626 200 20682 800 0 FreeSans 224 90 0 0 chanx_left_in[7]
port 22 nsew signal input
flabel metal3 s 39200 27888 39800 28008 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 23 nsew signal input
flabel metal3 s 39200 12248 39800 12368 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 24 nsew signal input
flabel metal2 s 15474 39200 15530 39800 0 FreeSans 224 90 0 0 chanx_left_out[0]
port 25 nsew signal tristate
flabel metal2 s 39302 200 39358 800 0 FreeSans 224 90 0 0 chanx_left_out[10]
port 26 nsew signal tristate
flabel metal2 s 32862 39200 32918 39800 0 FreeSans 224 90 0 0 chanx_left_out[11]
port 27 nsew signal tristate
flabel metal2 s 17406 200 17462 800 0 FreeSans 224 90 0 0 chanx_left_out[12]
port 28 nsew signal tristate
flabel metal2 s 3238 39200 3294 39800 0 FreeSans 224 90 0 0 chanx_left_out[13]
port 29 nsew signal tristate
flabel metal2 s 10966 200 11022 800 0 FreeSans 224 90 0 0 chanx_left_out[14]
port 30 nsew signal tristate
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 31 nsew signal tristate
flabel metal2 s 25134 200 25190 800 0 FreeSans 224 90 0 0 chanx_left_out[16]
port 32 nsew signal tristate
flabel metal3 s 39200 12928 39800 13048 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 33 nsew signal tristate
flabel metal3 s 39200 27208 39800 27328 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 34 nsew signal tristate
flabel metal2 s 34794 200 34850 800 0 FreeSans 224 90 0 0 chanx_left_out[1]
port 35 nsew signal tristate
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chanx_left_out[2]
port 36 nsew signal tristate
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 chanx_left_out[3]
port 37 nsew signal tristate
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chanx_left_out[4]
port 38 nsew signal tristate
flabel metal2 s 33506 200 33562 800 0 FreeSans 224 90 0 0 chanx_left_out[5]
port 39 nsew signal tristate
flabel metal3 s 39200 16328 39800 16448 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 40 nsew signal tristate
flabel metal2 s 7746 39200 7802 39800 0 FreeSans 224 90 0 0 chanx_left_out[7]
port 41 nsew signal tristate
flabel metal3 s 39200 23808 39800 23928 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 42 nsew signal tristate
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 chanx_left_out[9]
port 43 nsew signal tristate
flabel metal3 s 39200 32648 39800 32768 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 44 nsew signal input
flabel metal3 s 200 4088 800 4208 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 45 nsew signal input
flabel metal3 s 39200 17688 39800 17808 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 46 nsew signal input
flabel metal3 s 200 31288 800 31408 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 47 nsew signal input
flabel metal3 s 200 35368 800 35488 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 48 nsew signal input
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 49 nsew signal input
flabel metal3 s 39200 1368 39800 1488 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 50 nsew signal input
flabel metal2 s 21270 39200 21326 39800 0 FreeSans 224 90 0 0 chanx_right_in[16]
port 51 nsew signal input
flabel metal2 s 18694 39200 18750 39800 0 FreeSans 224 90 0 0 chanx_right_in[17]
port 52 nsew signal input
flabel metal2 s 30930 39200 30986 39800 0 FreeSans 224 90 0 0 chanx_right_in[18]
port 53 nsew signal input
flabel metal3 s 39200 37408 39800 37528 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 54 nsew signal input
flabel metal2 s 23202 39200 23258 39800 0 FreeSans 224 90 0 0 chanx_right_in[2]
port 55 nsew signal input
flabel metal2 s 9678 200 9734 800 0 FreeSans 224 90 0 0 chanx_right_in[3]
port 56 nsew signal input
flabel metal3 s 200 17008 800 17128 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 57 nsew signal input
flabel metal3 s 200 7488 800 7608 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 58 nsew signal input
flabel metal2 s 31574 200 31630 800 0 FreeSans 224 90 0 0 chanx_right_in[6]
port 59 nsew signal input
flabel metal3 s 39200 688 39800 808 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 60 nsew signal input
flabel metal3 s 200 14968 800 15088 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 61 nsew signal input
flabel metal3 s 39200 7488 39800 7608 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 62 nsew signal input
flabel metal2 s 10966 39200 11022 39800 0 FreeSans 224 90 0 0 chanx_right_out[0]
port 63 nsew signal tristate
flabel metal3 s 200 38768 800 38888 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 64 nsew signal tristate
flabel metal3 s 200 21768 800 21888 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 65 nsew signal tristate
flabel metal2 s 16118 200 16174 800 0 FreeSans 224 90 0 0 chanx_right_out[12]
port 66 nsew signal tristate
flabel metal3 s 200 25168 800 25288 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 67 nsew signal tristate
flabel metal2 s 34150 39200 34206 39800 0 FreeSans 224 90 0 0 chanx_right_out[14]
port 68 nsew signal tristate
flabel metal2 s 22558 200 22614 800 0 FreeSans 224 90 0 0 chanx_right_out[15]
port 69 nsew signal tristate
flabel metal2 s 29642 200 29698 800 0 FreeSans 224 90 0 0 chanx_right_out[16]
port 70 nsew signal tristate
flabel metal3 s 39200 24488 39800 24608 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 71 nsew signal tristate
flabel metal3 s 39200 4768 39800 4888 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 72 nsew signal tristate
flabel metal2 s 27710 39200 27766 39800 0 FreeSans 224 90 0 0 chanx_right_out[1]
port 73 nsew signal tristate
flabel metal3 s 39200 38768 39800 38888 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 74 nsew signal tristate
flabel metal2 s 17406 39200 17462 39800 0 FreeSans 224 90 0 0 chanx_right_out[3]
port 75 nsew signal tristate
flabel metal2 s 662 200 718 800 0 FreeSans 224 90 0 0 chanx_right_out[4]
port 76 nsew signal tristate
flabel metal2 s 5170 200 5226 800 0 FreeSans 224 90 0 0 chanx_right_out[5]
port 77 nsew signal tristate
flabel metal2 s 13542 39200 13598 39800 0 FreeSans 224 90 0 0 chanx_right_out[6]
port 78 nsew signal tristate
flabel metal2 s 9034 39200 9090 39800 0 FreeSans 224 90 0 0 chanx_right_out[7]
port 79 nsew signal tristate
flabel metal3 s 39200 21088 39800 21208 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 80 nsew signal tristate
flabel metal3 s 39200 14288 39800 14408 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 81 nsew signal tristate
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 82 nsew signal input
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 83 nsew signal input
flabel metal3 s 39200 2728 39800 2848 0 FreeSans 480 0 0 0 chany_bottom_in[11]
port 84 nsew signal input
flabel metal3 s 39200 15648 39800 15768 0 FreeSans 480 0 0 0 chany_bottom_in[12]
port 85 nsew signal input
flabel metal3 s 200 27208 800 27328 0 FreeSans 480 0 0 0 chany_bottom_in[13]
port 86 nsew signal input
flabel metal2 s 2594 39200 2650 39800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 87 nsew signal input
flabel metal2 s 36726 200 36782 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 88 nsew signal input
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 chany_bottom_in[16]
port 89 nsew signal input
flabel metal2 s 18 39200 74 39800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 90 nsew signal input
flabel metal2 s 38658 39200 38714 39800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 91 nsew signal input
flabel metal2 s 8390 200 8446 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 92 nsew signal input
flabel metal3 s 200 18368 800 18488 0 FreeSans 480 0 0 0 chany_bottom_in[2]
port 93 nsew signal input
flabel metal2 s 23846 200 23902 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 94 nsew signal input
flabel metal2 s 38014 200 38070 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 95 nsew signal input
flabel metal2 s 14186 39200 14242 39800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 96 nsew signal input
flabel metal2 s 30286 200 30342 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 97 nsew signal input
flabel metal2 s 3882 200 3938 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 98 nsew signal input
flabel metal3 s 200 13608 800 13728 0 FreeSans 480 0 0 0 chany_bottom_in[8]
port 99 nsew signal input
flabel metal3 s 39200 4088 39800 4208 0 FreeSans 480 0 0 0 chany_bottom_in[9]
port 100 nsew signal input
flabel metal3 s 39200 29248 39800 29368 0 FreeSans 480 0 0 0 chany_bottom_out[0]
port 101 nsew signal tristate
flabel metal3 s 39200 20408 39800 20528 0 FreeSans 480 0 0 0 chany_bottom_out[10]
port 102 nsew signal tristate
flabel metal2 s 32862 200 32918 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 103 nsew signal tristate
flabel metal3 s 200 23808 800 23928 0 FreeSans 480 0 0 0 chany_bottom_out[12]
port 104 nsew signal tristate
flabel metal3 s 39200 9528 39800 9648 0 FreeSans 480 0 0 0 chany_bottom_out[13]
port 105 nsew signal tristate
flabel metal3 s 200 31968 800 32088 0 FreeSans 480 0 0 0 chany_bottom_out[14]
port 106 nsew signal tristate
flabel metal3 s 39200 22448 39800 22568 0 FreeSans 480 0 0 0 chany_bottom_out[15]
port 107 nsew signal tristate
flabel metal3 s 39200 34008 39800 34128 0 FreeSans 480 0 0 0 chany_bottom_out[16]
port 108 nsew signal tristate
flabel metal2 s 36082 200 36138 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 109 nsew signal tristate
flabel metal3 s 39200 36048 39800 36168 0 FreeSans 480 0 0 0 chany_bottom_out[18]
port 110 nsew signal tristate
flabel metal3 s 200 33328 800 33448 0 FreeSans 480 0 0 0 chany_bottom_out[1]
port 111 nsew signal tristate
flabel metal3 s 200 2048 800 2168 0 FreeSans 480 0 0 0 chany_bottom_out[2]
port 112 nsew signal tristate
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 chany_bottom_out[3]
port 113 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 114 nsew signal tristate
flabel metal2 s 25778 200 25834 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 115 nsew signal tristate
flabel metal3 s 200 38088 800 38208 0 FreeSans 480 0 0 0 chany_bottom_out[6]
port 116 nsew signal tristate
flabel metal2 s 9678 39200 9734 39800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 117 nsew signal tristate
flabel metal2 s 24490 39200 24546 39800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 118 nsew signal tristate
flabel metal3 s 200 29928 800 30048 0 FreeSans 480 0 0 0 chany_bottom_out[9]
port 119 nsew signal tristate
flabel metal2 s 6458 200 6514 800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 120 nsew signal input
flabel metal2 s 1950 200 2006 800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 121 nsew signal input
flabel metal3 s 200 8848 800 8968 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 122 nsew signal input
flabel metal2 s 21914 39200 21970 39800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 123 nsew signal input
flabel metal2 s 18050 200 18106 800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 124 nsew signal input
flabel metal2 s 35438 39200 35494 39800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 125 nsew signal input
flabel metal3 s 39200 6128 39800 6248 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
port 126 nsew signal input
flabel metal3 s 200 36728 800 36848 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
port 127 nsew signal input
flabel metal3 s 200 11568 800 11688 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
port 128 nsew signal input
flabel metal2 s 7102 200 7158 800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
port 129 nsew signal input
flabel metal2 s 14186 200 14242 800 0 FreeSans 224 90 0 0 pReset
port 130 nsew signal input
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 prog_clk
port 131 nsew signal input
flabel metal3 s 39200 25848 39800 25968 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 132 nsew signal input
flabel metal2 s 21914 200 21970 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 133 nsew signal input
flabel metal2 s 29642 39200 29698 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 134 nsew signal input
flabel metal2 s 28354 39200 28410 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 135 nsew signal input
flabel metal2 s 1306 39200 1362 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 136 nsew signal input
flabel metal2 s 6458 39200 6514 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 137 nsew signal input
flabel metal2 s 27066 200 27122 800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
port 138 nsew signal input
flabel metal3 s 200 10208 800 10328 0 FreeSans 480 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
port 139 nsew signal input
flabel metal3 s 200 34688 800 34808 0 FreeSans 480 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
port 140 nsew signal input
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
port 141 nsew signal input
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 142 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 142 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 143 nsew ground bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal2 15594 3264 15594 3264 0 _0000_
rlabel metal2 21206 6273 21206 6273 0 _0001_
rlabel metal2 15318 5372 15318 5372 0 _0002_
rlabel metal1 19550 4624 19550 4624 0 _0003_
rlabel metal2 8694 6001 8694 6001 0 _0004_
rlabel metal3 16284 1700 16284 1700 0 _0005_
rlabel via2 12098 3995 12098 3995 0 _0006_
rlabel metal2 9246 11560 9246 11560 0 _0007_
rlabel metal1 9936 15334 9936 15334 0 _0008_
rlabel metal2 14490 17374 14490 17374 0 _0009_
rlabel metal1 11737 11050 11737 11050 0 _0010_
rlabel metal1 21344 4454 21344 4454 0 _0011_
rlabel metal2 17618 4913 17618 4913 0 _0012_
rlabel metal2 12558 1768 12558 1768 0 _0013_
rlabel metal1 16107 3434 16107 3434 0 _0014_
rlabel metal1 5382 2822 5382 2822 0 _0015_
rlabel metal2 14030 3570 14030 3570 0 _0016_
rlabel metal2 24058 3111 24058 3111 0 _0017_
rlabel metal1 16291 2346 16291 2346 0 _0018_
rlabel metal2 18262 3876 18262 3876 0 _0019_
rlabel metal1 17940 3094 17940 3094 0 _0020_
rlabel metal1 16107 7786 16107 7786 0 _0021_
rlabel metal1 15686 6807 15686 6807 0 _0022_
rlabel metal2 13846 5525 13846 5525 0 _0023_
rlabel metal2 6210 14790 6210 14790 0 _0024_
rlabel via2 4094 16405 4094 16405 0 _0025_
rlabel metal1 7774 12342 7774 12342 0 _0026_
rlabel metal2 2668 19210 2668 19210 0 _0027_
rlabel metal1 4692 8466 4692 8466 0 _0028_
rlabel metal2 4186 7548 4186 7548 0 _0029_
rlabel metal3 6187 18156 6187 18156 0 _0030_
rlabel metal1 5474 24786 5474 24786 0 _0031_
rlabel metal2 11454 16184 11454 16184 0 _0032_
rlabel metal1 11553 12138 11553 12138 0 _0033_
rlabel metal1 15686 11159 15686 11159 0 _0034_
rlabel metal1 9200 8330 9200 8330 0 _0035_
rlabel metal1 4048 4794 4048 4794 0 _0036_
rlabel metal1 3496 5338 3496 5338 0 _0037_
rlabel metal1 4041 12886 4041 12886 0 _0038_
rlabel metal1 5198 24106 5198 24106 0 _0039_
rlabel metal1 2576 24038 2576 24038 0 _0040_
rlabel metal1 3457 16490 3457 16490 0 _0041_
rlabel metal1 4055 4522 4055 4522 0 _0042_
rlabel metal1 4002 6834 4002 6834 0 _0043_
rlabel metal1 22540 4998 22540 4998 0 _0044_
rlabel metal1 5106 4454 5106 4454 0 _0045_
rlabel metal2 8280 19380 8280 19380 0 _0046_
rlabel metal1 14306 9146 14306 9146 0 _0047_
rlabel metal1 14674 18054 14674 18054 0 _0048_
rlabel metal2 9522 19822 9522 19822 0 _0049_
rlabel metal2 9844 18666 9844 18666 0 _0050_
rlabel via3 7659 17884 7659 17884 0 _0051_
rlabel metal2 16974 16796 16974 16796 0 _0052_
rlabel via3 3197 12308 3197 12308 0 _0053_
rlabel metal1 7905 12886 7905 12886 0 _0054_
rlabel metal1 16836 19686 16836 19686 0 _0055_
rlabel metal3 7107 13260 7107 13260 0 _0056_
rlabel metal2 11086 18292 11086 18292 0 _0057_
rlabel metal1 9890 8806 9890 8806 0 _0058_
rlabel metal2 12650 9554 12650 9554 0 _0059_
rlabel metal1 6578 19414 6578 19414 0 _0060_
rlabel metal1 12466 11764 12466 11764 0 _0061_
rlabel metal2 16238 15164 16238 15164 0 _0062_
rlabel metal1 13393 13226 13393 13226 0 _0063_
rlabel metal1 8556 9622 8556 9622 0 _0064_
rlabel via2 6854 11781 6854 11781 0 _0065_
rlabel metal2 20286 10863 20286 10863 0 _0066_
rlabel metal2 18722 13532 18722 13532 0 _0067_
rlabel metal2 19504 9996 19504 9996 0 _0068_
rlabel metal2 14398 10438 14398 10438 0 _0069_
rlabel metal3 13248 1836 13248 1836 0 _0070_
rlabel metal1 9752 2618 9752 2618 0 _0071_
rlabel via2 9614 4165 9614 4165 0 _0072_
rlabel metal1 7781 4522 7781 4522 0 _0073_
rlabel metal1 8464 2822 8464 2822 0 _0074_
rlabel via2 21574 4029 21574 4029 0 _0075_
rlabel via3 2139 19244 2139 19244 0 _0076_
rlabel metal2 1978 27013 1978 27013 0 _0077_
rlabel metal1 1748 26826 1748 26826 0 _0078_
rlabel metal1 1564 26758 1564 26758 0 _0079_
rlabel metal1 7222 9146 7222 9146 0 _0080_
rlabel metal2 7774 19652 7774 19652 0 _0081_
rlabel metal1 2484 10166 2484 10166 0 _0082_
rlabel metal2 690 19686 690 19686 0 _0083_
rlabel metal1 6663 7446 6663 7446 0 _0084_
rlabel metal1 7038 8058 7038 8058 0 _0085_
rlabel metal1 4784 6426 4784 6426 0 _0086_
rlabel metal2 6026 9554 6026 9554 0 _0087_
rlabel metal1 12926 15368 12926 15368 0 _0088_
rlabel metal1 11868 14246 11868 14246 0 _0089_
rlabel metal1 6854 11866 6854 11866 0 _0090_
rlabel metal1 7721 18326 7721 18326 0 _0091_
rlabel metal1 19688 11798 19688 11798 0 _0092_
rlabel metal1 13524 6834 13524 6834 0 _0093_
rlabel metal1 15831 8874 15831 8874 0 _0094_
rlabel metal1 11316 6970 11316 6970 0 _0095_
rlabel metal1 12436 8534 12436 8534 0 _0096_
rlabel metal1 11500 3094 11500 3094 0 _0097_
rlabel metal1 21804 6834 21804 6834 0 _0098_
rlabel metal1 17158 2618 17158 2618 0 _0099_
rlabel metal1 22080 3366 22080 3366 0 _0100_
rlabel metal1 18492 2618 18492 2618 0 _0101_
rlabel metal2 21482 7021 21482 7021 0 _0102_
rlabel metal1 10672 11526 10672 11526 0 _0103_
rlabel metal2 13662 14110 13662 14110 0 _0104_
rlabel metal1 16974 13974 16974 13974 0 _0105_
rlabel metal1 17572 17102 17572 17102 0 _0106_
rlabel metal1 12512 10778 12512 10778 0 _0107_
rlabel metal1 5796 8398 5796 8398 0 _0108_
rlabel metal1 4561 13974 4561 13974 0 _0109_
rlabel metal2 7498 19788 7498 19788 0 _0110_
rlabel metal1 7268 18598 7268 18598 0 _0111_
rlabel metal2 12650 16626 12650 16626 0 _0112_
rlabel metal1 12243 16490 12243 16490 0 _0113_
rlabel metal2 15042 15096 15042 15096 0 _0114_
rlabel metal1 6486 9078 6486 9078 0 _0115_
rlabel metal2 9706 3230 9706 3230 0 _0116_
rlabel metal1 10396 2550 10396 2550 0 _0117_
rlabel metal2 9430 3043 9430 3043 0 _0118_
rlabel metal2 24702 2074 24702 2074 0 _0119_
rlabel metal1 6256 20774 6256 20774 0 _0120_
rlabel metal2 7774 2482 7774 2482 0 _0121_
rlabel metal2 21206 10948 21206 10948 0 _0122_
rlabel metal2 18078 3179 18078 3179 0 _0123_
rlabel metal1 4462 8432 4462 8432 0 _0124_
rlabel metal3 4140 12716 4140 12716 0 _0125_
rlabel metal1 16698 19822 16698 19822 0 _0126_
rlabel metal2 14306 18564 14306 18564 0 _0127_
rlabel metal1 18124 8534 18124 8534 0 _0128_
rlabel metal1 25024 23086 25024 23086 0 _0129_
rlabel metal2 28290 17476 28290 17476 0 _0130_
rlabel metal2 27830 20876 27830 20876 0 _0131_
rlabel metal2 11914 29308 11914 29308 0 _0132_
rlabel metal2 13202 26996 13202 26996 0 _0133_
rlabel metal2 17710 29308 17710 29308 0 _0134_
rlabel metal2 22218 21148 22218 21148 0 _0135_
rlabel metal1 27968 12818 27968 12818 0 _0136_
rlabel metal2 28014 15164 28014 15164 0 _0137_
rlabel metal2 10718 25670 10718 25670 0 _0138_
rlabel metal1 9338 24752 9338 24752 0 _0139_
rlabel metal1 16192 24582 16192 24582 0 _0140_
rlabel metal2 10074 26044 10074 26044 0 _0141_
rlabel metal1 18998 27642 18998 27642 0 _0142_
rlabel metal2 15870 21318 15870 21318 0 _0143_
rlabel metal1 25852 19346 25852 19346 0 _0144_
rlabel metal2 13754 21114 13754 21114 0 _0145_
rlabel metal1 16790 26384 16790 26384 0 _0146_
rlabel metal2 22126 14586 22126 14586 0 _0147_
rlabel metal1 15502 25908 15502 25908 0 _0148_
rlabel metal2 13938 23800 13938 23800 0 _0149_
rlabel metal1 8970 28016 8970 28016 0 _0150_
rlabel metal2 19366 15844 19366 15844 0 _0151_
rlabel metal1 24288 7378 24288 7378 0 _0152_
rlabel metal2 19642 14586 19642 14586 0 _0153_
rlabel metal1 4922 2482 4922 2482 0 _0154_
rlabel metal2 20102 7888 20102 7888 0 _0155_
rlabel metal1 1288 10030 1288 10030 0 _0156_
rlabel metal1 21114 11696 21114 11696 0 _0157_
rlabel metal1 16882 2346 16882 2346 0 _0158_
rlabel metal1 5336 20502 5336 20502 0 _0159_
rlabel metal1 5382 26350 5382 26350 0 _0160_
rlabel metal2 6670 23970 6670 23970 0 _0161_
rlabel metal1 12880 21590 12880 21590 0 _0162_
rlabel metal1 20286 18394 20286 18394 0 _0163_
rlabel metal1 5888 19482 5888 19482 0 _0164_
rlabel metal1 1794 20536 1794 20536 0 _0165_
rlabel metal1 19642 15538 19642 15538 0 _0166_
rlabel metal1 3036 19414 3036 19414 0 _0167_
rlabel metal2 4002 20332 4002 20332 0 _0168_
rlabel metal1 7406 21862 7406 21862 0 _0169_
rlabel metal1 17250 23800 17250 23800 0 _0170_
rlabel metal1 15456 15130 15456 15130 0 _0171_
rlabel metal2 13294 10744 13294 10744 0 _0172_
rlabel metal2 22862 8670 22862 8670 0 _0173_
rlabel metal2 9614 24752 9614 24752 0 _0174_
rlabel metal2 14674 22406 14674 22406 0 _0175_
rlabel metal1 18354 22678 18354 22678 0 _0176_
rlabel metal1 5106 21896 5106 21896 0 _0177_
rlabel metal2 5842 15079 5842 15079 0 _0178_
rlabel metal1 6904 19754 6904 19754 0 _0179_
rlabel metal2 7406 16728 7406 16728 0 _0180_
rlabel metal1 19684 16490 19684 16490 0 _0181_
rlabel metal1 16054 23766 16054 23766 0 _0182_
rlabel metal2 20378 8194 20378 8194 0 _0183_
rlabel metal2 22310 17136 22310 17136 0 _0184_
rlabel metal2 20930 13464 20930 13464 0 _0185_
rlabel metal2 21022 13464 21022 13464 0 _0186_
rlabel metal2 19918 13447 19918 13447 0 _0187_
rlabel metal1 20746 12920 20746 12920 0 _0188_
rlabel metal1 21390 15674 21390 15674 0 _0189_
rlabel via2 16698 7803 16698 7803 0 _0190_
rlabel metal1 22586 7820 22586 7820 0 _0191_
rlabel metal1 18170 10744 18170 10744 0 _0192_
rlabel metal2 16238 6324 16238 6324 0 _0193_
rlabel metal2 9246 20230 9246 20230 0 _0194_
rlabel metal1 17526 8942 17526 8942 0 _0195_
rlabel metal1 20240 9622 20240 9622 0 _0196_
rlabel metal1 17986 3706 17986 3706 0 _0197_
rlabel metal1 21666 12138 21666 12138 0 _0198_
rlabel metal2 13570 18377 13570 18377 0 _0199_
rlabel metal1 13800 19414 13800 19414 0 _0200_
rlabel metal1 20378 20434 20378 20434 0 _0201_
rlabel metal1 17480 21114 17480 21114 0 _0202_
rlabel metal1 12650 22984 12650 22984 0 _0203_
rlabel metal1 16652 15062 16652 15062 0 _0204_
rlabel metal2 14490 14008 14490 14008 0 _0205_
rlabel metal1 10212 20842 10212 20842 0 _0206_
rlabel metal2 11822 21461 11822 21461 0 _0207_
rlabel metal2 1886 21250 1886 21250 0 _0208_
rlabel metal1 7590 22712 7590 22712 0 _0209_
rlabel metal2 14766 14654 14766 14654 0 _0210_
rlabel metal1 18354 12886 18354 12886 0 _0211_
rlabel metal1 20470 25466 20470 25466 0 _0212_
rlabel metal2 12466 21794 12466 21794 0 _0213_
rlabel metal2 21574 20264 21574 20264 0 _0214_
rlabel metal2 17986 24990 17986 24990 0 _0215_
rlabel metal1 10994 21930 10994 21930 0 _0216_
rlabel metal1 14122 24854 14122 24854 0 _0217_
rlabel metal1 15410 22950 15410 22950 0 _0218_
rlabel metal2 21114 3740 21114 3740 0 _0219_
rlabel metal1 19458 3094 19458 3094 0 _0220_
rlabel metal1 20378 5882 20378 5882 0 _0221_
rlabel metal1 18446 7752 18446 7752 0 _0222_
rlabel metal1 18814 13974 18814 13974 0 _0223_
rlabel metal1 18584 3706 18584 3706 0 _0224_
rlabel metal2 23414 7582 23414 7582 0 _0225_
rlabel metal1 19182 19414 19182 19414 0 _0226_
rlabel metal1 19826 5678 19826 5678 0 _0227_
rlabel metal2 20746 7922 20746 7922 0 _0228_
rlabel metal2 20930 6562 20930 6562 0 _0229_
rlabel metal1 20976 16218 20976 16218 0 _0230_
rlabel metal2 13294 6664 13294 6664 0 _0231_
rlabel metal2 20470 2145 20470 2145 0 _0232_
rlabel metal1 15778 3128 15778 3128 0 _0233_
rlabel metal1 18722 16150 18722 16150 0 _0234_
rlabel metal1 10672 22678 10672 22678 0 _0235_
rlabel metal1 18722 23290 18722 23290 0 _0236_
rlabel metal1 16238 18394 16238 18394 0 _0237_
rlabel metal2 14490 23256 14490 23256 0 _0238_
rlabel viali 8782 21590 8782 21590 0 _0239_
rlabel metal1 14904 12750 14904 12750 0 _0240_
rlabel metal1 7544 16218 7544 16218 0 _0241_
rlabel metal1 11040 16218 11040 16218 0 _0242_
rlabel metal1 23000 10098 23000 10098 0 _0243_
rlabel metal2 22218 4488 22218 4488 0 _0244_
rlabel metal1 20194 3910 20194 3910 0 _0245_
rlabel metal1 18354 15368 18354 15368 0 _0246_
rlabel metal1 18032 14314 18032 14314 0 _0247_
rlabel metal1 15870 6358 15870 6358 0 _0248_
rlabel metal1 19366 5610 19366 5610 0 _0249_
rlabel metal2 19090 9996 19090 9996 0 _0250_
rlabel metal1 20148 4250 20148 4250 0 _0251_
rlabel metal1 21114 8840 21114 8840 0 _0252_
rlabel metal1 20240 6222 20240 6222 0 _0253_
rlabel metal2 17066 5032 17066 5032 0 _0254_
rlabel metal1 17802 6086 17802 6086 0 _0255_
rlabel metal1 15916 11798 15916 11798 0 _0256_
rlabel metal1 19228 17306 19228 17306 0 _0257_
rlabel metal3 19642 13668 19642 13668 0 _0258_
rlabel metal1 20516 11866 20516 11866 0 _0259_
rlabel metal1 1886 10778 1886 10778 0 _0260_
rlabel metal2 2254 25126 2254 25126 0 _0261_
rlabel via3 4715 20740 4715 20740 0 _0262_
rlabel metal1 10396 15878 10396 15878 0 _0263_
rlabel metal2 2576 19108 2576 19108 0 _0264_
rlabel metal1 13064 20298 13064 20298 0 _0265_
rlabel metal1 21022 20570 21022 20570 0 _0266_
rlabel metal2 9982 21726 9982 21726 0 _0267_
rlabel metal2 2990 23358 2990 23358 0 _0268_
rlabel metal2 9706 10591 9706 10591 0 _0269_
rlabel metal1 8740 20026 8740 20026 0 _0270_
rlabel metal1 19136 20434 19136 20434 0 _0271_
rlabel metal2 9522 22005 9522 22005 0 _0272_
rlabel metal2 17066 19550 17066 19550 0 _0273_
rlabel metal2 1886 24072 1886 24072 0 _0274_
rlabel metal2 2530 25772 2530 25772 0 _0275_
rlabel metal1 2576 20842 2576 20842 0 _0276_
rlabel metal1 4232 20842 4232 20842 0 _0277_
rlabel metal2 3358 23086 3358 23086 0 _0278_
rlabel metal1 15180 17578 15180 17578 0 _0279_
rlabel metal1 1932 21590 1932 21590 0 _0280_
rlabel metal2 12558 20910 12558 20910 0 _0281_
rlabel metal1 14398 2550 14398 2550 0 _0282_
rlabel metal1 18124 14450 18124 14450 0 _0283_
rlabel metal2 22770 3723 22770 3723 0 _0284_
rlabel metal1 12926 10608 12926 10608 0 _0285_
rlabel metal1 21022 7242 21022 7242 0 _0286_
rlabel metal1 17526 16762 17526 16762 0 _0287_
rlabel metal2 22218 8364 22218 8364 0 _0288_
rlabel metal2 20930 10846 20930 10846 0 _0289_
rlabel metal2 8234 26316 8234 26316 0 _0290_
rlabel metal1 16514 24072 16514 24072 0 _0291_
rlabel metal2 7866 26860 7866 26860 0 _0292_
rlabel metal1 12098 22678 12098 22678 0 _0293_
rlabel metal1 14214 25194 14214 25194 0 _0294_
rlabel metal1 19918 14586 19918 14586 0 _0295_
rlabel metal1 13524 24106 13524 24106 0 _0296_
rlabel metal1 21068 14246 21068 14246 0 _0297_
rlabel metal1 16514 25194 16514 25194 0 _0298_
rlabel metal1 13616 20434 13616 20434 0 _0299_
rlabel metal2 15226 24990 15226 24990 0 _0300_
rlabel metal1 14168 20978 14168 20978 0 _0301_
rlabel metal1 24840 18666 24840 18666 0 _0302_
rlabel metal2 14030 20944 14030 20944 0 _0303_
rlabel metal2 23506 18904 23506 18904 0 _0304_
rlabel metal2 10074 18513 10074 18513 0 _0305_
rlabel metal2 17894 26894 17894 26894 0 _0306_
rlabel metal2 9522 24140 9522 24140 0 _0307_
rlabel metal2 17066 27438 17066 27438 0 _0308_
rlabel metal1 11684 27982 11684 27982 0 _0309_
rlabel metal1 8786 23698 8786 23698 0 _0310_
rlabel metal2 14490 24616 14490 24616 0 _0311_
rlabel metal1 9890 25772 9890 25772 0 _0312_
rlabel metal2 6210 25500 6210 25500 0 _0313_
rlabel metal2 15594 19550 15594 19550 0 _0314_
rlabel metal1 6164 23154 6164 23154 0 _0315_
rlabel metal2 27554 13124 27554 13124 0 _0316_
rlabel metal2 26174 14620 26174 14620 0 _0317_
rlabel metal2 22402 20740 22402 20740 0 _0318_
rlabel metal1 26036 12274 26036 12274 0 _0319_
rlabel metal1 25070 14348 25070 14348 0 _0320_
rlabel metal1 24840 21454 24840 21454 0 _0321_
rlabel metal2 12742 27166 12742 27166 0 _0322_
rlabel metal1 17296 28594 17296 28594 0 _0323_
rlabel metal2 10626 28254 10626 28254 0 _0324_
rlabel metal2 12190 26520 12190 26520 0 _0325_
rlabel metal1 18584 26894 18584 26894 0 _0326_
rlabel metal1 17342 27506 17342 27506 0 _0327_
rlabel metal2 27370 17340 27370 17340 0 _0328_
rlabel metal2 26818 20060 26818 20060 0 _0329_
rlabel metal1 23644 22950 23644 22950 0 _0330_
rlabel metal1 26726 16218 26726 16218 0 _0331_
rlabel metal2 27370 18428 27370 18428 0 _0332_
rlabel metal1 24058 23630 24058 23630 0 _0333_
rlabel metal1 13248 16490 13248 16490 0 _0334_
rlabel metal1 4554 19754 4554 19754 0 _0335_
rlabel metal1 9108 12410 9108 12410 0 _0336_
rlabel metal2 2530 22712 2530 22712 0 _0337_
rlabel metal1 22218 9622 22218 9622 0 _0338_
rlabel metal1 14490 19720 14490 19720 0 _0339_
rlabel metal1 24426 18326 24426 18326 0 _0340_
rlabel metal2 13846 20077 13846 20077 0 _0341_
rlabel metal2 13018 17000 13018 17000 0 _0342_
rlabel metal1 4416 22066 4416 22066 0 _0343_
rlabel metal2 21758 10268 21758 10268 0 _0344_
rlabel metal1 24748 22406 24748 22406 0 _0345_
rlabel metal1 13984 4046 13984 4046 0 _0346_
rlabel metal2 18354 4760 18354 4760 0 _0347_
rlabel metal1 20930 2482 20930 2482 0 _0348_
rlabel metal1 20470 4658 20470 4658 0 _0349_
rlabel metal2 6716 22236 6716 22236 0 _0350_
rlabel metal1 16330 16218 16330 16218 0 _0351_
rlabel metal1 7452 20842 7452 20842 0 _0352_
rlabel metal1 18262 8840 18262 8840 0 _0353_
rlabel metal1 10488 3570 10488 3570 0 _0354_
rlabel metal2 11086 5440 11086 5440 0 _0355_
rlabel metal1 6900 14042 6900 14042 0 _0356_
rlabel metal1 16330 8398 16330 8398 0 _0357_
rlabel metal3 1234 28628 1234 28628 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
rlabel metal1 5934 37230 5934 37230 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
rlabel metal2 12788 3910 12788 3910 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
rlabel metal1 23598 2448 23598 2448 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
rlabel metal2 3450 27319 3450 27319 0 ccff_head
rlabel metal3 1234 6868 1234 6868 0 ccff_tail
rlabel via2 37490 30685 37490 30685 0 chanx_left_in[0]
rlabel metal2 11638 1554 11638 1554 0 chanx_left_in[10]
rlabel metal1 25346 37230 25346 37230 0 chanx_left_in[11]
rlabel metal2 38134 8347 38134 8347 0 chanx_left_in[12]
rlabel metal3 1188 748 1188 748 0 chanx_left_in[13]
rlabel metal2 38134 35547 38134 35547 0 chanx_left_in[14]
rlabel metal3 1763 19108 1763 19108 0 chanx_left_in[15]
rlabel metal1 26864 37230 26864 37230 0 chanx_left_in[16]
rlabel metal3 1188 23188 1188 23188 0 chanx_left_in[17]
rlabel metal1 12558 37230 12558 37230 0 chanx_left_in[18]
rlabel metal1 37352 11118 37352 11118 0 chanx_left_in[1]
rlabel metal2 28382 1554 28382 1554 0 chanx_left_in[2]
rlabel metal1 4784 37230 4784 37230 0 chanx_left_in[3]
rlabel metal1 36202 37230 36202 37230 0 chanx_left_in[4]
rlabel metal1 37490 37230 37490 37230 0 chanx_left_in[5]
rlabel metal3 1050 5508 1050 5508 0 chanx_left_in[6]
rlabel metal2 20654 1588 20654 1588 0 chanx_left_in[7]
rlabel via2 37490 27965 37490 27965 0 chanx_left_in[8]
rlabel metal2 38134 12563 38134 12563 0 chanx_left_in[9]
rlabel metal1 15640 37094 15640 37094 0 chanx_left_out[0]
rlabel metal2 39330 1520 39330 1520 0 chanx_left_out[10]
rlabel metal1 33212 37094 33212 37094 0 chanx_left_out[11]
rlabel metal2 17434 1520 17434 1520 0 chanx_left_out[12]
rlabel metal1 3726 37094 3726 37094 0 chanx_left_out[13]
rlabel metal2 10994 1520 10994 1520 0 chanx_left_out[14]
rlabel metal2 2806 14875 2806 14875 0 chanx_left_out[15]
rlabel metal2 25162 1520 25162 1520 0 chanx_left_out[16]
rlabel metal2 38226 13073 38226 13073 0 chanx_left_out[17]
rlabel via2 38226 27285 38226 27285 0 chanx_left_out[18]
rlabel metal2 34822 1520 34822 1520 0 chanx_left_out[1]
rlabel metal2 14858 1520 14858 1520 0 chanx_left_out[2]
rlabel metal1 32384 37094 32384 37094 0 chanx_left_out[3]
rlabel metal1 20148 37094 20148 37094 0 chanx_left_out[4]
rlabel metal2 33534 1792 33534 1792 0 chanx_left_out[5]
rlabel via2 38226 16405 38226 16405 0 chanx_left_out[6]
rlabel metal1 7912 37094 7912 37094 0 chanx_left_out[7]
rlabel metal2 38226 23953 38226 23953 0 chanx_left_out[8]
rlabel metal1 16928 36890 16928 36890 0 chanx_left_out[9]
rlabel metal2 38134 32759 38134 32759 0 chanx_right_in[0]
rlabel metal3 1188 4148 1188 4148 0 chanx_right_in[10]
rlabel metal2 38318 18003 38318 18003 0 chanx_right_in[11]
rlabel metal3 1142 31348 1142 31348 0 chanx_right_in[12]
rlabel metal3 1142 35428 1142 35428 0 chanx_right_in[13]
rlabel metal2 38134 32215 38134 32215 0 chanx_right_in[14]
rlabel metal2 36938 2227 36938 2227 0 chanx_right_in[15]
rlabel metal1 21666 37298 21666 37298 0 chanx_right_in[16]
rlabel metal2 18722 38226 18722 38226 0 chanx_right_in[17]
rlabel metal1 31096 37230 31096 37230 0 chanx_right_in[18]
rlabel metal2 38134 37145 38134 37145 0 chanx_right_in[1]
rlabel metal1 23276 36754 23276 36754 0 chanx_right_in[2]
rlabel metal2 9706 1843 9706 1843 0 chanx_right_in[3]
rlabel metal2 2806 18241 2806 18241 0 chanx_right_in[4]
rlabel metal3 1050 7548 1050 7548 0 chanx_right_in[5]
rlabel metal2 31602 1588 31602 1588 0 chanx_right_in[6]
rlabel metal2 37674 2125 37674 2125 0 chanx_right_in[7]
rlabel metal2 3542 14671 3542 14671 0 chanx_right_in[8]
rlabel metal2 37490 7701 37490 7701 0 chanx_right_in[9]
rlabel metal1 11500 37094 11500 37094 0 chanx_right_out[0]
rlabel metal2 1794 38131 1794 38131 0 chanx_right_out[10]
rlabel metal2 1794 21471 1794 21471 0 chanx_right_out[11]
rlabel metal2 16146 1656 16146 1656 0 chanx_right_out[12]
rlabel metal3 1234 25228 1234 25228 0 chanx_right_out[13]
rlabel metal1 34822 37094 34822 37094 0 chanx_right_out[14]
rlabel metal2 22586 1520 22586 1520 0 chanx_right_out[15]
rlabel metal2 29670 1520 29670 1520 0 chanx_right_out[16]
rlabel via2 38226 24565 38226 24565 0 chanx_right_out[17]
rlabel metal2 38226 4913 38226 4913 0 chanx_right_out[18]
rlabel metal1 27922 37094 27922 37094 0 chanx_right_out[1]
rlabel metal1 37352 36346 37352 36346 0 chanx_right_out[2]
rlabel metal1 17572 37094 17572 37094 0 chanx_right_out[3]
rlabel metal2 690 1792 690 1792 0 chanx_right_out[4]
rlabel metal2 5198 1520 5198 1520 0 chanx_right_out[5]
rlabel metal1 14168 37094 14168 37094 0 chanx_right_out[6]
rlabel metal1 9200 36890 9200 36890 0 chanx_right_out[7]
rlabel metal2 38226 21233 38226 21233 0 chanx_right_out[8]
rlabel metal2 38226 14297 38226 14297 0 chanx_right_out[9]
rlabel metal1 38134 36754 38134 36754 0 chany_bottom_in[0]
rlabel metal1 3220 6766 3220 6766 0 chany_bottom_in[10]
rlabel metal2 38318 2907 38318 2907 0 chany_bottom_in[11]
rlabel metal2 38318 15895 38318 15895 0 chany_bottom_in[12]
rlabel metal2 4094 27659 4094 27659 0 chany_bottom_in[13]
rlabel metal1 2852 37230 2852 37230 0 chany_bottom_in[14]
rlabel metal2 36754 1928 36754 1928 0 chany_bottom_in[15]
rlabel metal2 3726 20349 3726 20349 0 chany_bottom_in[16]
rlabel metal1 3174 36788 3174 36788 0 chany_bottom_in[17]
rlabel metal1 38502 35054 38502 35054 0 chany_bottom_in[18]
rlabel metal2 8418 1707 8418 1707 0 chany_bottom_in[1]
rlabel metal3 1878 18428 1878 18428 0 chany_bottom_in[2]
rlabel metal2 23874 1214 23874 1214 0 chany_bottom_in[3]
rlabel metal2 38042 1367 38042 1367 0 chany_bottom_in[4]
rlabel metal1 13984 37230 13984 37230 0 chany_bottom_in[5]
rlabel metal2 30314 1588 30314 1588 0 chany_bottom_in[6]
rlabel metal1 2162 3570 2162 3570 0 chany_bottom_in[7]
rlabel metal1 2254 8500 2254 8500 0 chany_bottom_in[8]
rlabel via2 38318 4131 38318 4131 0 chany_bottom_in[9]
rlabel metal2 38226 29393 38226 29393 0 chany_bottom_out[0]
rlabel metal2 38226 20621 38226 20621 0 chany_bottom_out[10]
rlabel metal2 32890 1520 32890 1520 0 chany_bottom_out[11]
rlabel metal3 1234 23868 1234 23868 0 chany_bottom_out[12]
rlabel metal2 38226 9741 38226 9741 0 chany_bottom_out[13]
rlabel metal3 1234 32028 1234 32028 0 chany_bottom_out[14]
rlabel via2 38226 22491 38226 22491 0 chany_bottom_out[15]
rlabel metal2 38226 34221 38226 34221 0 chany_bottom_out[16]
rlabel metal2 36110 1520 36110 1520 0 chany_bottom_out[17]
rlabel metal2 38226 36057 38226 36057 0 chany_bottom_out[18]
rlabel metal3 1234 33388 1234 33388 0 chany_bottom_out[1]
rlabel metal3 1602 2108 1602 2108 0 chany_bottom_out[2]
rlabel metal1 5980 12614 5980 12614 0 chany_bottom_out[3]
rlabel metal2 46 1656 46 1656 0 chany_bottom_out[4]
rlabel metal2 25806 1520 25806 1520 0 chany_bottom_out[5]
rlabel metal1 1748 36890 1748 36890 0 chany_bottom_out[6]
rlabel metal1 9844 37094 9844 37094 0 chany_bottom_out[7]
rlabel metal1 24656 37094 24656 37094 0 chany_bottom_out[8]
rlabel metal3 1234 29988 1234 29988 0 chany_bottom_out[9]
rlabel metal1 15870 13192 15870 13192 0 clknet_0_prog_clk
rlabel metal2 1610 5168 1610 5168 0 clknet_4_0_0_prog_clk
rlabel metal1 1794 17102 1794 17102 0 clknet_4_10_0_prog_clk
rlabel metal1 5934 18156 5934 18156 0 clknet_4_11_0_prog_clk
rlabel metal1 7498 12852 7498 12852 0 clknet_4_12_0_prog_clk
rlabel metal1 14444 12274 14444 12274 0 clknet_4_13_0_prog_clk
rlabel metal2 6854 14382 6854 14382 0 clknet_4_14_0_prog_clk
rlabel metal2 9062 14688 9062 14688 0 clknet_4_15_0_prog_clk
rlabel metal1 6624 7310 6624 7310 0 clknet_4_1_0_prog_clk
rlabel metal1 1978 8398 1978 8398 0 clknet_4_2_0_prog_clk
rlabel metal1 6486 9996 6486 9996 0 clknet_4_3_0_prog_clk
rlabel metal2 9062 7072 9062 7072 0 clknet_4_4_0_prog_clk
rlabel metal1 14030 2482 14030 2482 0 clknet_4_5_0_prog_clk
rlabel metal2 9798 10948 9798 10948 0 clknet_4_6_0_prog_clk
rlabel metal1 15824 10098 15824 10098 0 clknet_4_7_0_prog_clk
rlabel metal1 2070 11798 2070 11798 0 clknet_4_8_0_prog_clk
rlabel metal1 4140 12614 4140 12614 0 clknet_4_9_0_prog_clk
rlabel metal1 4692 4046 4692 4046 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal2 1978 1928 1978 1928 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal2 4002 8721 4002 8721 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 22172 36754 22172 36754 0 left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 27370 2074 27370 2074 0 left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 35604 36754 35604 36754 0 left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 38318 6239 38318 6239 0 left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal3 1602 36788 1602 36788 0 left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal2 2806 10285 2806 10285 0 left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal2 7130 1761 7130 1761 0 left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal1 16698 5066 16698 5066 0 mem_bottom_track_1.DFFR_0_.D
rlabel metal1 15594 6086 15594 6086 0 mem_bottom_track_1.DFFR_0_.Q
rlabel metal1 16284 6902 16284 6902 0 mem_bottom_track_1.DFFR_1_.Q
rlabel metal2 16468 14790 16468 14790 0 mem_bottom_track_1.DFFR_2_.Q
rlabel metal1 15870 8262 15870 8262 0 mem_bottom_track_1.DFFR_3_.Q
rlabel metal1 17572 1938 17572 1938 0 mem_bottom_track_1.DFFR_4_.Q
rlabel metal1 16422 2618 16422 2618 0 mem_bottom_track_1.DFFR_5_.Q
rlabel metal1 10810 3400 10810 3400 0 mem_bottom_track_11.DFFR_0_.D
rlabel metal1 19458 14994 19458 14994 0 mem_bottom_track_11.DFFR_0_.Q
rlabel metal1 15916 7718 15916 7718 0 mem_bottom_track_11.DFFR_1_.Q
rlabel metal2 14306 13112 14306 13112 0 mem_bottom_track_13.DFFR_0_.Q
rlabel metal2 9062 17272 9062 17272 0 mem_bottom_track_13.DFFR_1_.Q
rlabel metal2 21298 14688 21298 14688 0 mem_bottom_track_15.DFFR_0_.Q
rlabel metal1 14122 25874 14122 25874 0 mem_bottom_track_15.DFFR_1_.Q
rlabel metal1 13248 21522 13248 21522 0 mem_bottom_track_17.DFFR_0_.Q
rlabel metal1 15594 25296 15594 25296 0 mem_bottom_track_17.DFFR_1_.Q
rlabel metal1 15870 19822 15870 19822 0 mem_bottom_track_19.DFFR_0_.Q
rlabel metal1 1656 12274 1656 12274 0 mem_bottom_track_19.DFFR_1_.Q
rlabel metal1 11638 17102 11638 17102 0 mem_bottom_track_21.DFFR_0_.Q
rlabel via2 19918 17595 19918 17595 0 mem_bottom_track_21.DFFR_1_.Q
rlabel metal2 27094 13821 27094 13821 0 mem_bottom_track_23.DFFR_0_.Q
rlabel metal1 11730 8058 11730 8058 0 mem_bottom_track_23.DFFR_1_.Q
rlabel metal1 15088 12818 15088 12818 0 mem_bottom_track_25.DFFR_0_.Q
rlabel metal1 11776 13226 11776 13226 0 mem_bottom_track_25.DFFR_1_.Q
rlabel metal1 14628 16490 14628 16490 0 mem_bottom_track_27.DFFR_0_.Q
rlabel metal1 16008 16422 16008 16422 0 mem_bottom_track_27.DFFR_1_.Q
rlabel metal1 18170 19856 18170 19856 0 mem_bottom_track_3.DFFR_0_.Q
rlabel metal1 15870 16626 15870 16626 0 mem_bottom_track_3.DFFR_1_.Q
rlabel via3 9131 16388 9131 16388 0 mem_bottom_track_3.DFFR_2_.Q
rlabel metal1 4600 17238 4600 17238 0 mem_bottom_track_3.DFFR_3_.Q
rlabel metal1 1932 14314 1932 14314 0 mem_bottom_track_3.DFFR_4_.Q
rlabel metal1 3404 14586 3404 14586 0 mem_bottom_track_3.DFFR_5_.Q
rlabel metal2 12650 27676 12650 27676 0 mem_bottom_track_37.DFFR_0_.Q
rlabel via3 13179 12444 13179 12444 0 mem_bottom_track_37.DFFR_1_.Q
rlabel via2 17342 17629 17342 17629 0 mem_bottom_track_5.DFFR_0_.Q
rlabel metal1 5382 17850 5382 17850 0 mem_bottom_track_5.DFFR_1_.Q
rlabel metal2 6394 14960 6394 14960 0 mem_bottom_track_5.DFFR_2_.Q
rlabel metal2 1886 26401 1886 26401 0 mem_bottom_track_5.DFFR_3_.Q
rlabel metal1 1886 7922 1886 7922 0 mem_bottom_track_5.DFFR_4_.Q
rlabel metal3 1127 24956 1127 24956 0 mem_bottom_track_5.DFFR_5_.Q
rlabel metal2 5152 13124 5152 13124 0 mem_bottom_track_7.DFFR_0_.Q
rlabel metal2 1886 13226 1886 13226 0 mem_bottom_track_7.DFFR_1_.Q
rlabel metal2 3358 15555 3358 15555 0 mem_bottom_track_7.DFFR_2_.Q
rlabel metal1 3726 15878 3726 15878 0 mem_bottom_track_7.DFFR_3_.Q
rlabel metal1 1886 10608 1886 10608 0 mem_bottom_track_7.DFFR_4_.Q
rlabel metal2 2530 27149 2530 27149 0 mem_bottom_track_7.DFFR_5_.Q
rlabel metal2 12558 14059 12558 14059 0 mem_bottom_track_9.DFFR_0_.Q
rlabel metal2 15042 10353 15042 10353 0 mem_left_track_1.DFFR_0_.Q
rlabel metal1 12742 10200 12742 10200 0 mem_left_track_1.DFFR_1_.Q
rlabel metal1 2622 23766 2622 23766 0 mem_left_track_1.DFFR_2_.Q
rlabel metal2 5612 13940 5612 13940 0 mem_left_track_1.DFFR_3_.Q
rlabel metal1 7268 11526 7268 11526 0 mem_left_track_1.DFFR_4_.Q
rlabel metal1 7084 14450 7084 14450 0 mem_left_track_1.DFFR_5_.Q
rlabel metal1 8602 9418 8602 9418 0 mem_left_track_17.DFFR_0_.D
rlabel metal1 20792 16082 20792 16082 0 mem_left_track_17.DFFR_0_.Q
rlabel metal2 12742 7684 12742 7684 0 mem_left_track_17.DFFR_1_.Q
rlabel metal1 19458 13906 19458 13906 0 mem_left_track_17.DFFR_2_.Q
rlabel metal2 16054 5236 16054 5236 0 mem_left_track_17.DFFR_3_.Q
rlabel metal2 12466 5984 12466 5984 0 mem_left_track_17.DFFR_4_.Q
rlabel metal2 13294 5253 13294 5253 0 mem_left_track_17.DFFR_5_.Q
rlabel metal1 18446 4216 18446 4216 0 mem_left_track_17.DFFR_6_.Q
rlabel metal1 19918 5746 19918 5746 0 mem_left_track_17.DFFR_7_.Q
rlabel metal1 10258 16082 10258 16082 0 mem_left_track_25.DFFR_0_.Q
rlabel metal2 13846 16065 13846 16065 0 mem_left_track_25.DFFR_1_.Q
rlabel metal2 12558 23970 12558 23970 0 mem_left_track_25.DFFR_2_.Q
rlabel metal2 18354 22661 18354 22661 0 mem_left_track_25.DFFR_3_.Q
rlabel metal2 8970 11390 8970 11390 0 mem_left_track_25.DFFR_4_.Q
rlabel metal1 6900 6834 6900 6834 0 mem_left_track_25.DFFR_5_.Q
rlabel metal1 5658 4998 5658 4998 0 mem_left_track_25.DFFR_6_.Q
rlabel via2 13018 3893 13018 3893 0 mem_left_track_25.DFFR_7_.Q
rlabel metal2 12650 7123 12650 7123 0 mem_left_track_33.DFFR_0_.Q
rlabel metal2 18078 6732 18078 6732 0 mem_left_track_33.DFFR_1_.Q
rlabel metal2 19274 4284 19274 4284 0 mem_left_track_33.DFFR_2_.Q
rlabel metal1 8050 3910 8050 3910 0 mem_left_track_33.DFFR_3_.Q
rlabel metal1 12650 4046 12650 4046 0 mem_left_track_33.DFFR_4_.Q
rlabel metal2 15042 20434 15042 20434 0 mem_left_track_9.DFFR_0_.Q
rlabel metal1 11592 21522 11592 21522 0 mem_left_track_9.DFFR_1_.Q
rlabel metal1 20562 14994 20562 14994 0 mem_left_track_9.DFFR_2_.Q
rlabel metal1 18998 25262 18998 25262 0 mem_left_track_9.DFFR_3_.Q
rlabel metal1 11224 14450 11224 14450 0 mem_left_track_9.DFFR_4_.Q
rlabel metal1 8694 17782 8694 17782 0 mem_left_track_9.DFFR_5_.Q
rlabel metal3 6647 21964 6647 21964 0 mem_left_track_9.DFFR_6_.Q
rlabel metal2 12650 23902 12650 23902 0 mem_right_track_0.DFFR_0_.Q
rlabel metal1 5612 17102 5612 17102 0 mem_right_track_0.DFFR_1_.Q
rlabel metal1 9236 14790 9236 14790 0 mem_right_track_0.DFFR_2_.Q
rlabel metal1 10350 14892 10350 14892 0 mem_right_track_0.DFFR_3_.Q
rlabel metal1 4370 15538 4370 15538 0 mem_right_track_0.DFFR_4_.Q
rlabel metal1 6118 15538 6118 15538 0 mem_right_track_0.DFFR_5_.Q
rlabel metal2 3726 18343 3726 18343 0 mem_right_track_0.DFFR_6_.Q
rlabel metal1 8050 18190 8050 18190 0 mem_right_track_0.DFFR_7_.Q
rlabel metal1 10120 8874 10120 8874 0 mem_right_track_16.DFFR_0_.D
rlabel metal3 7544 19380 7544 19380 0 mem_right_track_16.DFFR_0_.Q
rlabel metal1 22034 13872 22034 13872 0 mem_right_track_16.DFFR_1_.Q
rlabel metal1 13754 8500 13754 8500 0 mem_right_track_16.DFFR_2_.Q
rlabel metal1 13754 8330 13754 8330 0 mem_right_track_16.DFFR_3_.Q
rlabel metal2 15778 9282 15778 9282 0 mem_right_track_16.DFFR_4_.Q
rlabel metal1 16054 9044 16054 9044 0 mem_right_track_16.DFFR_5_.Q
rlabel via2 14582 12155 14582 12155 0 mem_right_track_16.DFFR_6_.Q
rlabel metal2 20102 12818 20102 12818 0 mem_right_track_16.DFFR_7_.Q
rlabel metal2 12558 14926 12558 14926 0 mem_right_track_24.DFFR_0_.Q
rlabel metal1 14214 17238 14214 17238 0 mem_right_track_24.DFFR_1_.Q
rlabel metal1 16100 16966 16100 16966 0 mem_right_track_24.DFFR_2_.Q
rlabel metal1 13156 19346 13156 19346 0 mem_right_track_24.DFFR_3_.Q
rlabel metal1 8510 10472 8510 10472 0 mem_right_track_24.DFFR_4_.Q
rlabel metal2 17250 7939 17250 7939 0 mem_right_track_24.DFFR_5_.Q
rlabel metal2 14490 9180 14490 9180 0 mem_right_track_24.DFFR_6_.Q
rlabel metal2 13478 3400 13478 3400 0 mem_right_track_24.DFFR_7_.Q
rlabel metal1 15042 2822 15042 2822 0 mem_right_track_32.DFFR_0_.Q
rlabel metal1 20746 15368 20746 15368 0 mem_right_track_32.DFFR_1_.Q
rlabel metal1 14444 3434 14444 3434 0 mem_right_track_32.DFFR_2_.Q
rlabel metal2 16054 3842 16054 3842 0 mem_right_track_32.DFFR_3_.Q
rlabel metal1 17572 5542 17572 5542 0 mem_right_track_32.DFFR_4_.Q
rlabel metal1 18860 19142 18860 19142 0 mem_right_track_8.DFFR_0_.Q
rlabel metal1 8050 13498 8050 13498 0 mem_right_track_8.DFFR_1_.Q
rlabel metal2 12558 17782 12558 17782 0 mem_right_track_8.DFFR_2_.Q
rlabel metal1 16974 22610 16974 22610 0 mem_right_track_8.DFFR_3_.Q
rlabel metal1 4876 9486 4876 9486 0 mem_right_track_8.DFFR_4_.Q
rlabel metal1 13938 15096 13938 15096 0 mem_right_track_8.DFFR_5_.Q
rlabel metal1 12466 9553 12466 9553 0 mem_right_track_8.DFFR_6_.Q
rlabel metal1 20562 17034 20562 17034 0 mux_bottom_track_1.INVTX1_0_.out
rlabel metal1 16146 11662 16146 11662 0 mux_bottom_track_1.INVTX1_1_.out
rlabel metal1 20194 19890 20194 19890 0 mux_bottom_track_1.INVTX1_2_.out
rlabel metal1 16974 5304 16974 5304 0 mux_bottom_track_1.INVTX1_3_.out
rlabel metal1 19642 17000 19642 17000 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 37398 26962 37398 26962 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 37582 27268 37582 27268 0 mux_bottom_track_1.out
rlabel metal1 21482 10540 21482 10540 0 mux_bottom_track_11.INVTX1_0_.out
rlabel metal2 16238 17442 16238 17442 0 mux_bottom_track_11.INVTX1_1_.out
rlabel metal2 21068 13804 21068 13804 0 mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 22770 7378 22770 7378 0 mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 22356 3026 22356 3026 0 mux_bottom_track_11.out
rlabel metal2 12282 24514 12282 24514 0 mux_bottom_track_13.INVTX1_0_.out
rlabel metal1 17986 22542 17986 22542 0 mux_bottom_track_13.INVTX1_1_.out
rlabel metal1 16008 24242 16008 24242 0 mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 8326 27846 8326 27846 0 mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 5152 34578 5152 34578 0 mux_bottom_track_13.out
rlabel metal1 19550 11016 19550 11016 0 mux_bottom_track_15.INVTX1_0_.out
rlabel metal1 19642 12750 19642 12750 0 mux_bottom_track_15.INVTX1_1_.out
rlabel metal2 18446 11696 18446 11696 0 mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 12374 32878 12374 32878 0 mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 10810 32572 10810 32572 0 mux_bottom_track_15.out
rlabel metal1 15456 20774 15456 20774 0 mux_bottom_track_17.INVTX1_0_.out
rlabel metal1 13708 20366 13708 20366 0 mux_bottom_track_17.INVTX1_1_.out
rlabel metal1 14812 20910 14812 20910 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 16974 26656 16974 26656 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 21804 33966 21804 33966 0 mux_bottom_track_17.out
rlabel metal2 7268 24004 7268 24004 0 mux_bottom_track_19.INVTX1_0_.out
rlabel metal1 17894 18598 17894 18598 0 mux_bottom_track_19.INVTX1_2_.out
rlabel metal1 6164 25262 6164 25262 0 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 15318 19210 15318 19210 0 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 7774 24854 7774 24854 0 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 7360 26010 7360 26010 0 mux_bottom_track_19.out
rlabel metal2 9430 21335 9430 21335 0 mux_bottom_track_21.INVTX1_0_.out
rlabel metal1 4876 18938 4876 18938 0 mux_bottom_track_21.INVTX1_1_.out
rlabel metal2 17250 18904 17250 18904 0 mux_bottom_track_21.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 34546 19244 34546 19244 0 mux_bottom_track_21.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 37490 19822 37490 19822 0 mux_bottom_track_21.out
rlabel metal1 23092 21454 23092 21454 0 mux_bottom_track_23.INVTX1_0_.out
rlabel metal2 17986 20587 17986 20587 0 mux_bottom_track_23.INVTX1_1_.out
rlabel metal1 22264 13498 22264 13498 0 mux_bottom_track_23.INVTX1_2_.out
rlabel metal1 23690 20774 23690 20774 0 mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 25944 14586 25944 14586 0 mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 26450 12925 26450 12925 0 mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 30406 5236 30406 5236 0 mux_bottom_track_23.out
rlabel metal1 19366 19482 19366 19482 0 mux_bottom_track_25.INVTX1_0_.out
rlabel metal1 3312 20366 3312 20366 0 mux_bottom_track_25.INVTX1_1_.out
rlabel metal2 22126 25398 22126 25398 0 mux_bottom_track_25.INVTX1_2_.out
rlabel metal2 12098 26996 12098 26996 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 17066 28662 17066 28662 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 12466 25092 12466 25092 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 7176 23834 7176 23834 0 mux_bottom_track_25.out
rlabel metal1 17572 24310 17572 24310 0 mux_bottom_track_27.INVTX1_0_.out
rlabel metal1 25438 26894 25438 26894 0 mux_bottom_track_27.INVTX1_1_.out
rlabel metal1 26128 17306 26128 17306 0 mux_bottom_track_27.INVTX1_2_.out
rlabel metal1 23874 19686 23874 19686 0 mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 27554 18326 27554 18326 0 mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 27646 16762 27646 16762 0 mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 30406 14654 30406 14654 0 mux_bottom_track_27.out
rlabel metal2 16698 20060 16698 20060 0 mux_bottom_track_3.INVTX1_0_.out
rlabel metal2 14674 11339 14674 11339 0 mux_bottom_track_3.INVTX1_1_.out
rlabel metal1 19458 21012 19458 21012 0 mux_bottom_track_3.INVTX1_3_.out
rlabel metal1 21114 31858 21114 31858 0 mux_bottom_track_3.INVTX1_4_.out
rlabel metal1 18998 20774 18998 20774 0 mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem2_0_out
rlabel metal2 17342 18513 17342 18513 0 mux_bottom_track_3.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 9660 22066 9660 22066 0 mux_bottom_track_3.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 5842 28900 5842 28900 0 mux_bottom_track_3.out
rlabel metal1 9016 33286 9016 33286 0 mux_bottom_track_37.INVTX1_1_.out
rlabel metal1 14674 26996 14674 26996 0 mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 17802 27030 17802 27030 0 mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 31970 32878 31970 32878 0 mux_bottom_track_37.out
rlabel metal1 21022 19720 21022 19720 0 mux_bottom_track_5.INVTX1_0_.out
rlabel metal2 15042 17170 15042 17170 0 mux_bottom_track_5.INVTX1_3_.out
rlabel metal1 1748 23018 1748 23018 0 mux_bottom_track_5.INVTX1_4_.out
rlabel metal1 15870 17782 15870 17782 0 mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem2_0_out
rlabel metal1 1794 21420 1794 21420 0 mux_bottom_track_5.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 2116 6290 2116 6290 0 mux_bottom_track_5.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 1978 6596 1978 6596 0 mux_bottom_track_5.out
rlabel metal2 12558 19278 12558 19278 0 mux_bottom_track_7.INVTX1_0_.out
rlabel metal1 13478 18156 13478 18156 0 mux_bottom_track_7.INVTX1_2_.out
rlabel metal1 8464 19142 8464 19142 0 mux_bottom_track_7.INVTX1_3_.out
rlabel metal2 12834 19856 12834 19856 0 mux_bottom_track_7.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 2024 21998 2024 21998 0 mux_bottom_track_7.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 1978 22066 1978 22066 0 mux_bottom_track_7.out
rlabel metal1 19964 10574 19964 10574 0 mux_bottom_track_9.INVTX1_0_.out
rlabel metal2 17802 14552 17802 14552 0 mux_bottom_track_9.INVTX1_1_.out
rlabel metal1 17664 14246 17664 14246 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 17250 2924 17250 2924 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 3542 6256 3542 6256 0 mux_bottom_track_9.out
rlabel metal2 21160 9690 21160 9690 0 mux_left_track_1.INVTX1_3_.out
rlabel metal2 21022 8738 21022 8738 0 mux_left_track_1.INVTX1_4_.out
rlabel metal2 14398 19703 14398 19703 0 mux_left_track_1.INVTX1_5_.out
rlabel metal2 2070 15368 2070 15368 0 mux_left_track_1.INVTX1_6_.out
rlabel metal2 5290 21529 5290 21529 0 mux_left_track_1.INVTX1_7_.out
rlabel metal2 17710 18496 17710 18496 0 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 15042 19635 15042 19635 0 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 3634 21692 3634 21692 0 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 13570 19159 13570 19159 0 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 14628 36754 14628 36754 0 mux_left_track_1.out
rlabel metal1 17020 5746 17020 5746 0 mux_left_track_17.INVTX1_3_.out
rlabel metal1 21528 7786 21528 7786 0 mux_left_track_17.INVTX1_4_.out
rlabel via2 26266 7939 26266 7939 0 mux_left_track_17.INVTX1_5_.out
rlabel metal2 17710 14637 17710 14637 0 mux_left_track_17.INVTX1_6_.out
rlabel metal2 14214 4828 14214 4828 0 mux_left_track_17.INVTX1_7_.out
rlabel metal2 18814 2210 18814 2210 0 mux_left_track_17.INVTX1_8_.out
rlabel metal1 19826 19278 19826 19278 0 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 17756 13124 17756 13124 0 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 21298 12789 21298 12789 0 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 36846 19958 36846 19958 0 mux_left_track_17.out
rlabel metal1 4048 18190 4048 18190 0 mux_left_track_25.INVTX1_3_.out
rlabel metal1 6302 3978 6302 3978 0 mux_left_track_25.INVTX1_4_.out
rlabel metal1 19826 16626 19826 16626 0 mux_left_track_25.INVTX1_5_.out
rlabel metal1 9614 23154 9614 23154 0 mux_left_track_25.INVTX1_6_.out
rlabel metal1 27968 31858 27968 31858 0 mux_left_track_25.INVTX1_7_.out
rlabel metal2 20102 3009 20102 3009 0 mux_left_track_25.INVTX1_8_.out
rlabel metal1 10488 21318 10488 21318 0 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 17802 10982 17802 10982 0 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 16238 10472 16238 10472 0 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 24794 2992 24794 2992 0 mux_left_track_25.out
rlabel metal2 18170 8738 18170 8738 0 mux_left_track_33.INVTX1_2_.out
rlabel metal2 2898 27251 2898 27251 0 mux_left_track_33.INVTX1_3_.out
rlabel metal1 6302 22066 6302 22066 0 mux_left_track_33.INVTX1_4_.out
rlabel metal2 17342 20910 17342 20910 0 mux_left_track_33.INVTX1_5_.out
rlabel metal2 16514 5661 16514 5661 0 mux_left_track_33.INVTX1_6_.out
rlabel metal2 14490 1836 14490 1836 0 mux_left_track_33.INVTX1_7_.out
rlabel metal2 18032 17068 18032 17068 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 18170 19805 18170 19805 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 18262 4828 18262 4828 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 17986 6834 17986 6834 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 22126 2414 22126 2414 0 mux_left_track_33.out
rlabel metal1 17756 24718 17756 24718 0 mux_left_track_9.INVTX1_3_.out
rlabel metal2 13386 27642 13386 27642 0 mux_left_track_9.INVTX1_4_.out
rlabel metal1 14122 13226 14122 13226 0 mux_left_track_9.INVTX1_5_.out
rlabel metal2 20654 11866 20654 11866 0 mux_left_track_9.INVTX1_6_.out
rlabel metal1 20746 32198 20746 32198 0 mux_left_track_9.INVTX1_7_.out
rlabel metal1 2392 25942 2392 25942 0 mux_left_track_9.INVTX1_8_.out
rlabel metal1 16238 20502 16238 20502 0 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 15824 21590 15824 21590 0 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 19458 29036 19458 29036 0 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 19964 36142 19964 36142 0 mux_left_track_9.out
rlabel metal1 21758 31994 21758 31994 0 mux_right_track_0.INVTX1_0_.out
rlabel metal1 1610 20536 1610 20536 0 mux_right_track_0.INVTX1_1_.out
rlabel metal1 18492 21454 18492 21454 0 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 20194 20604 20194 20604 0 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 6026 20536 6026 20536 0 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 8832 30906 8832 30906 0 mux_right_track_0.out
rlabel metal1 8556 30634 8556 30634 0 mux_right_track_16.INVTX1_0_.out
rlabel metal1 22586 16014 22586 16014 0 mux_right_track_16.INVTX1_1_.out
rlabel metal1 13110 19924 13110 19924 0 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 20424 12750 20424 12750 0 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 21482 16048 21482 16048 0 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 31418 21318 31418 21318 0 mux_right_track_16.out
rlabel metal1 9936 32742 9936 32742 0 mux_right_track_24.INVTX1_0_.out
rlabel metal2 31142 22168 31142 22168 0 mux_right_track_24.INVTX1_1_.out
rlabel metal1 17848 21454 17848 21454 0 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 14398 18734 14398 18734 0 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 22402 16932 22402 16932 0 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 13570 1938 13570 1938 0 mux_right_track_24.out
rlabel metal2 20194 5814 20194 5814 0 mux_right_track_32.INVTX1_0_.out
rlabel metal2 15686 6137 15686 6137 0 mux_right_track_32.INVTX1_1_.out
rlabel metal1 22816 6222 22816 6222 0 mux_right_track_32.mux_2level_tapbuf_basis_input2_mem2_0_out
rlabel metal1 17388 5882 17388 5882 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 20056 14314 20056 14314 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 23230 5984 23230 5984 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 26450 5372 26450 5372 0 mux_right_track_32.out
rlabel metal2 23598 32062 23598 32062 0 mux_right_track_8.INVTX1_0_.out
rlabel metal1 4738 30022 4738 30022 0 mux_right_track_8.INVTX1_1_.out
rlabel metal1 6532 19278 6532 19278 0 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 20516 16490 20516 16490 0 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 16146 15572 16146 15572 0 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 3450 4726 3450 4726 0 mux_right_track_8.out
rlabel metal2 4738 26809 4738 26809 0 net1
rlabel metal1 1656 2618 1656 2618 0 net10
rlabel metal2 38042 16286 38042 16286 0 net100
rlabel metal1 17158 36856 17158 36856 0 net101
rlabel metal2 37766 22372 37766 22372 0 net102
rlabel metal2 16882 33014 16882 33014 0 net103
rlabel metal1 10626 37162 10626 37162 0 net104
rlabel metal1 2024 37230 2024 37230 0 net105
rlabel metal1 1932 20910 1932 20910 0 net106
rlabel metal2 18262 2244 18262 2244 0 net107
rlabel via2 2254 25245 2254 25245 0 net108
rlabel metal1 34868 37230 34868 37230 0 net109
rlabel metal1 37950 35462 37950 35462 0 net11
rlabel metal2 22678 2040 22678 2040 0 net110
rlabel metal1 29624 2414 29624 2414 0 net111
rlabel metal2 32706 24310 32706 24310 0 net112
rlabel metal1 37996 5202 37996 5202 0 net113
rlabel metal1 26956 30906 26956 30906 0 net114
rlabel metal1 37950 21114 37950 21114 0 net115
rlabel metal1 18308 37162 18308 37162 0 net116
rlabel metal1 2070 3026 2070 3026 0 net117
rlabel metal3 6371 2652 6371 2652 0 net118
rlabel metal2 14306 36924 14306 36924 0 net119
rlabel via3 1909 19244 1909 19244 0 net12
rlabel metal2 9154 34247 9154 34247 0 net120
rlabel metal1 36961 21522 36961 21522 0 net121
rlabel metal1 37904 21862 37904 21862 0 net122
rlabel metal2 37398 28594 37398 28594 0 net123
rlabel metal1 37904 20026 37904 20026 0 net124
rlabel metal1 33350 2414 33350 2414 0 net125
rlabel metal1 1610 24276 1610 24276 0 net126
rlabel metal2 36938 11594 36938 11594 0 net127
rlabel metal2 2254 32096 2254 32096 0 net128
rlabel metal2 37858 21046 37858 21046 0 net129
rlabel metal1 30130 37298 30130 37298 0 net13
rlabel metal1 38042 18938 38042 18938 0 net130
rlabel metal1 36041 2414 36041 2414 0 net131
rlabel metal1 38042 36108 38042 36108 0 net132
rlabel metal1 2852 33490 2852 33490 0 net133
rlabel metal1 2300 6630 2300 6630 0 net134
rlabel metal1 1380 24582 1380 24582 0 net135
rlabel metal1 3220 6086 3220 6086 0 net136
rlabel metal1 25944 2414 25944 2414 0 net137
rlabel metal1 2852 36686 2852 36686 0 net138
rlabel metal1 10212 32538 10212 32538 0 net139
rlabel metal2 12742 24514 12742 24514 0 net14
rlabel metal1 23230 37162 23230 37162 0 net140
rlabel metal1 1610 30192 1610 30192 0 net141
rlabel metal2 7038 24480 7038 24480 0 net142
rlabel metal1 20010 6834 20010 6834 0 net143
rlabel metal2 20470 14110 20470 14110 0 net144
rlabel metal1 17710 6188 17710 6188 0 net145
rlabel metal2 7498 22814 7498 22814 0 net146
rlabel metal1 21114 7922 21114 7922 0 net147
rlabel metal1 15686 3128 15686 3128 0 net148
rlabel metal1 22494 9690 22494 9690 0 net149
rlabel metal2 12466 33898 12466 33898 0 net15
rlabel metal2 24978 9758 24978 9758 0 net150
rlabel metal1 2760 18802 2760 18802 0 net151
rlabel metal2 2898 23902 2898 23902 0 net152
rlabel metal1 2760 20978 2760 20978 0 net153
rlabel metal1 6946 3672 6946 3672 0 net154
rlabel metal2 20838 7888 20838 7888 0 net155
rlabel metal1 8096 24786 8096 24786 0 net156
rlabel metal1 12650 25194 12650 25194 0 net157
rlabel metal2 16330 25568 16330 25568 0 net158
rlabel metal2 24702 19040 24702 19040 0 net159
rlabel metal1 37490 20910 37490 20910 0 net16
rlabel metal2 17802 26078 17802 26078 0 net160
rlabel metal2 14398 24684 14398 24684 0 net161
rlabel metal2 25990 14688 25990 14688 0 net162
rlabel metal2 16974 28356 16974 28356 0 net163
rlabel metal1 26312 19822 26312 19822 0 net164
rlabel metal2 2438 23392 2438 23392 0 net165
rlabel metal1 21390 4522 21390 4522 0 net166
rlabel metal1 17250 17170 17250 17170 0 net17
rlabel metal2 4738 35292 4738 35292 0 net18
rlabel metal2 36386 27744 36386 27744 0 net19
rlabel metal1 6118 37094 6118 37094 0 net2
rlabel metal1 18630 36754 18630 36754 0 net20
rlabel metal1 1886 5066 1886 5066 0 net21
rlabel metal1 21298 2618 21298 2618 0 net22
rlabel metal2 38042 22372 38042 22372 0 net23
rlabel metal2 38226 12665 38226 12665 0 net24
rlabel metal2 38180 29580 38180 29580 0 net25
rlabel metal1 1978 4114 1978 4114 0 net26
rlabel metal1 38088 18394 38088 18394 0 net27
rlabel metal1 3772 27098 3772 27098 0 net28
rlabel metal1 4692 35598 4692 35598 0 net29
rlabel metal2 18078 5440 18078 5440 0 net3
rlabel metal1 38088 32198 38088 32198 0 net30
rlabel metal2 30590 10234 30590 10234 0 net31
rlabel metal1 21896 37230 21896 37230 0 net32
rlabel metal1 18722 37298 18722 37298 0 net33
rlabel metal1 29670 37162 29670 37162 0 net34
rlabel metal1 38364 36618 38364 36618 0 net35
rlabel metal1 22862 36686 22862 36686 0 net36
rlabel metal2 2714 2397 2714 2397 0 net37
rlabel metal1 10810 13906 10810 13906 0 net38
rlabel via2 1886 7259 1886 7259 0 net39
rlabel via2 23414 2533 23414 2533 0 net4
rlabel metal1 28382 2482 28382 2482 0 net40
rlabel metal1 37582 18734 37582 18734 0 net41
rlabel metal1 16882 29138 16882 29138 0 net42
rlabel metal1 37904 4590 37904 4590 0 net43
rlabel metal1 34960 36618 34960 36618 0 net44
rlabel metal1 7314 5678 7314 5678 0 net45
rlabel metal1 38134 2924 38134 2924 0 net46
rlabel metal2 29762 15674 29762 15674 0 net47
rlabel metal1 5152 22610 5152 22610 0 net48
rlabel metal1 4784 37162 4784 37162 0 net49
rlabel metal4 1012 20604 1012 20604 0 net5
rlabel metal2 27186 5270 27186 5270 0 net50
rlabel metal1 4094 26384 4094 26384 0 net51
rlabel metal1 4416 36550 4416 36550 0 net52
rlabel metal2 37306 32878 37306 32878 0 net53
rlabel metal2 15686 6528 15686 6528 0 net54
rlabel metal2 2622 10438 2622 10438 0 net55
rlabel metal1 21298 6732 21298 6732 0 net56
rlabel metal2 38134 4420 38134 4420 0 net57
rlabel metal1 13248 37094 13248 37094 0 net58
rlabel metal1 30314 2618 30314 2618 0 net59
rlabel metal1 36823 30770 36823 30770 0 net6
rlabel metal2 6578 3910 6578 3910 0 net60
rlabel via2 1610 8619 1610 8619 0 net61
rlabel metal2 31418 6766 31418 6766 0 net62
rlabel metal2 4002 3468 4002 3468 0 net63
rlabel metal2 4922 4522 4922 4522 0 net64
rlabel metal2 1978 8772 1978 8772 0 net65
rlabel metal1 21390 36550 21390 36550 0 net66
rlabel metal2 27186 2329 27186 2329 0 net67
rlabel metal1 31786 31790 31786 31790 0 net68
rlabel metal1 37007 6426 37007 6426 0 net69
rlabel metal1 11592 2618 11592 2618 0 net7
rlabel metal2 2346 33626 2346 33626 0 net70
rlabel metal3 1863 18972 1863 18972 0 net71
rlabel metal1 3956 3366 3956 3366 0 net72
rlabel metal1 18032 10030 18032 10030 0 net73
rlabel metal2 34546 25330 34546 25330 0 net74
rlabel metal2 22678 3332 22678 3332 0 net75
rlabel metal1 28198 36210 28198 36210 0 net76
rlabel metal1 26082 32402 26082 32402 0 net77
rlabel metal1 2116 36006 2116 36006 0 net78
rlabel metal2 6578 34986 6578 34986 0 net79
rlabel metal1 24932 31858 24932 31858 0 net8
rlabel metal1 26542 4590 26542 4590 0 net80
rlabel via2 2622 28067 2622 28067 0 net81
rlabel metal2 2714 32572 2714 32572 0 net82
rlabel metal2 38134 18428 38134 18428 0 net83
rlabel metal2 1610 6324 1610 6324 0 net84
rlabel metal2 14858 37060 14858 37060 0 net85
rlabel metal2 38042 3434 38042 3434 0 net86
rlabel metal1 32752 37230 32752 37230 0 net87
rlabel metal1 19826 2516 19826 2516 0 net88
rlabel metal1 3588 35258 3588 35258 0 net89
rlabel metal2 38226 17715 38226 17715 0 net9
rlabel via3 10925 2652 10925 2652 0 net90
rlabel metal2 2254 14433 2254 14433 0 net91
rlabel metal2 25254 2516 25254 2516 0 net92
rlabel metal2 37306 13872 37306 13872 0 net93
rlabel metal2 38042 26452 38042 26452 0 net94
rlabel metal1 34868 2414 34868 2414 0 net95
rlabel via3 13501 2652 13501 2652 0 net96
rlabel metal1 29762 36890 29762 36890 0 net97
rlabel metal1 19918 36346 19918 36346 0 net98
rlabel metal2 33626 3230 33626 3230 0 net99
rlabel metal2 14214 1775 14214 1775 0 pReset
rlabel metal2 4094 3519 4094 3519 0 prog_clk
rlabel metal3 38786 25908 38786 25908 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal2 21942 1860 21942 1860 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal1 29808 37230 29808 37230 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 28612 37230 28612 37230 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 1564 36142 1564 36142 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 6624 37230 6624 37230 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 27094 1554 27094 1554 0 right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal2 3818 9979 3818 9979 0 right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal3 1234 34748 1234 34748 0 right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal2 38318 18921 38318 18921 0 right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
