// This is the unpowered netlist.
module sb_4__0_ (ccff_head,
    ccff_tail,
    left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_,
    left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_,
    left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_,
    left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_,
    left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_,
    left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_,
    left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_,
    left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_,
    left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_,
    left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_,
    pReset,
    prog_clk,
    top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_,
    top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_,
    top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
    top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
    top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
    top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
    top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_,
    top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_,
    top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_,
    top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_,
    chanx_left_in,
    chanx_left_out,
    chany_top_in,
    chany_top_out);
 input ccff_head;
 output ccff_tail;
 input left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
 input left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
 input left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
 input left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
 input left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
 input left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
 input left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
 input left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
 input left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_;
 input left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_;
 input pReset;
 input prog_clk;
 input top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_;
 input top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_;
 input top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
 input top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
 input top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
 input top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
 input top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
 input top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
 input top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
 input top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
 input [0:18] chanx_left_in;
 output [0:18] chanx_left_out;
 input [0:18] chany_top_in;
 output [0:18] chany_top_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire clknet_0_prog_clk;
 wire \mem_left_track_1.DFFR_0_.D ;
 wire \mem_left_track_1.DFFR_0_.Q ;
 wire \mem_left_track_1.DFFR_1_.Q ;
 wire \mem_left_track_11.DFFR_0_.D ;
 wire \mem_left_track_11.DFFR_0_.Q ;
 wire \mem_left_track_11.DFFR_1_.Q ;
 wire \mem_left_track_13.DFFR_0_.Q ;
 wire \mem_left_track_13.DFFR_1_.Q ;
 wire \mem_left_track_15.DFFR_0_.Q ;
 wire \mem_left_track_15.DFFR_1_.Q ;
 wire \mem_left_track_17.DFFR_0_.Q ;
 wire \mem_left_track_17.DFFR_1_.Q ;
 wire \mem_left_track_19.DFFR_0_.Q ;
 wire \mem_left_track_19.DFFR_1_.Q ;
 wire \mem_left_track_21.DFFR_0_.Q ;
 wire \mem_left_track_21.DFFR_1_.Q ;
 wire \mem_left_track_23.DFFR_0_.Q ;
 wire \mem_left_track_23.DFFR_1_.Q ;
 wire \mem_left_track_25.DFFR_0_.Q ;
 wire \mem_left_track_25.DFFR_1_.Q ;
 wire \mem_left_track_27.DFFR_0_.Q ;
 wire \mem_left_track_27.DFFR_1_.Q ;
 wire \mem_left_track_29.DFFR_0_.Q ;
 wire \mem_left_track_29.DFFR_1_.Q ;
 wire \mem_left_track_3.DFFR_0_.Q ;
 wire \mem_left_track_3.DFFR_1_.Q ;
 wire \mem_left_track_31.DFFR_0_.Q ;
 wire \mem_left_track_31.DFFR_1_.Q ;
 wire \mem_left_track_33.DFFR_0_.Q ;
 wire \mem_left_track_33.DFFR_1_.Q ;
 wire \mem_left_track_35.DFFR_0_.Q ;
 wire \mem_left_track_35.DFFR_1_.Q ;
 wire \mem_left_track_37.DFFR_0_.Q ;
 wire \mem_left_track_5.DFFR_0_.Q ;
 wire \mem_left_track_5.DFFR_1_.Q ;
 wire \mem_left_track_7.DFFR_0_.Q ;
 wire \mem_left_track_7.DFFR_1_.Q ;
 wire \mem_left_track_9.DFFR_0_.Q ;
 wire \mem_top_track_0.DFFR_0_.Q ;
 wire \mem_top_track_0.DFFR_1_.Q ;
 wire \mem_top_track_10.DFFR_0_.D ;
 wire \mem_top_track_10.DFFR_0_.Q ;
 wire \mem_top_track_10.DFFR_1_.Q ;
 wire \mem_top_track_12.DFFR_0_.Q ;
 wire \mem_top_track_12.DFFR_1_.Q ;
 wire \mem_top_track_14.DFFR_0_.Q ;
 wire \mem_top_track_14.DFFR_1_.Q ;
 wire \mem_top_track_16.DFFR_0_.Q ;
 wire \mem_top_track_16.DFFR_1_.Q ;
 wire \mem_top_track_18.DFFR_0_.Q ;
 wire \mem_top_track_18.DFFR_1_.Q ;
 wire \mem_top_track_2.DFFR_0_.Q ;
 wire \mem_top_track_2.DFFR_1_.Q ;
 wire \mem_top_track_20.DFFR_0_.Q ;
 wire \mem_top_track_20.DFFR_1_.Q ;
 wire \mem_top_track_22.DFFR_0_.Q ;
 wire \mem_top_track_22.DFFR_1_.Q ;
 wire \mem_top_track_24.DFFR_0_.Q ;
 wire \mem_top_track_24.DFFR_1_.Q ;
 wire \mem_top_track_26.DFFR_0_.Q ;
 wire \mem_top_track_26.DFFR_1_.Q ;
 wire \mem_top_track_28.DFFR_0_.Q ;
 wire \mem_top_track_28.DFFR_1_.Q ;
 wire \mem_top_track_30.DFFR_0_.Q ;
 wire \mem_top_track_30.DFFR_1_.Q ;
 wire \mem_top_track_32.DFFR_0_.Q ;
 wire \mem_top_track_32.DFFR_1_.Q ;
 wire \mem_top_track_34.DFFR_0_.Q ;
 wire \mem_top_track_34.DFFR_1_.Q ;
 wire \mem_top_track_36.DFFR_0_.Q ;
 wire \mem_top_track_4.DFFR_0_.Q ;
 wire \mem_top_track_4.DFFR_1_.Q ;
 wire \mem_top_track_6.DFFR_0_.Q ;
 wire \mem_top_track_6.DFFR_1_.Q ;
 wire \mem_top_track_8.DFFR_0_.Q ;
 wire \mux_left_track_1.INVTX1_0_.out ;
 wire \mux_left_track_1.INVTX1_1_.out ;
 wire \mux_left_track_1.INVTX1_2_.out ;
 wire \mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_left_track_1.out ;
 wire \mux_left_track_11.INVTX1_0_.out ;
 wire \mux_left_track_11.INVTX1_1_.out ;
 wire \mux_left_track_11.INVTX1_2_.out ;
 wire \mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_left_track_11.out ;
 wire \mux_left_track_13.INVTX1_0_.out ;
 wire \mux_left_track_13.INVTX1_2_.out ;
 wire \mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_left_track_13.out ;
 wire \mux_left_track_15.INVTX1_0_.out ;
 wire \mux_left_track_15.INVTX1_2_.out ;
 wire \mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_left_track_15.out ;
 wire \mux_left_track_17.INVTX1_0_.out ;
 wire \mux_left_track_17.INVTX1_2_.out ;
 wire \mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_left_track_17.out ;
 wire \mux_left_track_19.INVTX1_0_.out ;
 wire \mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_left_track_19.out ;
 wire \mux_left_track_21.INVTX1_0_.out ;
 wire \mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_left_track_21.out ;
 wire \mux_left_track_23.INVTX1_0_.out ;
 wire \mux_left_track_23.INVTX1_1_.out ;
 wire \mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_left_track_23.out ;
 wire \mux_left_track_25.INVTX1_0_.out ;
 wire \mux_left_track_25.INVTX1_1_.out ;
 wire \mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_left_track_25.out ;
 wire \mux_left_track_27.INVTX1_0_.out ;
 wire \mux_left_track_27.INVTX1_1_.out ;
 wire \mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_left_track_27.out ;
 wire \mux_left_track_29.INVTX1_0_.out ;
 wire \mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_left_track_29.out ;
 wire \mux_left_track_3.INVTX1_0_.out ;
 wire \mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_left_track_3.out ;
 wire \mux_left_track_31.INVTX1_0_.out ;
 wire \mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_left_track_31.out ;
 wire \mux_left_track_33.INVTX1_0_.out ;
 wire \mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_left_track_33.out ;
 wire \mux_left_track_35.INVTX1_0_.out ;
 wire \mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_left_track_35.out ;
 wire \mux_left_track_37.INVTX1_0_.out ;
 wire \mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_left_track_37.out ;
 wire \mux_left_track_5.INVTX1_0_.out ;
 wire \mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_left_track_5.out ;
 wire \mux_left_track_7.INVTX1_0_.out ;
 wire \mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_left_track_7.out ;
 wire \mux_left_track_9.INVTX1_0_.out ;
 wire \mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_left_track_9.out ;
 wire \mux_top_track_0.INVTX1_0_.out ;
 wire \mux_top_track_0.INVTX1_1_.out ;
 wire \mux_top_track_0.INVTX1_2_.out ;
 wire \mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_top_track_0.out ;
 wire \mux_top_track_10.INVTX1_0_.out ;
 wire \mux_top_track_10.INVTX1_1_.out ;
 wire \mux_top_track_10.INVTX1_2_.out ;
 wire \mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_top_track_10.out ;
 wire \mux_top_track_12.INVTX1_1_.out ;
 wire \mux_top_track_12.INVTX1_2_.out ;
 wire \mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_top_track_12.out ;
 wire \mux_top_track_14.INVTX1_1_.out ;
 wire \mux_top_track_14.INVTX1_2_.out ;
 wire \mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_top_track_14.out ;
 wire \mux_top_track_16.INVTX1_1_.out ;
 wire \mux_top_track_16.INVTX1_2_.out ;
 wire \mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_top_track_16.out ;
 wire \mux_top_track_18.INVTX1_2_.out ;
 wire \mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_top_track_18.out ;
 wire \mux_top_track_2.INVTX1_1_.out ;
 wire \mux_top_track_2.INVTX1_2_.out ;
 wire \mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_top_track_2.out ;
 wire \mux_top_track_20.INVTX1_1_.out ;
 wire \mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_top_track_20.out ;
 wire \mux_top_track_22.INVTX1_1_.out ;
 wire \mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_top_track_22.out ;
 wire \mux_top_track_24.INVTX1_0_.out ;
 wire \mux_top_track_24.INVTX1_1_.out ;
 wire \mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_top_track_24.out ;
 wire \mux_top_track_26.INVTX1_0_.out ;
 wire \mux_top_track_26.INVTX1_1_.out ;
 wire \mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_top_track_26.out ;
 wire \mux_top_track_28.INVTX1_1_.out ;
 wire \mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_top_track_28.out ;
 wire \mux_top_track_30.INVTX1_1_.out ;
 wire \mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_top_track_30.out ;
 wire \mux_top_track_32.INVTX1_1_.out ;
 wire \mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_top_track_32.out ;
 wire \mux_top_track_34.INVTX1_1_.out ;
 wire \mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_top_track_34.out ;
 wire \mux_top_track_36.INVTX1_2_.out ;
 wire \mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_top_track_36.out ;
 wire \mux_top_track_4.INVTX1_2_.out ;
 wire \mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_top_track_4.out ;
 wire \mux_top_track_6.INVTX1_2_.out ;
 wire \mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_top_track_6.out ;
 wire \mux_top_track_8.INVTX1_2_.out ;
 wire \mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_top_track_8.out ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire clknet_3_0__leaf_prog_clk;
 wire clknet_3_1__leaf_prog_clk;
 wire clknet_3_2__leaf_prog_clk;
 wire clknet_3_3__leaf_prog_clk;
 wire clknet_3_4__leaf_prog_clk;
 wire clknet_3_5__leaf_prog_clk;
 wire clknet_3_6__leaf_prog_clk;
 wire clknet_3_7__leaf_prog_clk;

 sky130_fd_sc_hd__inv_2 _0416_ (.A(\mem_left_track_35.DFFR_1_.Q ),
    .Y(_0376_));
 sky130_fd_sc_hd__inv_2 _0417_ (.A(\mem_left_track_35.DFFR_0_.Q ),
    .Y(_0377_));
 sky130_fd_sc_hd__clkbuf_1 _0418_ (.A(\mem_left_track_35.DFFR_0_.Q ),
    .X(_0076_));
 sky130_fd_sc_hd__clkbuf_1 _0419_ (.A(_0076_),
    .X(_0375_));
 sky130_fd_sc_hd__clkbuf_1 _0420_ (.A(\mem_left_track_35.DFFR_1_.Q ),
    .X(_0077_));
 sky130_fd_sc_hd__clkbuf_1 _0421_ (.A(_0077_),
    .X(_0374_));
 sky130_fd_sc_hd__inv_2 _0422_ (.A(\mem_left_track_33.DFFR_1_.Q ),
    .Y(_0372_));
 sky130_fd_sc_hd__inv_2 _0423_ (.A(\mem_left_track_33.DFFR_0_.Q ),
    .Y(_0373_));
 sky130_fd_sc_hd__clkbuf_1 _0424_ (.A(\mem_left_track_33.DFFR_0_.Q ),
    .X(_0078_));
 sky130_fd_sc_hd__clkbuf_1 _0425_ (.A(_0078_),
    .X(_0371_));
 sky130_fd_sc_hd__clkbuf_1 _0426_ (.A(\mem_left_track_33.DFFR_1_.Q ),
    .X(_0079_));
 sky130_fd_sc_hd__clkbuf_1 _0427_ (.A(_0079_),
    .X(_0370_));
 sky130_fd_sc_hd__inv_2 _0428_ (.A(\mem_left_track_31.DFFR_1_.Q ),
    .Y(_0368_));
 sky130_fd_sc_hd__inv_2 _0429_ (.A(\mem_left_track_31.DFFR_0_.Q ),
    .Y(_0369_));
 sky130_fd_sc_hd__clkbuf_1 _0430_ (.A(\mem_left_track_31.DFFR_0_.Q ),
    .X(_0080_));
 sky130_fd_sc_hd__clkbuf_1 _0431_ (.A(_0080_),
    .X(_0367_));
 sky130_fd_sc_hd__clkbuf_1 _0432_ (.A(\mem_left_track_31.DFFR_1_.Q ),
    .X(_0081_));
 sky130_fd_sc_hd__clkbuf_1 _0433_ (.A(_0081_),
    .X(_0366_));
 sky130_fd_sc_hd__inv_2 _0434_ (.A(\mem_left_track_29.DFFR_1_.Q ),
    .Y(_0364_));
 sky130_fd_sc_hd__inv_2 _0435_ (.A(\mem_left_track_29.DFFR_0_.Q ),
    .Y(_0365_));
 sky130_fd_sc_hd__clkbuf_1 _0436_ (.A(\mem_left_track_29.DFFR_0_.Q ),
    .X(_0082_));
 sky130_fd_sc_hd__clkbuf_1 _0437_ (.A(_0082_),
    .X(_0363_));
 sky130_fd_sc_hd__clkbuf_1 _0438_ (.A(\mem_left_track_29.DFFR_1_.Q ),
    .X(_0083_));
 sky130_fd_sc_hd__clkbuf_1 _0439_ (.A(_0083_),
    .X(_0362_));
 sky130_fd_sc_hd__inv_2 _0440_ (.A(\mem_left_track_27.DFFR_1_.Q ),
    .Y(_0360_));
 sky130_fd_sc_hd__inv_2 _0441_ (.A(\mem_left_track_27.DFFR_0_.Q ),
    .Y(_0361_));
 sky130_fd_sc_hd__clkbuf_1 _0442_ (.A(\mem_left_track_27.DFFR_0_.Q ),
    .X(_0084_));
 sky130_fd_sc_hd__clkbuf_1 _0443_ (.A(_0084_),
    .X(_0359_));
 sky130_fd_sc_hd__clkbuf_1 _0444_ (.A(\mem_left_track_27.DFFR_1_.Q ),
    .X(_0085_));
 sky130_fd_sc_hd__clkbuf_1 _0445_ (.A(_0085_),
    .X(_0358_));
 sky130_fd_sc_hd__inv_2 _0446_ (.A(\mem_left_track_25.DFFR_1_.Q ),
    .Y(_0356_));
 sky130_fd_sc_hd__inv_2 _0447_ (.A(\mem_left_track_25.DFFR_0_.Q ),
    .Y(_0357_));
 sky130_fd_sc_hd__clkbuf_1 _0448_ (.A(\mem_left_track_25.DFFR_0_.Q ),
    .X(_0086_));
 sky130_fd_sc_hd__clkbuf_1 _0449_ (.A(_0086_),
    .X(_0355_));
 sky130_fd_sc_hd__clkbuf_1 _0450_ (.A(\mem_left_track_25.DFFR_1_.Q ),
    .X(_0087_));
 sky130_fd_sc_hd__clkbuf_1 _0451_ (.A(_0087_),
    .X(_0354_));
 sky130_fd_sc_hd__inv_2 _0452_ (.A(\mem_left_track_23.DFFR_1_.Q ),
    .Y(_0352_));
 sky130_fd_sc_hd__inv_2 _0453_ (.A(\mem_left_track_23.DFFR_0_.Q ),
    .Y(_0353_));
 sky130_fd_sc_hd__clkbuf_1 _0454_ (.A(\mem_left_track_23.DFFR_0_.Q ),
    .X(_0088_));
 sky130_fd_sc_hd__clkbuf_1 _0455_ (.A(_0088_),
    .X(_0351_));
 sky130_fd_sc_hd__clkbuf_1 _0456_ (.A(\mem_top_track_0.DFFR_1_.Q ),
    .X(_0089_));
 sky130_fd_sc_hd__clkbuf_1 _0457_ (.A(_0089_),
    .X(_0182_));
 sky130_fd_sc_hd__clkbuf_1 _0458_ (.A(\mem_left_track_23.DFFR_1_.Q ),
    .X(_0090_));
 sky130_fd_sc_hd__clkbuf_1 _0459_ (.A(_0090_),
    .X(_0350_));
 sky130_fd_sc_hd__inv_2 _0460_ (.A(\mem_left_track_21.DFFR_1_.Q ),
    .Y(_0348_));
 sky130_fd_sc_hd__inv_2 _0461_ (.A(\mem_left_track_21.DFFR_0_.Q ),
    .Y(_0349_));
 sky130_fd_sc_hd__clkbuf_1 _0462_ (.A(\mem_left_track_21.DFFR_0_.Q ),
    .X(_0091_));
 sky130_fd_sc_hd__clkbuf_1 _0463_ (.A(_0091_),
    .X(_0347_));
 sky130_fd_sc_hd__clkbuf_1 _0464_ (.A(\mem_left_track_21.DFFR_1_.Q ),
    .X(_0092_));
 sky130_fd_sc_hd__clkbuf_1 _0465_ (.A(_0092_),
    .X(_0346_));
 sky130_fd_sc_hd__inv_2 _0466_ (.A(\mem_top_track_34.DFFR_1_.Q ),
    .Y(_0344_));
 sky130_fd_sc_hd__inv_2 _0467_ (.A(\mem_top_track_34.DFFR_0_.Q ),
    .Y(_0345_));
 sky130_fd_sc_hd__clkbuf_1 _0468_ (.A(\mem_top_track_34.DFFR_0_.Q ),
    .X(_0093_));
 sky130_fd_sc_hd__clkbuf_1 _0469_ (.A(_0093_),
    .X(_0343_));
 sky130_fd_sc_hd__clkbuf_1 _0470_ (.A(\mem_top_track_34.DFFR_1_.Q ),
    .X(_0094_));
 sky130_fd_sc_hd__clkbuf_1 _0471_ (.A(_0094_),
    .X(_0342_));
 sky130_fd_sc_hd__inv_2 _0472_ (.A(\mem_top_track_32.DFFR_1_.Q ),
    .Y(_0340_));
 sky130_fd_sc_hd__inv_2 _0473_ (.A(\mem_top_track_32.DFFR_0_.Q ),
    .Y(_0341_));
 sky130_fd_sc_hd__clkbuf_1 _0474_ (.A(\mem_top_track_32.DFFR_0_.Q ),
    .X(_0095_));
 sky130_fd_sc_hd__clkbuf_1 _0475_ (.A(_0095_),
    .X(_0339_));
 sky130_fd_sc_hd__clkbuf_1 _0476_ (.A(\mem_top_track_32.DFFR_1_.Q ),
    .X(_0096_));
 sky130_fd_sc_hd__clkbuf_1 _0477_ (.A(_0096_),
    .X(_0338_));
 sky130_fd_sc_hd__inv_2 _0478_ (.A(\mem_top_track_30.DFFR_1_.Q ),
    .Y(_0336_));
 sky130_fd_sc_hd__inv_2 _0479_ (.A(\mem_top_track_30.DFFR_0_.Q ),
    .Y(_0337_));
 sky130_fd_sc_hd__clkbuf_1 _0480_ (.A(\mem_top_track_30.DFFR_0_.Q ),
    .X(_0097_));
 sky130_fd_sc_hd__clkbuf_1 _0481_ (.A(_0097_),
    .X(_0335_));
 sky130_fd_sc_hd__clkbuf_1 _0482_ (.A(\mem_top_track_30.DFFR_1_.Q ),
    .X(_0098_));
 sky130_fd_sc_hd__clkbuf_1 _0483_ (.A(_0098_),
    .X(_0334_));
 sky130_fd_sc_hd__inv_2 _0484_ (.A(\mem_top_track_28.DFFR_1_.Q ),
    .Y(_0332_));
 sky130_fd_sc_hd__inv_2 _0485_ (.A(\mem_top_track_28.DFFR_0_.Q ),
    .Y(_0333_));
 sky130_fd_sc_hd__clkbuf_1 _0486_ (.A(\mem_top_track_28.DFFR_0_.Q ),
    .X(_0099_));
 sky130_fd_sc_hd__clkbuf_1 _0487_ (.A(_0099_),
    .X(_0331_));
 sky130_fd_sc_hd__clkbuf_1 _0488_ (.A(\mem_top_track_28.DFFR_1_.Q ),
    .X(_0100_));
 sky130_fd_sc_hd__clkbuf_1 _0489_ (.A(_0100_),
    .X(_0330_));
 sky130_fd_sc_hd__inv_2 _0490_ (.A(\mem_top_track_26.DFFR_1_.Q ),
    .Y(_0328_));
 sky130_fd_sc_hd__inv_2 _0491_ (.A(\mem_top_track_26.DFFR_0_.Q ),
    .Y(_0329_));
 sky130_fd_sc_hd__clkbuf_1 _0492_ (.A(\mem_top_track_26.DFFR_0_.Q ),
    .X(_0101_));
 sky130_fd_sc_hd__clkbuf_1 _0493_ (.A(_0101_),
    .X(_0327_));
 sky130_fd_sc_hd__clkbuf_1 _0494_ (.A(\mem_top_track_26.DFFR_1_.Q ),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_1 _0495_ (.A(_0102_),
    .X(_0326_));
 sky130_fd_sc_hd__inv_2 _0496_ (.A(\mem_top_track_24.DFFR_1_.Q ),
    .Y(_0324_));
 sky130_fd_sc_hd__inv_2 _0497_ (.A(\mem_top_track_24.DFFR_0_.Q ),
    .Y(_0325_));
 sky130_fd_sc_hd__clkbuf_1 _0498_ (.A(\mem_top_track_24.DFFR_0_.Q ),
    .X(_0103_));
 sky130_fd_sc_hd__clkbuf_1 _0499_ (.A(_0103_),
    .X(_0323_));
 sky130_fd_sc_hd__clkbuf_1 _0500_ (.A(\mem_top_track_24.DFFR_1_.Q ),
    .X(_0104_));
 sky130_fd_sc_hd__clkbuf_1 _0501_ (.A(_0104_),
    .X(_0322_));
 sky130_fd_sc_hd__inv_2 _0502_ (.A(\mem_top_track_22.DFFR_1_.Q ),
    .Y(_0320_));
 sky130_fd_sc_hd__inv_2 _0503_ (.A(\mem_top_track_22.DFFR_0_.Q ),
    .Y(_0321_));
 sky130_fd_sc_hd__clkbuf_1 _0504_ (.A(\mem_top_track_22.DFFR_0_.Q ),
    .X(_0105_));
 sky130_fd_sc_hd__clkbuf_1 _0505_ (.A(_0105_),
    .X(_0319_));
 sky130_fd_sc_hd__clkbuf_1 _0506_ (.A(\mem_top_track_22.DFFR_1_.Q ),
    .X(_0106_));
 sky130_fd_sc_hd__clkbuf_1 _0507_ (.A(_0106_),
    .X(_0318_));
 sky130_fd_sc_hd__inv_2 _0508_ (.A(\mem_top_track_20.DFFR_1_.Q ),
    .Y(_0316_));
 sky130_fd_sc_hd__inv_2 _0509_ (.A(\mem_top_track_20.DFFR_0_.Q ),
    .Y(_0317_));
 sky130_fd_sc_hd__clkbuf_1 _0510_ (.A(\mem_top_track_20.DFFR_0_.Q ),
    .X(_0107_));
 sky130_fd_sc_hd__clkbuf_1 _0511_ (.A(_0107_),
    .X(_0315_));
 sky130_fd_sc_hd__clkbuf_1 _0512_ (.A(\mem_top_track_20.DFFR_1_.Q ),
    .X(_0108_));
 sky130_fd_sc_hd__clkbuf_1 _0513_ (.A(_0108_),
    .X(_0314_));
 sky130_fd_sc_hd__inv_2 _0514_ (.A(net61),
    .Y(_0311_));
 sky130_fd_sc_hd__inv_2 _0515_ (.A(\mem_left_track_37.DFFR_0_.Q ),
    .Y(_0313_));
 sky130_fd_sc_hd__clkbuf_1 _0516_ (.A(\mem_left_track_37.DFFR_0_.Q ),
    .X(_0109_));
 sky130_fd_sc_hd__clkbuf_1 _0517_ (.A(_0109_),
    .X(_0310_));
 sky130_fd_sc_hd__clkbuf_1 _0518_ (.A(net61),
    .X(_0110_));
 sky130_fd_sc_hd__clkbuf_1 _0519_ (.A(_0110_),
    .X(_0308_));
 sky130_fd_sc_hd__inv_2 _0520_ (.A(\mem_left_track_37.DFFR_0_.Q ),
    .Y(_0312_));
 sky130_fd_sc_hd__clkbuf_1 _0521_ (.A(\mem_left_track_37.DFFR_0_.Q ),
    .X(_0111_));
 sky130_fd_sc_hd__clkbuf_1 _0522_ (.A(_0111_),
    .X(_0309_));
 sky130_fd_sc_hd__inv_2 _0523_ (.A(\mem_left_track_19.DFFR_1_.Q ),
    .Y(_0305_));
 sky130_fd_sc_hd__inv_2 _0524_ (.A(\mem_left_track_19.DFFR_0_.Q ),
    .Y(_0307_));
 sky130_fd_sc_hd__clkbuf_1 _0525_ (.A(\mem_left_track_19.DFFR_0_.Q ),
    .X(_0112_));
 sky130_fd_sc_hd__clkbuf_1 _0526_ (.A(_0112_),
    .X(_0304_));
 sky130_fd_sc_hd__clkbuf_1 _0527_ (.A(\mem_left_track_19.DFFR_1_.Q ),
    .X(_0113_));
 sky130_fd_sc_hd__clkbuf_1 _0528_ (.A(_0113_),
    .X(_0302_));
 sky130_fd_sc_hd__inv_2 _0529_ (.A(\mem_left_track_19.DFFR_0_.Q ),
    .Y(_0306_));
 sky130_fd_sc_hd__clkbuf_1 _0530_ (.A(\mem_left_track_19.DFFR_0_.Q ),
    .X(_0114_));
 sky130_fd_sc_hd__clkbuf_1 _0531_ (.A(_0114_),
    .X(_0303_));
 sky130_fd_sc_hd__inv_2 _0532_ (.A(\mem_left_track_17.DFFR_1_.Q ),
    .Y(_0299_));
 sky130_fd_sc_hd__inv_2 _0533_ (.A(\mem_left_track_17.DFFR_0_.Q ),
    .Y(_0301_));
 sky130_fd_sc_hd__clkbuf_1 _0534_ (.A(\mem_left_track_17.DFFR_0_.Q ),
    .X(_0115_));
 sky130_fd_sc_hd__clkbuf_1 _0535_ (.A(_0115_),
    .X(_0298_));
 sky130_fd_sc_hd__clkbuf_1 _0536_ (.A(\mem_left_track_17.DFFR_1_.Q ),
    .X(_0116_));
 sky130_fd_sc_hd__clkbuf_1 _0537_ (.A(_0116_),
    .X(_0296_));
 sky130_fd_sc_hd__inv_2 _0538_ (.A(\mem_left_track_17.DFFR_0_.Q ),
    .Y(_0300_));
 sky130_fd_sc_hd__clkbuf_1 _0539_ (.A(\mem_left_track_17.DFFR_0_.Q ),
    .X(_0117_));
 sky130_fd_sc_hd__clkbuf_1 _0540_ (.A(_0117_),
    .X(_0297_));
 sky130_fd_sc_hd__inv_2 _0541_ (.A(\mem_left_track_15.DFFR_1_.Q ),
    .Y(_0293_));
 sky130_fd_sc_hd__inv_2 _0542_ (.A(\mem_left_track_15.DFFR_0_.Q ),
    .Y(_0295_));
 sky130_fd_sc_hd__clkbuf_1 _0543_ (.A(\mem_left_track_15.DFFR_0_.Q ),
    .X(_0118_));
 sky130_fd_sc_hd__clkbuf_1 _0544_ (.A(_0118_),
    .X(_0292_));
 sky130_fd_sc_hd__clkbuf_1 _0545_ (.A(\mem_left_track_15.DFFR_1_.Q ),
    .X(_0119_));
 sky130_fd_sc_hd__clkbuf_1 _0546_ (.A(_0119_),
    .X(_0290_));
 sky130_fd_sc_hd__inv_2 _0547_ (.A(\mem_left_track_15.DFFR_0_.Q ),
    .Y(_0294_));
 sky130_fd_sc_hd__clkbuf_1 _0548_ (.A(\mem_left_track_15.DFFR_0_.Q ),
    .X(_0120_));
 sky130_fd_sc_hd__clkbuf_1 _0549_ (.A(_0120_),
    .X(_0291_));
 sky130_fd_sc_hd__inv_2 _0550_ (.A(\mem_left_track_13.DFFR_1_.Q ),
    .Y(_0287_));
 sky130_fd_sc_hd__inv_2 _0551_ (.A(\mem_left_track_13.DFFR_0_.Q ),
    .Y(_0289_));
 sky130_fd_sc_hd__clkbuf_1 _0552_ (.A(\mem_left_track_13.DFFR_0_.Q ),
    .X(_0121_));
 sky130_fd_sc_hd__clkbuf_1 _0553_ (.A(_0121_),
    .X(_0286_));
 sky130_fd_sc_hd__clkbuf_1 _0554_ (.A(\mem_left_track_13.DFFR_1_.Q ),
    .X(_0122_));
 sky130_fd_sc_hd__clkbuf_1 _0555_ (.A(_0122_),
    .X(_0284_));
 sky130_fd_sc_hd__inv_2 _0556_ (.A(\mem_left_track_13.DFFR_0_.Q ),
    .Y(_0288_));
 sky130_fd_sc_hd__clkbuf_1 _0557_ (.A(\mem_left_track_13.DFFR_0_.Q ),
    .X(_0123_));
 sky130_fd_sc_hd__clkbuf_1 _0558_ (.A(_0123_),
    .X(_0285_));
 sky130_fd_sc_hd__inv_2 _0559_ (.A(\mem_left_track_11.DFFR_1_.Q ),
    .Y(_0281_));
 sky130_fd_sc_hd__inv_2 _0560_ (.A(\mem_left_track_11.DFFR_0_.Q ),
    .Y(_0283_));
 sky130_fd_sc_hd__clkbuf_1 _0561_ (.A(\mem_left_track_11.DFFR_0_.Q ),
    .X(_0124_));
 sky130_fd_sc_hd__clkbuf_1 _0562_ (.A(_0124_),
    .X(_0280_));
 sky130_fd_sc_hd__clkbuf_1 _0563_ (.A(\mem_left_track_11.DFFR_1_.Q ),
    .X(_0125_));
 sky130_fd_sc_hd__clkbuf_1 _0564_ (.A(_0125_),
    .X(_0278_));
 sky130_fd_sc_hd__inv_2 _0565_ (.A(\mem_left_track_11.DFFR_0_.Q ),
    .Y(_0282_));
 sky130_fd_sc_hd__clkbuf_1 _0566_ (.A(\mem_left_track_11.DFFR_0_.Q ),
    .X(_0126_));
 sky130_fd_sc_hd__clkbuf_1 _0567_ (.A(_0126_),
    .X(_0279_));
 sky130_fd_sc_hd__inv_2 _0568_ (.A(\mem_left_track_11.DFFR_0_.D ),
    .Y(_0275_));
 sky130_fd_sc_hd__inv_2 _0569_ (.A(\mem_left_track_9.DFFR_0_.Q ),
    .Y(_0277_));
 sky130_fd_sc_hd__clkbuf_1 _0570_ (.A(\mem_left_track_9.DFFR_0_.Q ),
    .X(_0127_));
 sky130_fd_sc_hd__clkbuf_1 _0571_ (.A(_0127_),
    .X(_0274_));
 sky130_fd_sc_hd__clkbuf_1 _0572_ (.A(\mem_left_track_11.DFFR_0_.D ),
    .X(_0128_));
 sky130_fd_sc_hd__clkbuf_1 _0573_ (.A(_0128_),
    .X(_0272_));
 sky130_fd_sc_hd__inv_2 _0574_ (.A(\mem_left_track_9.DFFR_0_.Q ),
    .Y(_0276_));
 sky130_fd_sc_hd__clkbuf_1 _0575_ (.A(\mem_left_track_9.DFFR_0_.Q ),
    .X(_0129_));
 sky130_fd_sc_hd__clkbuf_1 _0576_ (.A(_0129_),
    .X(_0273_));
 sky130_fd_sc_hd__inv_2 _0577_ (.A(\mem_left_track_7.DFFR_1_.Q ),
    .Y(_0269_));
 sky130_fd_sc_hd__inv_2 _0578_ (.A(\mem_left_track_7.DFFR_0_.Q ),
    .Y(_0271_));
 sky130_fd_sc_hd__clkbuf_1 _0579_ (.A(\mem_left_track_7.DFFR_0_.Q ),
    .X(_0130_));
 sky130_fd_sc_hd__clkbuf_1 _0580_ (.A(_0130_),
    .X(_0268_));
 sky130_fd_sc_hd__clkbuf_1 _0581_ (.A(\mem_left_track_7.DFFR_1_.Q ),
    .X(_0131_));
 sky130_fd_sc_hd__clkbuf_1 _0582_ (.A(_0131_),
    .X(_0266_));
 sky130_fd_sc_hd__inv_2 _0583_ (.A(\mem_left_track_7.DFFR_0_.Q ),
    .Y(_0270_));
 sky130_fd_sc_hd__clkbuf_1 _0584_ (.A(\mem_left_track_7.DFFR_0_.Q ),
    .X(_0132_));
 sky130_fd_sc_hd__clkbuf_1 _0585_ (.A(_0132_),
    .X(_0267_));
 sky130_fd_sc_hd__inv_2 _0586_ (.A(\mem_left_track_5.DFFR_1_.Q ),
    .Y(_0263_));
 sky130_fd_sc_hd__inv_2 _0587_ (.A(\mem_left_track_5.DFFR_0_.Q ),
    .Y(_0265_));
 sky130_fd_sc_hd__clkbuf_1 _0588_ (.A(\mem_left_track_5.DFFR_0_.Q ),
    .X(_0133_));
 sky130_fd_sc_hd__clkbuf_1 _0589_ (.A(_0133_),
    .X(_0262_));
 sky130_fd_sc_hd__clkbuf_1 _0590_ (.A(\mem_left_track_5.DFFR_1_.Q ),
    .X(_0134_));
 sky130_fd_sc_hd__clkbuf_1 _0591_ (.A(_0134_),
    .X(_0260_));
 sky130_fd_sc_hd__inv_2 _0592_ (.A(\mem_left_track_5.DFFR_0_.Q ),
    .Y(_0264_));
 sky130_fd_sc_hd__clkbuf_1 _0593_ (.A(\mem_left_track_5.DFFR_0_.Q ),
    .X(_0135_));
 sky130_fd_sc_hd__clkbuf_1 _0594_ (.A(_0135_),
    .X(_0261_));
 sky130_fd_sc_hd__inv_2 _0595_ (.A(\mem_left_track_3.DFFR_1_.Q ),
    .Y(_0257_));
 sky130_fd_sc_hd__inv_2 _0596_ (.A(\mem_left_track_3.DFFR_0_.Q ),
    .Y(_0259_));
 sky130_fd_sc_hd__clkbuf_1 _0597_ (.A(\mem_left_track_3.DFFR_0_.Q ),
    .X(_0136_));
 sky130_fd_sc_hd__clkbuf_1 _0598_ (.A(_0136_),
    .X(_0256_));
 sky130_fd_sc_hd__clkbuf_1 _0599_ (.A(\mem_left_track_3.DFFR_1_.Q ),
    .X(_0137_));
 sky130_fd_sc_hd__clkbuf_1 _0600_ (.A(_0137_),
    .X(_0254_));
 sky130_fd_sc_hd__inv_2 _0601_ (.A(\mem_left_track_3.DFFR_0_.Q ),
    .Y(_0258_));
 sky130_fd_sc_hd__clkbuf_1 _0602_ (.A(\mem_left_track_3.DFFR_0_.Q ),
    .X(_0138_));
 sky130_fd_sc_hd__clkbuf_1 _0603_ (.A(_0138_),
    .X(_0255_));
 sky130_fd_sc_hd__inv_2 _0604_ (.A(\mem_left_track_1.DFFR_1_.Q ),
    .Y(_0251_));
 sky130_fd_sc_hd__inv_2 _0605_ (.A(\mem_left_track_1.DFFR_0_.Q ),
    .Y(_0253_));
 sky130_fd_sc_hd__clkbuf_1 _0606_ (.A(\mem_left_track_1.DFFR_0_.Q ),
    .X(_0139_));
 sky130_fd_sc_hd__clkbuf_1 _0607_ (.A(_0139_),
    .X(_0250_));
 sky130_fd_sc_hd__clkbuf_1 _0608_ (.A(\mem_left_track_1.DFFR_1_.Q ),
    .X(_0140_));
 sky130_fd_sc_hd__clkbuf_1 _0609_ (.A(_0140_),
    .X(_0248_));
 sky130_fd_sc_hd__inv_2 _0610_ (.A(\mem_left_track_1.DFFR_0_.Q ),
    .Y(_0252_));
 sky130_fd_sc_hd__clkbuf_1 _0611_ (.A(\mem_left_track_1.DFFR_0_.Q ),
    .X(_0141_));
 sky130_fd_sc_hd__clkbuf_1 _0612_ (.A(_0141_),
    .X(_0249_));
 sky130_fd_sc_hd__inv_2 _0613_ (.A(\mem_left_track_1.DFFR_0_.D ),
    .Y(_0245_));
 sky130_fd_sc_hd__inv_2 _0614_ (.A(\mem_top_track_36.DFFR_0_.Q ),
    .Y(_0247_));
 sky130_fd_sc_hd__clkbuf_1 _0615_ (.A(\mem_top_track_36.DFFR_0_.Q ),
    .X(_0142_));
 sky130_fd_sc_hd__clkbuf_1 _0616_ (.A(_0142_),
    .X(_0244_));
 sky130_fd_sc_hd__clkbuf_1 _0617_ (.A(\mem_left_track_1.DFFR_0_.D ),
    .X(_0143_));
 sky130_fd_sc_hd__clkbuf_1 _0618_ (.A(_0143_),
    .X(_0242_));
 sky130_fd_sc_hd__inv_2 _0619_ (.A(\mem_top_track_36.DFFR_0_.Q ),
    .Y(_0246_));
 sky130_fd_sc_hd__clkbuf_1 _0620_ (.A(\mem_top_track_36.DFFR_0_.Q ),
    .X(_0144_));
 sky130_fd_sc_hd__clkbuf_1 _0621_ (.A(_0144_),
    .X(_0243_));
 sky130_fd_sc_hd__inv_2 _0622_ (.A(\mem_top_track_18.DFFR_1_.Q ),
    .Y(_0239_));
 sky130_fd_sc_hd__inv_2 _0623_ (.A(\mem_top_track_18.DFFR_0_.Q ),
    .Y(_0241_));
 sky130_fd_sc_hd__clkbuf_1 _0624_ (.A(\mem_top_track_18.DFFR_0_.Q ),
    .X(_0145_));
 sky130_fd_sc_hd__clkbuf_1 _0625_ (.A(_0145_),
    .X(_0238_));
 sky130_fd_sc_hd__clkbuf_1 _0626_ (.A(\mem_top_track_18.DFFR_1_.Q ),
    .X(_0146_));
 sky130_fd_sc_hd__clkbuf_1 _0627_ (.A(_0146_),
    .X(_0236_));
 sky130_fd_sc_hd__inv_2 _0628_ (.A(\mem_top_track_18.DFFR_0_.Q ),
    .Y(_0240_));
 sky130_fd_sc_hd__clkbuf_1 _0629_ (.A(\mem_top_track_18.DFFR_0_.Q ),
    .X(_0147_));
 sky130_fd_sc_hd__clkbuf_1 _0630_ (.A(_0147_),
    .X(_0237_));
 sky130_fd_sc_hd__inv_2 _0631_ (.A(\mem_top_track_16.DFFR_1_.Q ),
    .Y(_0233_));
 sky130_fd_sc_hd__inv_2 _0632_ (.A(\mem_top_track_16.DFFR_0_.Q ),
    .Y(_0235_));
 sky130_fd_sc_hd__clkbuf_1 _0633_ (.A(\mem_top_track_16.DFFR_0_.Q ),
    .X(_0148_));
 sky130_fd_sc_hd__clkbuf_1 _0634_ (.A(_0148_),
    .X(_0232_));
 sky130_fd_sc_hd__clkbuf_1 _0635_ (.A(\mem_top_track_16.DFFR_1_.Q ),
    .X(_0149_));
 sky130_fd_sc_hd__clkbuf_1 _0636_ (.A(_0149_),
    .X(_0230_));
 sky130_fd_sc_hd__inv_2 _0637_ (.A(\mem_top_track_16.DFFR_0_.Q ),
    .Y(_0234_));
 sky130_fd_sc_hd__clkbuf_1 _0638_ (.A(\mem_top_track_16.DFFR_0_.Q ),
    .X(_0150_));
 sky130_fd_sc_hd__clkbuf_1 _0639_ (.A(_0150_),
    .X(_0231_));
 sky130_fd_sc_hd__inv_2 _0640_ (.A(\mem_top_track_14.DFFR_1_.Q ),
    .Y(_0227_));
 sky130_fd_sc_hd__inv_2 _0641_ (.A(\mem_top_track_14.DFFR_0_.Q ),
    .Y(_0229_));
 sky130_fd_sc_hd__clkbuf_1 _0642_ (.A(\mem_top_track_14.DFFR_0_.Q ),
    .X(_0151_));
 sky130_fd_sc_hd__clkbuf_1 _0643_ (.A(_0151_),
    .X(_0226_));
 sky130_fd_sc_hd__clkbuf_1 _0644_ (.A(\mem_top_track_14.DFFR_1_.Q ),
    .X(_0152_));
 sky130_fd_sc_hd__clkbuf_1 _0645_ (.A(_0152_),
    .X(_0224_));
 sky130_fd_sc_hd__inv_2 _0646_ (.A(\mem_top_track_14.DFFR_0_.Q ),
    .Y(_0228_));
 sky130_fd_sc_hd__clkbuf_1 _0647_ (.A(\mem_top_track_14.DFFR_0_.Q ),
    .X(_0153_));
 sky130_fd_sc_hd__clkbuf_1 _0648_ (.A(_0153_),
    .X(_0225_));
 sky130_fd_sc_hd__inv_2 _0649_ (.A(\mem_top_track_12.DFFR_1_.Q ),
    .Y(_0221_));
 sky130_fd_sc_hd__inv_2 _0650_ (.A(\mem_top_track_12.DFFR_0_.Q ),
    .Y(_0223_));
 sky130_fd_sc_hd__clkbuf_1 _0651_ (.A(\mem_top_track_12.DFFR_0_.Q ),
    .X(_0154_));
 sky130_fd_sc_hd__clkbuf_1 _0652_ (.A(_0154_),
    .X(_0220_));
 sky130_fd_sc_hd__clkbuf_1 _0653_ (.A(\mem_top_track_12.DFFR_1_.Q ),
    .X(_0155_));
 sky130_fd_sc_hd__clkbuf_1 _0654_ (.A(_0155_),
    .X(_0218_));
 sky130_fd_sc_hd__inv_2 _0655_ (.A(\mem_top_track_12.DFFR_0_.Q ),
    .Y(_0222_));
 sky130_fd_sc_hd__clkbuf_1 _0656_ (.A(\mem_top_track_12.DFFR_0_.Q ),
    .X(_0156_));
 sky130_fd_sc_hd__clkbuf_1 _0657_ (.A(_0156_),
    .X(_0219_));
 sky130_fd_sc_hd__inv_2 _0658_ (.A(\mem_top_track_10.DFFR_1_.Q ),
    .Y(_0215_));
 sky130_fd_sc_hd__inv_2 _0659_ (.A(\mem_top_track_10.DFFR_0_.Q ),
    .Y(_0217_));
 sky130_fd_sc_hd__clkbuf_1 _0660_ (.A(\mem_top_track_10.DFFR_0_.Q ),
    .X(_0157_));
 sky130_fd_sc_hd__clkbuf_1 _0661_ (.A(_0157_),
    .X(_0214_));
 sky130_fd_sc_hd__clkbuf_1 _0662_ (.A(\mem_top_track_10.DFFR_1_.Q ),
    .X(_0158_));
 sky130_fd_sc_hd__clkbuf_1 _0663_ (.A(_0158_),
    .X(_0212_));
 sky130_fd_sc_hd__inv_2 _0664_ (.A(\mem_top_track_10.DFFR_0_.Q ),
    .Y(_0216_));
 sky130_fd_sc_hd__clkbuf_1 _0665_ (.A(\mem_top_track_10.DFFR_0_.Q ),
    .X(_0159_));
 sky130_fd_sc_hd__clkbuf_1 _0666_ (.A(_0159_),
    .X(_0213_));
 sky130_fd_sc_hd__inv_2 _0667_ (.A(\mem_top_track_10.DFFR_0_.D ),
    .Y(_0209_));
 sky130_fd_sc_hd__inv_2 _0668_ (.A(\mem_top_track_8.DFFR_0_.Q ),
    .Y(_0211_));
 sky130_fd_sc_hd__clkbuf_1 _0669_ (.A(\mem_top_track_8.DFFR_0_.Q ),
    .X(_0160_));
 sky130_fd_sc_hd__clkbuf_1 _0670_ (.A(_0160_),
    .X(_0208_));
 sky130_fd_sc_hd__clkbuf_1 _0671_ (.A(\mem_top_track_10.DFFR_0_.D ),
    .X(_0161_));
 sky130_fd_sc_hd__clkbuf_1 _0672_ (.A(_0161_),
    .X(_0206_));
 sky130_fd_sc_hd__inv_2 _0673_ (.A(\mem_top_track_8.DFFR_0_.Q ),
    .Y(_0210_));
 sky130_fd_sc_hd__clkbuf_1 _0674_ (.A(\mem_top_track_8.DFFR_0_.Q ),
    .X(_0162_));
 sky130_fd_sc_hd__clkbuf_1 _0675_ (.A(_0162_),
    .X(_0207_));
 sky130_fd_sc_hd__inv_2 _0676_ (.A(\mem_top_track_6.DFFR_1_.Q ),
    .Y(_0203_));
 sky130_fd_sc_hd__inv_2 _0677_ (.A(\mem_top_track_6.DFFR_0_.Q ),
    .Y(_0205_));
 sky130_fd_sc_hd__clkbuf_1 _0678_ (.A(\mem_top_track_6.DFFR_0_.Q ),
    .X(_0163_));
 sky130_fd_sc_hd__clkbuf_1 _0679_ (.A(_0163_),
    .X(_0202_));
 sky130_fd_sc_hd__clkbuf_1 _0680_ (.A(\mem_top_track_6.DFFR_1_.Q ),
    .X(_0164_));
 sky130_fd_sc_hd__clkbuf_1 _0681_ (.A(_0164_),
    .X(_0200_));
 sky130_fd_sc_hd__inv_2 _0682_ (.A(\mem_top_track_6.DFFR_0_.Q ),
    .Y(_0204_));
 sky130_fd_sc_hd__clkbuf_1 _0683_ (.A(\mem_top_track_6.DFFR_0_.Q ),
    .X(_0165_));
 sky130_fd_sc_hd__clkbuf_1 _0684_ (.A(_0165_),
    .X(_0201_));
 sky130_fd_sc_hd__inv_2 _0685_ (.A(\mem_top_track_4.DFFR_1_.Q ),
    .Y(_0197_));
 sky130_fd_sc_hd__inv_2 _0686_ (.A(\mem_top_track_4.DFFR_0_.Q ),
    .Y(_0199_));
 sky130_fd_sc_hd__clkbuf_1 _0687_ (.A(\mem_top_track_4.DFFR_0_.Q ),
    .X(_0166_));
 sky130_fd_sc_hd__clkbuf_1 _0688_ (.A(_0166_),
    .X(_0196_));
 sky130_fd_sc_hd__clkbuf_1 _0689_ (.A(\mem_top_track_4.DFFR_1_.Q ),
    .X(_0167_));
 sky130_fd_sc_hd__clkbuf_1 _0690_ (.A(_0167_),
    .X(_0194_));
 sky130_fd_sc_hd__inv_2 _0691_ (.A(\mem_top_track_4.DFFR_0_.Q ),
    .Y(_0198_));
 sky130_fd_sc_hd__clkbuf_1 _0692_ (.A(\mem_top_track_4.DFFR_0_.Q ),
    .X(_0168_));
 sky130_fd_sc_hd__clkbuf_1 _0693_ (.A(_0168_),
    .X(_0195_));
 sky130_fd_sc_hd__inv_2 _0694_ (.A(\mem_top_track_2.DFFR_1_.Q ),
    .Y(_0191_));
 sky130_fd_sc_hd__inv_2 _0695_ (.A(\mem_top_track_2.DFFR_0_.Q ),
    .Y(_0193_));
 sky130_fd_sc_hd__clkbuf_1 _0696_ (.A(\mem_top_track_2.DFFR_1_.Q ),
    .X(_0169_));
 sky130_fd_sc_hd__clkbuf_1 _0697_ (.A(_0169_),
    .X(_0190_));
 sky130_fd_sc_hd__inv_2 _0698_ (.A(\mem_top_track_2.DFFR_0_.Q ),
    .Y(_0192_));
 sky130_fd_sc_hd__clkbuf_1 _0699_ (.A(\mem_top_track_2.DFFR_0_.Q ),
    .X(_0170_));
 sky130_fd_sc_hd__clkbuf_1 _0700_ (.A(_0170_),
    .X(_0189_));
 sky130_fd_sc_hd__clkbuf_1 _0701_ (.A(\mem_top_track_2.DFFR_0_.Q ),
    .X(_0171_));
 sky130_fd_sc_hd__clkbuf_1 _0702_ (.A(_0171_),
    .X(_0188_));
 sky130_fd_sc_hd__inv_2 _0703_ (.A(\mem_top_track_0.DFFR_0_.Q ),
    .Y(_0187_));
 sky130_fd_sc_hd__inv_2 _0704_ (.A(\mem_top_track_0.DFFR_1_.Q ),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_2 _0705_ (.A(\mem_top_track_0.DFFR_0_.Q ),
    .Y(_0186_));
 sky130_fd_sc_hd__clkbuf_1 _0706_ (.A(\mem_top_track_0.DFFR_0_.Q ),
    .X(_0172_));
 sky130_fd_sc_hd__clkbuf_1 _0707_ (.A(_0172_),
    .X(_0184_));
 sky130_fd_sc_hd__clkbuf_1 _0708_ (.A(\mem_top_track_0.DFFR_0_.Q ),
    .X(_0173_));
 sky130_fd_sc_hd__clkbuf_1 _0709_ (.A(_0173_),
    .X(_0183_));
 sky130_fd_sc_hd__inv_2 _0710_ (.A(net51),
    .Y(\mux_top_track_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0711_ (.A(net52),
    .Y(\mux_top_track_0.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0712_ (.A(\mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_top_track_0.out ));
 sky130_fd_sc_hd__inv_2 _0713_ (.A(net2),
    .Y(\mux_top_track_0.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0714_ (.A(net53),
    .Y(\mux_top_track_2.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0715_ (.A(\mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_top_track_2.out ));
 sky130_fd_sc_hd__inv_2 _0716_ (.A(net11),
    .Y(\mux_top_track_2.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0717_ (.A(\mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_top_track_4.out ));
 sky130_fd_sc_hd__inv_2 _0718_ (.A(net10),
    .Y(\mux_top_track_4.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0719_ (.A(\mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_top_track_6.out ));
 sky130_fd_sc_hd__inv_2 _0720_ (.A(net9),
    .Y(\mux_top_track_6.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0721_ (.A(\mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_top_track_8.out ));
 sky130_fd_sc_hd__inv_2 _0722_ (.A(net8),
    .Y(\mux_top_track_8.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0723_ (.A(\mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_top_track_10.out ));
 sky130_fd_sc_hd__inv_2 _0724_ (.A(net57),
    .Y(\mux_top_track_10.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0725_ (.A(net56),
    .Y(\mux_top_track_10.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0726_ (.A(net7),
    .Y(\mux_top_track_10.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0727_ (.A(\mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_top_track_12.out ));
 sky130_fd_sc_hd__inv_2 _0728_ (.A(net58),
    .Y(\mux_top_track_12.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0729_ (.A(net6),
    .Y(\mux_top_track_12.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0730_ (.A(\mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_top_track_14.out ));
 sky130_fd_sc_hd__inv_2 _0731_ (.A(net59),
    .Y(\mux_top_track_14.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0732_ (.A(net5),
    .Y(\mux_top_track_14.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0733_ (.A(\mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_top_track_16.out ));
 sky130_fd_sc_hd__inv_2 _0734_ (.A(net60),
    .Y(\mux_top_track_16.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0735_ (.A(net4),
    .Y(\mux_top_track_16.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0736_ (.A(\mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_top_track_18.out ));
 sky130_fd_sc_hd__inv_2 _0737_ (.A(net3),
    .Y(\mux_top_track_18.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0738_ (.A(\mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_top_track_36.out ));
 sky130_fd_sc_hd__inv_2 _0739_ (.A(net12),
    .Y(\mux_top_track_36.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0740_ (.A(\mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_left_track_1.out ));
 sky130_fd_sc_hd__inv_2 _0741_ (.A(net48),
    .Y(\mux_left_track_1.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0742_ (.A(net21),
    .Y(\mux_left_track_1.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0743_ (.A(net49),
    .Y(\mux_left_track_1.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0744_ (.A(\mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_left_track_3.out ));
 sky130_fd_sc_hd__inv_2 _0745_ (.A(net30),
    .Y(\mux_left_track_3.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0746_ (.A(\mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_left_track_5.out ));
 sky130_fd_sc_hd__inv_2 _0747_ (.A(net29),
    .Y(\mux_left_track_5.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0748_ (.A(\mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_left_track_7.out ));
 sky130_fd_sc_hd__inv_2 _0749_ (.A(net28),
    .Y(\mux_left_track_7.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0750_ (.A(\mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_left_track_9.out ));
 sky130_fd_sc_hd__inv_2 _0751_ (.A(net27),
    .Y(\mux_left_track_9.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0752_ (.A(\mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_left_track_11.out ));
 sky130_fd_sc_hd__inv_2 _0753_ (.A(net43),
    .Y(\mux_left_track_11.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0754_ (.A(net26),
    .Y(\mux_left_track_11.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0755_ (.A(net44),
    .Y(\mux_left_track_11.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0756_ (.A(\mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_left_track_13.out ));
 sky130_fd_sc_hd__inv_2 _0757_ (.A(net25),
    .Y(\mux_left_track_13.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0758_ (.A(net45),
    .Y(\mux_left_track_13.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0759_ (.A(\mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_left_track_15.out ));
 sky130_fd_sc_hd__inv_2 _0760_ (.A(net24),
    .Y(\mux_left_track_15.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0761_ (.A(net46),
    .Y(\mux_left_track_15.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0762_ (.A(\mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_left_track_17.out ));
 sky130_fd_sc_hd__inv_2 _0763_ (.A(net23),
    .Y(\mux_left_track_17.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0764_ (.A(net47),
    .Y(\mux_left_track_17.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0765_ (.A(\mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_left_track_19.out ));
 sky130_fd_sc_hd__inv_2 _0766_ (.A(net22),
    .Y(\mux_left_track_19.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0767_ (.A(\mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_left_track_37.out ));
 sky130_fd_sc_hd__inv_2 _0768_ (.A(net31),
    .Y(\mux_left_track_37.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0769_ (.A(\mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_top_track_20.out ));
 sky130_fd_sc_hd__inv_2 _0770_ (.A(net20),
    .Y(\mux_top_track_20.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0771_ (.A(\mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_top_track_22.out ));
 sky130_fd_sc_hd__inv_2 _0772_ (.A(net19),
    .Y(\mux_top_track_22.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0773_ (.A(\mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_top_track_24.out ));
 sky130_fd_sc_hd__inv_2 _0774_ (.A(net54),
    .Y(\mux_top_track_24.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0775_ (.A(net18),
    .Y(\mux_top_track_24.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0776_ (.A(\mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_top_track_26.out ));
 sky130_fd_sc_hd__inv_2 _0777_ (.A(net55),
    .Y(\mux_top_track_26.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0778_ (.A(net17),
    .Y(\mux_top_track_26.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0779_ (.A(\mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_top_track_28.out ));
 sky130_fd_sc_hd__inv_2 _0780_ (.A(net16),
    .Y(\mux_top_track_28.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0781_ (.A(\mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_top_track_30.out ));
 sky130_fd_sc_hd__inv_2 _0782_ (.A(net15),
    .Y(\mux_top_track_30.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0783_ (.A(\mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_top_track_32.out ));
 sky130_fd_sc_hd__inv_2 _0784_ (.A(net14),
    .Y(\mux_top_track_32.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0785_ (.A(\mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_top_track_34.out ));
 sky130_fd_sc_hd__inv_2 _0786_ (.A(net13),
    .Y(\mux_top_track_34.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0787_ (.A(\mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_left_track_21.out ));
 sky130_fd_sc_hd__inv_2 _0788_ (.A(net39),
    .Y(\mux_left_track_21.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0789_ (.A(\mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_left_track_23.out ));
 sky130_fd_sc_hd__inv_2 _0790_ (.A(net38),
    .Y(\mux_left_track_23.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0791_ (.A(net40),
    .Y(\mux_left_track_23.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0792_ (.A(\mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_left_track_25.out ));
 sky130_fd_sc_hd__inv_2 _0793_ (.A(net37),
    .Y(\mux_left_track_25.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0794_ (.A(net41),
    .Y(\mux_left_track_25.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0795_ (.A(\mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_left_track_27.out ));
 sky130_fd_sc_hd__inv_2 _0796_ (.A(net36),
    .Y(\mux_left_track_27.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0797_ (.A(net42),
    .Y(\mux_left_track_27.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0798_ (.A(\mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_left_track_29.out ));
 sky130_fd_sc_hd__inv_2 _0799_ (.A(net35),
    .Y(\mux_left_track_29.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0800_ (.A(\mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_left_track_31.out ));
 sky130_fd_sc_hd__inv_2 _0801_ (.A(net34),
    .Y(\mux_left_track_31.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0802_ (.A(\mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_left_track_33.out ));
 sky130_fd_sc_hd__inv_2 _0803_ (.A(net33),
    .Y(\mux_left_track_33.INVTX1_0_.out ));
 sky130_fd_sc_hd__clkinv_2 _0804_ (.A(\mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_left_track_35.out ));
 sky130_fd_sc_hd__inv_2 _0805_ (.A(net32),
    .Y(\mux_left_track_35.INVTX1_0_.out ));
 sky130_fd_sc_hd__buf_4 _0806_ (.A(net50),
    .X(_0174_));
 sky130_fd_sc_hd__buf_4 _0807_ (.A(_0174_),
    .X(_0175_));
 sky130_fd_sc_hd__inv_2 _0808_ (.A(_0175_),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _0809_ (.A(_0175_),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _0810_ (.A(_0175_),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _0811_ (.A(_0175_),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _0812_ (.A(_0175_),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _0813_ (.A(_0175_),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _0814_ (.A(_0175_),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _0815_ (.A(_0175_),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _0816_ (.A(_0175_),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _0817_ (.A(_0175_),
    .Y(_0064_));
 sky130_fd_sc_hd__buf_4 _0818_ (.A(_0174_),
    .X(_0176_));
 sky130_fd_sc_hd__inv_2 _0819_ (.A(_0176_),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _0820_ (.A(_0176_),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _0821_ (.A(_0176_),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _0822_ (.A(_0176_),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _0823_ (.A(_0176_),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _0824_ (.A(_0176_),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _0825_ (.A(_0176_),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _0826_ (.A(_0176_),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _0827_ (.A(_0176_),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _0828_ (.A(_0176_),
    .Y(_0074_));
 sky130_fd_sc_hd__buf_4 _0829_ (.A(_0174_),
    .X(_0177_));
 sky130_fd_sc_hd__inv_2 _0830_ (.A(_0177_),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _0831_ (.A(_0177_),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_2 _0832_ (.A(_0177_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _0833_ (.A(_0177_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _0834_ (.A(_0177_),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _0835_ (.A(_0177_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _0836_ (.A(_0177_),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _0837_ (.A(_0177_),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _0838_ (.A(_0177_),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _0839_ (.A(_0177_),
    .Y(_0008_));
 sky130_fd_sc_hd__buf_4 _0840_ (.A(_0174_),
    .X(_0178_));
 sky130_fd_sc_hd__inv_2 _0841_ (.A(_0178_),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _0842_ (.A(_0178_),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _0843_ (.A(_0178_),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _0844_ (.A(_0178_),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _0845_ (.A(_0178_),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _0846_ (.A(_0178_),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _0847_ (.A(_0178_),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _0848_ (.A(_0178_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _0849_ (.A(_0178_),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _0850_ (.A(_0178_),
    .Y(_0018_));
 sky130_fd_sc_hd__buf_4 _0851_ (.A(net50),
    .X(_0179_));
 sky130_fd_sc_hd__inv_2 _0852_ (.A(_0179_),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _0853_ (.A(_0179_),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _0854_ (.A(_0179_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _0855_ (.A(_0179_),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _0856_ (.A(_0179_),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _0857_ (.A(_0179_),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _0858_ (.A(_0179_),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _0859_ (.A(_0179_),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _0860_ (.A(_0179_),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _0861_ (.A(_0179_),
    .Y(_0028_));
 sky130_fd_sc_hd__buf_4 _0862_ (.A(net50),
    .X(_0180_));
 sky130_fd_sc_hd__inv_2 _0863_ (.A(_0180_),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _0864_ (.A(_0180_),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _0865_ (.A(_0180_),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _0866_ (.A(_0180_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _0867_ (.A(_0180_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _0868_ (.A(_0180_),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _0869_ (.A(_0180_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _0870_ (.A(_0180_),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _0871_ (.A(_0180_),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _0872_ (.A(_0180_),
    .Y(_0038_));
 sky130_fd_sc_hd__buf_4 _0873_ (.A(net50),
    .X(_0181_));
 sky130_fd_sc_hd__inv_2 _0874_ (.A(_0181_),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _0875_ (.A(_0181_),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _0876_ (.A(_0181_),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _0877_ (.A(_0181_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _0878_ (.A(_0181_),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _0879_ (.A(_0181_),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _0880_ (.A(_0181_),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _0881_ (.A(_0181_),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _0882_ (.A(_0181_),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _0883_ (.A(_0181_),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _0884_ (.A(_0174_),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _0885_ (.A(_0174_),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _0886_ (.A(_0174_),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _0887_ (.A(_0174_),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _0888_ (.A(_0174_),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _0889_ (.A(_0174_),
    .Y(_0054_));
 sky130_fd_sc_hd__dfrtp_1 _0890_ (.CLK(clknet_3_6__leaf_prog_clk),
    .D(\mem_top_track_0.DFFR_0_.Q ),
    .RESET_B(_0055_),
    .Q(\mem_top_track_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0891_ (.CLK(clknet_3_5__leaf_prog_clk),
    .D(net1),
    .RESET_B(_0056_),
    .Q(\mem_top_track_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0892_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_top_track_2.DFFR_0_.Q ),
    .RESET_B(_0057_),
    .Q(\mem_top_track_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0893_ (.CLK(clknet_3_1__leaf_prog_clk),
    .D(\mem_top_track_0.DFFR_1_.Q ),
    .RESET_B(_0058_),
    .Q(\mem_top_track_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0894_ (.CLK(clknet_3_5__leaf_prog_clk),
    .D(\mem_top_track_4.DFFR_0_.Q ),
    .RESET_B(_0059_),
    .Q(\mem_top_track_4.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0895_ (.CLK(clknet_3_1__leaf_prog_clk),
    .D(\mem_top_track_2.DFFR_1_.Q ),
    .RESET_B(_0060_),
    .Q(\mem_top_track_4.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0896_ (.CLK(clknet_3_2__leaf_prog_clk),
    .D(\mem_top_track_6.DFFR_0_.Q ),
    .RESET_B(_0061_),
    .Q(\mem_top_track_6.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0897_ (.CLK(clknet_3_1__leaf_prog_clk),
    .D(\mem_top_track_4.DFFR_1_.Q ),
    .RESET_B(_0062_),
    .Q(\mem_top_track_6.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0898_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_top_track_8.DFFR_0_.Q ),
    .RESET_B(_0063_),
    .Q(\mem_top_track_10.DFFR_0_.D ));
 sky130_fd_sc_hd__dfrtp_4 _0899_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_top_track_6.DFFR_1_.Q ),
    .RESET_B(_0064_),
    .Q(\mem_top_track_8.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0900_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_top_track_10.DFFR_0_.Q ),
    .RESET_B(_0065_),
    .Q(\mem_top_track_10.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0901_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_top_track_10.DFFR_0_.D ),
    .RESET_B(_0066_),
    .Q(\mem_top_track_10.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0902_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_top_track_12.DFFR_0_.Q ),
    .RESET_B(_0067_),
    .Q(\mem_top_track_12.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0903_ (.CLK(clknet_3_1__leaf_prog_clk),
    .D(\mem_top_track_10.DFFR_1_.Q ),
    .RESET_B(_0068_),
    .Q(\mem_top_track_12.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0904_ (.CLK(clknet_3_5__leaf_prog_clk),
    .D(\mem_top_track_14.DFFR_0_.Q ),
    .RESET_B(_0069_),
    .Q(\mem_top_track_14.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0905_ (.CLK(clknet_3_3__leaf_prog_clk),
    .D(\mem_top_track_12.DFFR_1_.Q ),
    .RESET_B(_0070_),
    .Q(\mem_top_track_14.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0906_ (.CLK(clknet_3_5__leaf_prog_clk),
    .D(\mem_top_track_16.DFFR_0_.Q ),
    .RESET_B(_0071_),
    .Q(\mem_top_track_16.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0907_ (.CLK(clknet_3_5__leaf_prog_clk),
    .D(\mem_top_track_14.DFFR_1_.Q ),
    .RESET_B(_0072_),
    .Q(\mem_top_track_16.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0908_ (.CLK(clknet_3_5__leaf_prog_clk),
    .D(\mem_top_track_18.DFFR_0_.Q ),
    .RESET_B(_0073_),
    .Q(\mem_top_track_18.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0909_ (.CLK(clknet_3_4__leaf_prog_clk),
    .D(\mem_top_track_16.DFFR_1_.Q ),
    .RESET_B(_0074_),
    .Q(\mem_top_track_18.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0910_ (.CLK(clknet_3_1__leaf_prog_clk),
    .D(\mem_top_track_36.DFFR_0_.Q ),
    .RESET_B(_0075_),
    .Q(\mem_left_track_1.DFFR_0_.D ));
 sky130_fd_sc_hd__dfrtp_4 _0911_ (.CLK(clknet_3_4__leaf_prog_clk),
    .D(\mem_top_track_34.DFFR_1_.Q ),
    .RESET_B(_0000_),
    .Q(\mem_top_track_36.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0912_ (.CLK(clknet_3_4__leaf_prog_clk),
    .D(\mem_left_track_1.DFFR_0_.Q ),
    .RESET_B(_0001_),
    .Q(\mem_left_track_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0913_ (.CLK(clknet_3_1__leaf_prog_clk),
    .D(\mem_left_track_1.DFFR_0_.D ),
    .RESET_B(_0002_),
    .Q(\mem_left_track_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0914_ (.CLK(clknet_3_4__leaf_prog_clk),
    .D(\mem_left_track_3.DFFR_0_.Q ),
    .RESET_B(_0003_),
    .Q(\mem_left_track_3.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0915_ (.CLK(clknet_3_6__leaf_prog_clk),
    .D(\mem_left_track_1.DFFR_1_.Q ),
    .RESET_B(_0004_),
    .Q(\mem_left_track_3.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0916_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_left_track_5.DFFR_0_.Q ),
    .RESET_B(_0005_),
    .Q(\mem_left_track_5.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0917_ (.CLK(clknet_3_1__leaf_prog_clk),
    .D(\mem_left_track_3.DFFR_1_.Q ),
    .RESET_B(_0006_),
    .Q(\mem_left_track_5.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0918_ (.CLK(clknet_3_1__leaf_prog_clk),
    .D(\mem_left_track_7.DFFR_0_.Q ),
    .RESET_B(_0007_),
    .Q(\mem_left_track_7.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0919_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_left_track_5.DFFR_1_.Q ),
    .RESET_B(_0008_),
    .Q(\mem_left_track_7.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0920_ (.CLK(clknet_3_4__leaf_prog_clk),
    .D(\mem_left_track_9.DFFR_0_.Q ),
    .RESET_B(_0009_),
    .Q(\mem_left_track_11.DFFR_0_.D ));
 sky130_fd_sc_hd__dfrtp_2 _0921_ (.CLK(clknet_3_4__leaf_prog_clk),
    .D(\mem_left_track_7.DFFR_1_.Q ),
    .RESET_B(_0010_),
    .Q(\mem_left_track_9.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0922_ (.CLK(clknet_3_4__leaf_prog_clk),
    .D(\mem_left_track_11.DFFR_0_.Q ),
    .RESET_B(_0011_),
    .Q(\mem_left_track_11.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0923_ (.CLK(clknet_3_5__leaf_prog_clk),
    .D(\mem_left_track_11.DFFR_0_.D ),
    .RESET_B(_0012_),
    .Q(\mem_left_track_11.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0924_ (.CLK(clknet_3_4__leaf_prog_clk),
    .D(\mem_left_track_13.DFFR_0_.Q ),
    .RESET_B(_0013_),
    .Q(\mem_left_track_13.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0925_ (.CLK(clknet_3_4__leaf_prog_clk),
    .D(\mem_left_track_11.DFFR_1_.Q ),
    .RESET_B(_0014_),
    .Q(\mem_left_track_13.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0926_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_left_track_15.DFFR_0_.Q ),
    .RESET_B(_0015_),
    .Q(\mem_left_track_15.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0927_ (.CLK(clknet_3_6__leaf_prog_clk),
    .D(\mem_left_track_13.DFFR_1_.Q ),
    .RESET_B(_0016_),
    .Q(\mem_left_track_15.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0928_ (.CLK(clknet_3_5__leaf_prog_clk),
    .D(\mem_left_track_17.DFFR_0_.Q ),
    .RESET_B(_0017_),
    .Q(\mem_left_track_17.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0929_ (.CLK(clknet_3_1__leaf_prog_clk),
    .D(\mem_left_track_15.DFFR_1_.Q ),
    .RESET_B(_0018_),
    .Q(\mem_left_track_17.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0930_ (.CLK(clknet_3_3__leaf_prog_clk),
    .D(\mem_left_track_19.DFFR_0_.Q ),
    .RESET_B(_0019_),
    .Q(\mem_left_track_19.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0931_ (.CLK(clknet_3_7__leaf_prog_clk),
    .D(\mem_left_track_17.DFFR_1_.Q ),
    .RESET_B(_0020_),
    .Q(\mem_left_track_19.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0932_ (.CLK(clknet_3_7__leaf_prog_clk),
    .D(\mem_left_track_37.DFFR_0_.Q ),
    .RESET_B(_0021_),
    .Q(net61));
 sky130_fd_sc_hd__dfrtp_2 _0933_ (.CLK(clknet_3_6__leaf_prog_clk),
    .D(\mem_left_track_35.DFFR_1_.Q ),
    .RESET_B(_0022_),
    .Q(\mem_left_track_37.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0934_ (.CLK(clknet_3_3__leaf_prog_clk),
    .D(\mem_top_track_20.DFFR_0_.Q ),
    .RESET_B(_0023_),
    .Q(\mem_top_track_20.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0935_ (.CLK(clknet_3_3__leaf_prog_clk),
    .D(\mem_top_track_18.DFFR_1_.Q ),
    .RESET_B(_0024_),
    .Q(\mem_top_track_20.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0936_ (.CLK(clknet_3_2__leaf_prog_clk),
    .D(\mem_top_track_22.DFFR_0_.Q ),
    .RESET_B(_0025_),
    .Q(\mem_top_track_22.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0937_ (.CLK(clknet_3_2__leaf_prog_clk),
    .D(\mem_top_track_20.DFFR_1_.Q ),
    .RESET_B(_0026_),
    .Q(\mem_top_track_22.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0938_ (.CLK(clknet_3_5__leaf_prog_clk),
    .D(\mem_top_track_24.DFFR_0_.Q ),
    .RESET_B(_0027_),
    .Q(\mem_top_track_24.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0939_ (.CLK(clknet_3_2__leaf_prog_clk),
    .D(\mem_top_track_22.DFFR_1_.Q ),
    .RESET_B(_0028_),
    .Q(\mem_top_track_24.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0940_ (.CLK(clknet_3_6__leaf_prog_clk),
    .D(\mem_top_track_26.DFFR_0_.Q ),
    .RESET_B(_0029_),
    .Q(\mem_top_track_26.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0941_ (.CLK(clknet_3_5__leaf_prog_clk),
    .D(\mem_top_track_24.DFFR_1_.Q ),
    .RESET_B(_0030_),
    .Q(\mem_top_track_26.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0942_ (.CLK(clknet_3_7__leaf_prog_clk),
    .D(\mem_top_track_28.DFFR_0_.Q ),
    .RESET_B(_0031_),
    .Q(\mem_top_track_28.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0943_ (.CLK(clknet_3_6__leaf_prog_clk),
    .D(\mem_top_track_26.DFFR_1_.Q ),
    .RESET_B(_0032_),
    .Q(\mem_top_track_28.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0944_ (.CLK(clknet_3_2__leaf_prog_clk),
    .D(\mem_top_track_30.DFFR_0_.Q ),
    .RESET_B(_0033_),
    .Q(\mem_top_track_30.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0945_ (.CLK(clknet_3_6__leaf_prog_clk),
    .D(\mem_top_track_28.DFFR_1_.Q ),
    .RESET_B(_0034_),
    .Q(\mem_top_track_30.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0946_ (.CLK(clknet_3_6__leaf_prog_clk),
    .D(\mem_top_track_32.DFFR_0_.Q ),
    .RESET_B(_0035_),
    .Q(\mem_top_track_32.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0947_ (.CLK(clknet_3_1__leaf_prog_clk),
    .D(\mem_top_track_30.DFFR_1_.Q ),
    .RESET_B(_0036_),
    .Q(\mem_top_track_32.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0948_ (.CLK(clknet_3_3__leaf_prog_clk),
    .D(\mem_top_track_34.DFFR_0_.Q ),
    .RESET_B(_0037_),
    .Q(\mem_top_track_34.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0949_ (.CLK(clknet_3_6__leaf_prog_clk),
    .D(\mem_top_track_32.DFFR_1_.Q ),
    .RESET_B(_0038_),
    .Q(\mem_top_track_34.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0950_ (.CLK(clknet_3_2__leaf_prog_clk),
    .D(\mem_left_track_21.DFFR_0_.Q ),
    .RESET_B(_0039_),
    .Q(\mem_left_track_21.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0951_ (.CLK(clknet_3_2__leaf_prog_clk),
    .D(\mem_left_track_19.DFFR_1_.Q ),
    .RESET_B(_0040_),
    .Q(\mem_left_track_21.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0952_ (.CLK(clknet_3_6__leaf_prog_clk),
    .D(\mem_left_track_23.DFFR_0_.Q ),
    .RESET_B(_0041_),
    .Q(\mem_left_track_23.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0953_ (.CLK(clknet_3_3__leaf_prog_clk),
    .D(\mem_left_track_21.DFFR_1_.Q ),
    .RESET_B(_0042_),
    .Q(\mem_left_track_23.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0954_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_left_track_25.DFFR_0_.Q ),
    .RESET_B(_0043_),
    .Q(\mem_left_track_25.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0955_ (.CLK(clknet_3_0__leaf_prog_clk),
    .D(\mem_left_track_23.DFFR_1_.Q ),
    .RESET_B(_0044_),
    .Q(\mem_left_track_25.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0956_ (.CLK(clknet_3_6__leaf_prog_clk),
    .D(\mem_left_track_27.DFFR_0_.Q ),
    .RESET_B(_0045_),
    .Q(\mem_left_track_27.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0957_ (.CLK(clknet_3_3__leaf_prog_clk),
    .D(\mem_left_track_25.DFFR_1_.Q ),
    .RESET_B(_0046_),
    .Q(\mem_left_track_27.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0958_ (.CLK(clknet_3_7__leaf_prog_clk),
    .D(\mem_left_track_29.DFFR_0_.Q ),
    .RESET_B(_0047_),
    .Q(\mem_left_track_29.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0959_ (.CLK(clknet_3_7__leaf_prog_clk),
    .D(\mem_left_track_27.DFFR_1_.Q ),
    .RESET_B(_0048_),
    .Q(\mem_left_track_29.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0960_ (.CLK(clknet_3_3__leaf_prog_clk),
    .D(\mem_left_track_31.DFFR_0_.Q ),
    .RESET_B(_0049_),
    .Q(\mem_left_track_31.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0961_ (.CLK(clknet_3_3__leaf_prog_clk),
    .D(\mem_left_track_29.DFFR_1_.Q ),
    .RESET_B(_0050_),
    .Q(\mem_left_track_31.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0962_ (.CLK(clknet_3_7__leaf_prog_clk),
    .D(\mem_left_track_33.DFFR_0_.Q ),
    .RESET_B(_0051_),
    .Q(\mem_left_track_33.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0963_ (.CLK(clknet_3_6__leaf_prog_clk),
    .D(\mem_left_track_31.DFFR_1_.Q ),
    .RESET_B(_0052_),
    .Q(\mem_left_track_33.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0964_ (.CLK(clknet_3_7__leaf_prog_clk),
    .D(\mem_left_track_35.DFFR_0_.Q ),
    .RESET_B(_0053_),
    .Q(\mem_left_track_35.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0965_ (.CLK(clknet_3_7__leaf_prog_clk),
    .D(\mem_left_track_33.DFFR_1_.Q ),
    .RESET_B(_0054_),
    .Q(\mem_left_track_35.DFFR_0_.Q ));
 sky130_fd_sc_hd__conb_1 _1049__101 (.HI(net101));
 sky130_fd_sc_hd__conb_1 _1055__102 (.HI(net102));
 sky130_fd_sc_hd__conb_1 _1061__103 (.HI(net103));
 sky130_fd_sc_hd__conb_1 _1067__104 (.HI(net104));
 sky130_fd_sc_hd__conb_1 _1073__105 (.HI(net105));
 sky130_fd_sc_hd__conb_1 _1079__106 (.HI(net106));
 sky130_fd_sc_hd__conb_1 _1085__107 (.HI(net107));
 sky130_fd_sc_hd__conb_1 _1091__108 (.HI(net108));
 sky130_fd_sc_hd__conb_1 _1097__109 (.HI(net109));
 sky130_fd_sc_hd__conb_1 _1103__110 (.HI(net110));
 sky130_fd_sc_hd__conb_1 _1109__111 (.HI(net111));
 sky130_fd_sc_hd__conb_1 _1115__112 (.HI(net112));
 sky130_fd_sc_hd__conb_1 _1121__113 (.HI(net113));
 sky130_fd_sc_hd__conb_1 _1127__114 (.HI(net114));
 sky130_fd_sc_hd__conb_1 _1133__115 (.HI(net115));
 sky130_fd_sc_hd__conb_1 _1139__116 (.HI(net116));
 sky130_fd_sc_hd__conb_1 _1145__117 (.HI(net117));
 sky130_fd_sc_hd__conb_1 _1151__118 (.HI(net118));
 sky130_fd_sc_hd__conb_1 _1157__119 (.HI(net119));
 sky130_fd_sc_hd__conb_1 _1163__120 (.HI(net120));
 sky130_fd_sc_hd__conb_1 _1169__121 (.HI(net121));
 sky130_fd_sc_hd__conb_1 _1174__122 (.HI(net122));
 sky130_fd_sc_hd__conb_1 _1178__123 (.HI(net123));
 sky130_fd_sc_hd__conb_1 _1182__124 (.HI(net124));
 sky130_fd_sc_hd__conb_1 _1186__125 (.HI(net125));
 sky130_fd_sc_hd__conb_1 _1190__126 (.HI(net126));
 sky130_fd_sc_hd__conb_1 _1194__127 (.HI(net127));
 sky130_fd_sc_hd__conb_1 _1198__128 (.HI(net128));
 sky130_fd_sc_hd__conb_1 _1202__129 (.HI(net129));
 sky130_fd_sc_hd__conb_1 _1206__130 (.HI(net130));
 sky130_fd_sc_hd__conb_1 _1210__131 (.HI(net131));
 sky130_fd_sc_hd__conb_1 _1214__132 (.HI(net132));
 sky130_fd_sc_hd__conb_1 _1218__133 (.HI(net133));
 sky130_fd_sc_hd__conb_1 _1222__134 (.HI(net134));
 sky130_fd_sc_hd__conb_1 _1226__135 (.HI(net135));
 sky130_fd_sc_hd__conb_1 _1230__136 (.HI(net136));
 sky130_fd_sc_hd__conb_1 _1234__137 (.HI(net137));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_prog_clk (.A(prog_clk),
    .X(clknet_0_prog_clk));
 sky130_fd_sc_hd__clkbuf_1 _1004_ (.A(\mux_left_track_37.out ),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 _1005_ (.A(\mux_left_track_35.out ),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 _1006_ (.A(\mux_left_track_33.out ),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 _1007_ (.A(\mux_left_track_31.out ),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 _1008_ (.A(\mux_left_track_29.out ),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 _1009_ (.A(\mux_left_track_27.out ),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 _1010_ (.A(\mux_left_track_25.out ),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 _1011_ (.A(\mux_left_track_23.out ),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 _1012_ (.A(\mux_left_track_21.out ),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 _1013_ (.A(\mux_left_track_19.out ),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _1014_ (.A(\mux_left_track_17.out ),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _1015_ (.A(\mux_left_track_15.out ),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 _1016_ (.A(\mux_left_track_13.out ),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 _1017_ (.A(\mux_left_track_11.out ),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _1018_ (.A(\mux_left_track_9.out ),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _1019_ (.A(\mux_left_track_7.out ),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 _1020_ (.A(\mux_left_track_5.out ),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 _1021_ (.A(\mux_left_track_3.out ),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 _1022_ (.A(\mux_left_track_1.out ),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 _1023_ (.A(\mux_top_track_36.out ),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 _1024_ (.A(\mux_top_track_34.out ),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 _1025_ (.A(\mux_top_track_32.out ),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 _1026_ (.A(\mux_top_track_30.out ),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 _1027_ (.A(\mux_top_track_28.out ),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 _1028_ (.A(\mux_top_track_26.out ),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 _1029_ (.A(\mux_top_track_24.out ),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 _1030_ (.A(\mux_top_track_22.out ),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 _1031_ (.A(\mux_top_track_20.out ),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 _1032_ (.A(\mux_top_track_18.out ),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 _1033_ (.A(\mux_top_track_16.out ),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 _1034_ (.A(\mux_top_track_14.out ),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 _1035_ (.A(\mux_top_track_12.out ),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 _1036_ (.A(\mux_top_track_10.out ),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 _1037_ (.A(\mux_top_track_8.out ),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 _1038_ (.A(\mux_top_track_6.out ),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 _1039_ (.A(\mux_top_track_4.out ),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 _1040_ (.A(\mux_top_track_2.out ),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 _1041_ (.A(\mux_top_track_0.out ),
    .X(net81));
 sky130_fd_sc_hd__ebufn_2 _1042_ (.A(\mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0182_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1043_ (.A(net100),
    .TE_B(_0183_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1044_ (.A(\mux_top_track_0.INVTX1_1_.out ),
    .TE_B(_0184_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1045_ (.A(\mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0185_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1046_ (.A(\mux_top_track_0.INVTX1_0_.out ),
    .TE_B(_0186_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1047_ (.A(\mux_top_track_0.INVTX1_2_.out ),
    .TE_B(_0187_),
    .Z(\mux_top_track_0.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1048_ (.A(\mux_top_track_2.INVTX1_1_.out ),
    .TE_B(_0188_),
    .Z(\mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1049_ (.A(net101),
    .TE_B(_0189_),
    .Z(\mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1050_ (.A(\mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0190_),
    .Z(\mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1051_ (.A(\mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0191_),
    .Z(\mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1052_ (.A(\mux_top_track_2.INVTX1_2_.out ),
    .TE_B(_0192_),
    .Z(\mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1053_ (.A(\mux_top_track_0.INVTX1_1_.out ),
    .TE_B(_0193_),
    .Z(\mux_top_track_2.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1054_ (.A(\mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0194_),
    .Z(\mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1055_ (.A(net102),
    .TE_B(_0195_),
    .Z(\mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1056_ (.A(\mux_top_track_24.INVTX1_0_.out ),
    .TE_B(_0196_),
    .Z(\mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1057_ (.A(\mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0197_),
    .Z(\mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1058_ (.A(\mux_top_track_4.INVTX1_2_.out ),
    .TE_B(_0198_),
    .Z(\mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1059_ (.A(\mux_top_track_2.INVTX1_1_.out ),
    .TE_B(_0199_),
    .Z(\mux_top_track_4.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1060_ (.A(\mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0200_),
    .Z(\mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1061_ (.A(net103),
    .TE_B(_0201_),
    .Z(\mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1062_ (.A(\mux_top_track_26.INVTX1_0_.out ),
    .TE_B(_0202_),
    .Z(\mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1063_ (.A(\mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0203_),
    .Z(\mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1064_ (.A(\mux_top_track_6.INVTX1_2_.out ),
    .TE_B(_0204_),
    .Z(\mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1065_ (.A(\mux_top_track_24.INVTX1_0_.out ),
    .TE_B(_0205_),
    .Z(\mux_top_track_6.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1066_ (.A(\mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0206_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1067_ (.A(net104),
    .TE_B(_0207_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1068_ (.A(\mux_top_track_10.INVTX1_0_.out ),
    .TE_B(_0208_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1069_ (.A(\mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0209_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1070_ (.A(\mux_top_track_8.INVTX1_2_.out ),
    .TE_B(_0210_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1071_ (.A(\mux_top_track_26.INVTX1_0_.out ),
    .TE_B(_0211_),
    .Z(\mux_top_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1072_ (.A(\mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0212_),
    .Z(\mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1073_ (.A(net105),
    .TE_B(_0213_),
    .Z(\mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1074_ (.A(\mux_top_track_10.INVTX1_1_.out ),
    .TE_B(_0214_),
    .Z(\mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1075_ (.A(\mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0215_),
    .Z(\mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1076_ (.A(\mux_top_track_10.INVTX1_2_.out ),
    .TE_B(_0216_),
    .Z(\mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1077_ (.A(\mux_top_track_10.INVTX1_0_.out ),
    .TE_B(_0217_),
    .Z(\mux_top_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1078_ (.A(\mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0218_),
    .Z(\mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1079_ (.A(net106),
    .TE_B(_0219_),
    .Z(\mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1080_ (.A(\mux_top_track_12.INVTX1_1_.out ),
    .TE_B(_0220_),
    .Z(\mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1081_ (.A(\mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0221_),
    .Z(\mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1082_ (.A(\mux_top_track_12.INVTX1_2_.out ),
    .TE_B(_0222_),
    .Z(\mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1083_ (.A(\mux_top_track_10.INVTX1_1_.out ),
    .TE_B(_0223_),
    .Z(\mux_top_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1084_ (.A(\mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0224_),
    .Z(\mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1085_ (.A(net107),
    .TE_B(_0225_),
    .Z(\mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1086_ (.A(\mux_top_track_14.INVTX1_1_.out ),
    .TE_B(_0226_),
    .Z(\mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1087_ (.A(\mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0227_),
    .Z(\mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1088_ (.A(\mux_top_track_14.INVTX1_2_.out ),
    .TE_B(_0228_),
    .Z(\mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1089_ (.A(\mux_top_track_12.INVTX1_1_.out ),
    .TE_B(_0229_),
    .Z(\mux_top_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1090_ (.A(\mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0230_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1091_ (.A(net108),
    .TE_B(_0231_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1092_ (.A(\mux_top_track_16.INVTX1_1_.out ),
    .TE_B(_0232_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1093_ (.A(\mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0233_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1094_ (.A(\mux_top_track_16.INVTX1_2_.out ),
    .TE_B(_0234_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1095_ (.A(\mux_top_track_14.INVTX1_1_.out ),
    .TE_B(_0235_),
    .Z(\mux_top_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1096_ (.A(\mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0236_),
    .Z(\mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1097_ (.A(net109),
    .TE_B(_0237_),
    .Z(\mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1098_ (.A(\mux_top_track_16.INVTX1_1_.out ),
    .TE_B(_0238_),
    .Z(\mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1099_ (.A(\mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0239_),
    .Z(\mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1100_ (.A(\mux_top_track_18.INVTX1_2_.out ),
    .TE_B(_0240_),
    .Z(\mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1101_ (.A(\mux_top_track_0.INVTX1_0_.out ),
    .TE_B(_0241_),
    .Z(\mux_top_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1102_ (.A(\mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0242_),
    .Z(\mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1103_ (.A(net110),
    .TE_B(_0243_),
    .Z(\mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1104_ (.A(\mux_top_track_16.INVTX1_1_.out ),
    .TE_B(_0244_),
    .Z(\mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1105_ (.A(\mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0245_),
    .Z(\mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1106_ (.A(\mux_top_track_36.INVTX1_2_.out ),
    .TE_B(_0246_),
    .Z(\mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1107_ (.A(\mux_top_track_0.INVTX1_0_.out ),
    .TE_B(_0247_),
    .Z(\mux_top_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1108_ (.A(\mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0248_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1109_ (.A(net111),
    .TE_B(_0249_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1110_ (.A(\mux_left_track_1.INVTX1_1_.out ),
    .TE_B(_0250_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1111_ (.A(\mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0251_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1112_ (.A(\mux_left_track_1.INVTX1_2_.out ),
    .TE_B(_0252_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1113_ (.A(\mux_left_track_1.INVTX1_0_.out ),
    .TE_B(_0253_),
    .Z(\mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1114_ (.A(\mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0254_),
    .Z(\mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1115_ (.A(net112),
    .TE_B(_0255_),
    .Z(\mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1116_ (.A(\mux_left_track_1.INVTX1_2_.out ),
    .TE_B(_0256_),
    .Z(\mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1117_ (.A(\mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0257_),
    .Z(\mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1118_ (.A(\mux_left_track_23.INVTX1_1_.out ),
    .TE_B(_0258_),
    .Z(\mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1119_ (.A(\mux_left_track_3.INVTX1_0_.out ),
    .TE_B(_0259_),
    .Z(\mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1120_ (.A(\mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0260_),
    .Z(\mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1121_ (.A(net113),
    .TE_B(_0261_),
    .Z(\mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1122_ (.A(\mux_left_track_23.INVTX1_1_.out ),
    .TE_B(_0262_),
    .Z(\mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1123_ (.A(\mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0263_),
    .Z(\mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1124_ (.A(\mux_left_track_25.INVTX1_1_.out ),
    .TE_B(_0264_),
    .Z(\mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1125_ (.A(\mux_left_track_5.INVTX1_0_.out ),
    .TE_B(_0265_),
    .Z(\mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1126_ (.A(\mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0266_),
    .Z(\mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1127_ (.A(net114),
    .TE_B(_0267_),
    .Z(\mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1128_ (.A(\mux_left_track_25.INVTX1_1_.out ),
    .TE_B(_0268_),
    .Z(\mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1129_ (.A(\mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0269_),
    .Z(\mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1130_ (.A(\mux_left_track_27.INVTX1_1_.out ),
    .TE_B(_0270_),
    .Z(\mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1131_ (.A(\mux_left_track_7.INVTX1_0_.out ),
    .TE_B(_0271_),
    .Z(\mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1132_ (.A(\mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0272_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1133_ (.A(net115),
    .TE_B(_0273_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1134_ (.A(\mux_left_track_27.INVTX1_1_.out ),
    .TE_B(_0274_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1135_ (.A(\mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0275_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1136_ (.A(\mux_left_track_11.INVTX1_1_.out ),
    .TE_B(_0276_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1137_ (.A(\mux_left_track_9.INVTX1_0_.out ),
    .TE_B(_0277_),
    .Z(\mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1138_ (.A(\mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0278_),
    .Z(\mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1139_ (.A(net116),
    .TE_B(_0279_),
    .Z(\mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1140_ (.A(\mux_left_track_11.INVTX1_1_.out ),
    .TE_B(_0280_),
    .Z(\mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1141_ (.A(\mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0281_),
    .Z(\mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1142_ (.A(\mux_left_track_11.INVTX1_2_.out ),
    .TE_B(_0282_),
    .Z(\mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1143_ (.A(\mux_left_track_11.INVTX1_0_.out ),
    .TE_B(_0283_),
    .Z(\mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1144_ (.A(\mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0284_),
    .Z(\mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1145_ (.A(net117),
    .TE_B(_0285_),
    .Z(\mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1146_ (.A(\mux_left_track_11.INVTX1_2_.out ),
    .TE_B(_0286_),
    .Z(\mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1147_ (.A(\mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0287_),
    .Z(\mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1148_ (.A(\mux_left_track_13.INVTX1_2_.out ),
    .TE_B(_0288_),
    .Z(\mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1149_ (.A(\mux_left_track_13.INVTX1_0_.out ),
    .TE_B(_0289_),
    .Z(\mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1150_ (.A(\mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0290_),
    .Z(\mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1151_ (.A(net118),
    .TE_B(_0291_),
    .Z(\mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1152_ (.A(\mux_left_track_13.INVTX1_2_.out ),
    .TE_B(_0292_),
    .Z(\mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1153_ (.A(\mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0293_),
    .Z(\mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1154_ (.A(\mux_left_track_15.INVTX1_2_.out ),
    .TE_B(_0294_),
    .Z(\mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1155_ (.A(\mux_left_track_15.INVTX1_0_.out ),
    .TE_B(_0295_),
    .Z(\mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1156_ (.A(\mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0296_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1157_ (.A(net119),
    .TE_B(_0297_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1158_ (.A(\mux_left_track_15.INVTX1_2_.out ),
    .TE_B(_0298_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1159_ (.A(\mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0299_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1160_ (.A(\mux_left_track_17.INVTX1_2_.out ),
    .TE_B(_0300_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1161_ (.A(\mux_left_track_17.INVTX1_0_.out ),
    .TE_B(_0301_),
    .Z(\mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1162_ (.A(\mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0302_),
    .Z(\mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1163_ (.A(net120),
    .TE_B(_0303_),
    .Z(\mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1164_ (.A(\mux_left_track_1.INVTX1_1_.out ),
    .TE_B(_0304_),
    .Z(\mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1165_ (.A(\mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0305_),
    .Z(\mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1166_ (.A(\mux_left_track_17.INVTX1_2_.out ),
    .TE_B(_0306_),
    .Z(\mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1167_ (.A(\mux_left_track_19.INVTX1_0_.out ),
    .TE_B(_0307_),
    .Z(\mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1168_ (.A(\mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0308_),
    .Z(\mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1169_ (.A(net121),
    .TE_B(_0309_),
    .Z(\mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1170_ (.A(\mux_left_track_1.INVTX1_1_.out ),
    .TE_B(_0310_),
    .Z(\mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1171_ (.A(\mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0311_),
    .Z(\mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1172_ (.A(\mux_left_track_17.INVTX1_2_.out ),
    .TE_B(_0312_),
    .Z(\mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1173_ (.A(\mux_left_track_37.INVTX1_0_.out ),
    .TE_B(_0313_),
    .Z(\mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1174_ (.A(net122),
    .TE_B(_0314_),
    .Z(\mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1175_ (.A(\mux_top_track_20.INVTX1_1_.out ),
    .TE_B(_0315_),
    .Z(\mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1176_ (.A(\mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0316_),
    .Z(\mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1177_ (.A(\mux_top_track_0.INVTX1_1_.out ),
    .TE_B(_0317_),
    .Z(\mux_top_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1178_ (.A(net123),
    .TE_B(_0318_),
    .Z(\mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1179_ (.A(\mux_top_track_22.INVTX1_1_.out ),
    .TE_B(_0319_),
    .Z(\mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1180_ (.A(\mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0320_),
    .Z(\mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1181_ (.A(\mux_top_track_2.INVTX1_1_.out ),
    .TE_B(_0321_),
    .Z(\mux_top_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1182_ (.A(net124),
    .TE_B(_0322_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1183_ (.A(\mux_top_track_24.INVTX1_1_.out ),
    .TE_B(_0323_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1184_ (.A(\mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0324_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1185_ (.A(\mux_top_track_24.INVTX1_0_.out ),
    .TE_B(_0325_),
    .Z(\mux_top_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1186_ (.A(net125),
    .TE_B(_0326_),
    .Z(\mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1187_ (.A(\mux_top_track_26.INVTX1_1_.out ),
    .TE_B(_0327_),
    .Z(\mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1188_ (.A(\mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0328_),
    .Z(\mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1189_ (.A(\mux_top_track_26.INVTX1_0_.out ),
    .TE_B(_0329_),
    .Z(\mux_top_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1190_ (.A(net126),
    .TE_B(_0330_),
    .Z(\mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1191_ (.A(\mux_top_track_28.INVTX1_1_.out ),
    .TE_B(_0331_),
    .Z(\mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1192_ (.A(\mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0332_),
    .Z(\mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1193_ (.A(\mux_top_track_10.INVTX1_0_.out ),
    .TE_B(_0333_),
    .Z(\mux_top_track_28.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1194_ (.A(net127),
    .TE_B(_0334_),
    .Z(\mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1195_ (.A(\mux_top_track_30.INVTX1_1_.out ),
    .TE_B(_0335_),
    .Z(\mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1196_ (.A(\mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0336_),
    .Z(\mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1197_ (.A(\mux_top_track_10.INVTX1_1_.out ),
    .TE_B(_0337_),
    .Z(\mux_top_track_30.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1198_ (.A(net128),
    .TE_B(_0338_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1199_ (.A(\mux_top_track_32.INVTX1_1_.out ),
    .TE_B(_0339_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1200_ (.A(\mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0340_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1201_ (.A(\mux_top_track_12.INVTX1_1_.out ),
    .TE_B(_0341_),
    .Z(\mux_top_track_32.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1202_ (.A(net129),
    .TE_B(_0342_),
    .Z(\mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1203_ (.A(\mux_top_track_34.INVTX1_1_.out ),
    .TE_B(_0343_),
    .Z(\mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1204_ (.A(\mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0344_),
    .Z(\mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1205_ (.A(\mux_top_track_14.INVTX1_1_.out ),
    .TE_B(_0345_),
    .Z(\mux_top_track_34.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1206_ (.A(net130),
    .TE_B(_0346_),
    .Z(\mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1207_ (.A(\mux_left_track_1.INVTX1_2_.out ),
    .TE_B(_0347_),
    .Z(\mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1208_ (.A(\mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0348_),
    .Z(\mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1209_ (.A(\mux_left_track_21.INVTX1_0_.out ),
    .TE_B(_0349_),
    .Z(\mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1210_ (.A(net131),
    .TE_B(_0350_),
    .Z(\mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1211_ (.A(\mux_left_track_23.INVTX1_1_.out ),
    .TE_B(_0351_),
    .Z(\mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1212_ (.A(\mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0352_),
    .Z(\mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1213_ (.A(\mux_left_track_23.INVTX1_0_.out ),
    .TE_B(_0353_),
    .Z(\mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1214_ (.A(net132),
    .TE_B(_0354_),
    .Z(\mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1215_ (.A(\mux_left_track_25.INVTX1_1_.out ),
    .TE_B(_0355_),
    .Z(\mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1216_ (.A(\mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0356_),
    .Z(\mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1217_ (.A(\mux_left_track_25.INVTX1_0_.out ),
    .TE_B(_0357_),
    .Z(\mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1218_ (.A(net133),
    .TE_B(_0358_),
    .Z(\mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1219_ (.A(\mux_left_track_27.INVTX1_1_.out ),
    .TE_B(_0359_),
    .Z(\mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1220_ (.A(\mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0360_),
    .Z(\mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1221_ (.A(\mux_left_track_27.INVTX1_0_.out ),
    .TE_B(_0361_),
    .Z(\mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1222_ (.A(net134),
    .TE_B(_0362_),
    .Z(\mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1223_ (.A(\mux_left_track_11.INVTX1_1_.out ),
    .TE_B(_0363_),
    .Z(\mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1224_ (.A(\mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0364_),
    .Z(\mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1225_ (.A(\mux_left_track_29.INVTX1_0_.out ),
    .TE_B(_0365_),
    .Z(\mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1226_ (.A(net135),
    .TE_B(_0366_),
    .Z(\mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1227_ (.A(\mux_left_track_11.INVTX1_2_.out ),
    .TE_B(_0367_),
    .Z(\mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1228_ (.A(\mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0368_),
    .Z(\mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1229_ (.A(\mux_left_track_31.INVTX1_0_.out ),
    .TE_B(_0369_),
    .Z(\mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1230_ (.A(net136),
    .TE_B(_0370_),
    .Z(\mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1231_ (.A(\mux_left_track_13.INVTX1_2_.out ),
    .TE_B(_0371_),
    .Z(\mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1232_ (.A(\mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0372_),
    .Z(\mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1233_ (.A(\mux_left_track_33.INVTX1_0_.out ),
    .TE_B(_0373_),
    .Z(\mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1234_ (.A(net137),
    .TE_B(_0374_),
    .Z(\mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1235_ (.A(\mux_left_track_15.INVTX1_2_.out ),
    .TE_B(_0375_),
    .Z(\mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1236_ (.A(\mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0376_),
    .Z(\mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1237_ (.A(\mux_left_track_35.INVTX1_0_.out ),
    .TE_B(_0377_),
    .Z(\mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(ccff_head),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(chanx_left_in[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(chanx_left_in[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(chanx_left_in[11]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(chanx_left_in[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(chanx_left_in[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(chanx_left_in[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(chanx_left_in[15]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(chanx_left_in[16]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(chanx_left_in[17]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(chanx_left_in[18]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(chanx_left_in[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(chanx_left_in[2]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(chanx_left_in[3]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(chanx_left_in[4]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(chanx_left_in[5]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(chanx_left_in[6]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(chanx_left_in[7]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(chanx_left_in[8]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(chanx_left_in[9]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(chany_top_in[0]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(chany_top_in[10]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(chany_top_in[11]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(chany_top_in[12]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(chany_top_in[13]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(chany_top_in[14]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(chany_top_in[15]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(chany_top_in[16]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(chany_top_in[17]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(chany_top_in[18]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(chany_top_in[1]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(chany_top_in[2]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(chany_top_in[3]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(chany_top_in[4]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(chany_top_in[5]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(chany_top_in[6]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(chany_top_in[7]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(chany_top_in[8]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(chany_top_in[9]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_),
    .X(net49));
 sky130_fd_sc_hd__dlymetal6s2s_1 input50 (.A(pReset),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_),
    .X(net60));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(ccff_tail));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(chanx_left_out[0]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(chanx_left_out[10]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(chanx_left_out[11]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(chanx_left_out[12]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(chanx_left_out[13]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(chanx_left_out[14]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(chanx_left_out[15]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(chanx_left_out[16]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(chanx_left_out[17]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(chanx_left_out[18]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(chanx_left_out[1]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(chanx_left_out[2]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(chanx_left_out[3]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(chanx_left_out[4]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(chanx_left_out[5]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(chanx_left_out[6]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(chanx_left_out[7]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(chanx_left_out[8]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(chanx_left_out[9]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(chany_top_out[0]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(chany_top_out[10]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(chany_top_out[11]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(chany_top_out[12]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(chany_top_out[13]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(chany_top_out[14]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(chany_top_out[15]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(chany_top_out[16]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(chany_top_out[17]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(chany_top_out[18]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(chany_top_out[1]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(chany_top_out[2]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(chany_top_out[3]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(chany_top_out[4]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(chany_top_out[5]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(chany_top_out[6]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(chany_top_out[7]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(chany_top_out[8]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(chany_top_out[9]));
 sky130_fd_sc_hd__conb_1 _1043__100 (.HI(net100));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_3_0__leaf_prog_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_3_1__leaf_prog_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_3_2__leaf_prog_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_3_3__leaf_prog_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_3_4__leaf_prog_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_3_5__leaf_prog_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_3_6__leaf_prog_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_prog_clk (.A(clknet_0_prog_clk),
    .X(clknet_3_7__leaf_prog_clk));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_405 ();
endmodule

